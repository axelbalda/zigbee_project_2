
module MSK_MODULATOR ( clk, reset, i_empty, i_data, o_ready, o_sinI, o_sinQ );
  output [3:0] o_sinI;
  output [3:0] o_sinQ;
  input clk, reset, i_empty, i_data;
  output o_ready;
  wire   clk_10M, N459, N460, N461, N462, N463, N464, N465, N466, N467, N468,
         N469, N470, N471, N472, N473, N474, N475, N476, \stateI[0] ,
         \stateQ[0] , IorQ, sin_was_positiveI, sin_was_positiveQ, isPositiveI,
         isPositiveQ, is9, old_i_data, my_clk_10M, N499, N501, N503, N504,
         N505, N506, N507, N508, N509, N510, N511, N512, N513, N514, N515,
         N516, N517, N518, N519, N520, N521, N522, N563, N564, N652, N692,
         N693, N694, N695, N696, N697, N698, N699, N700, N701, N702, N703,
         N704, N705, N706, N707, N708, N709, N767, N768, N769, N770, N771,
         N772, N773, N774, N775, N776, N777, N778, N779, N780, N781, N782,
         N783, N784, N785, N786, N787, N790, N791, N792, N793, N794, N795,
         N934, N974, N975, N976, N977, N978, N979, N980, N981, N982, N983,
         N984, N985, N986, N987, N988, N989, N990, N991, N1050, N1051, N1052,
         N1053, N1054, N1055, N1056, N1057, N1058, N1059, N1060, N1061, N1062,
         N1063, N1064, N1065, N1066, N1067, N1068, N1069, N1070, N1071, N1072,
         N1073, N1075, N1076, N1077, N1078, N1079, N1080, N1081, N1083, N1084,
         N1085, N1092, N1098, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n232, n233, n234, n235, n236, n237, n238,
         n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249,
         n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260,
         n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271,
         n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282,
         n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293,
         n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417;
  wire   [19:0] c;
  wire   [19:0] i;
  wire   [19:0] j;
  wire   [19:2] \add_236/carry ;
  wire   [19:2] \add_173/carry ;
  wire   [19:2] \add_78/carry ;

  OAI222 U12 ( .A(n295), .B(n278), .C(n132), .D(n133), .Q(N795) );
  OAI222 U14 ( .A(n135), .B(n278), .C(n136), .D(n378), .Q(N794) );
  OAI222 U16 ( .A(n139), .B(n140), .C(n141), .D(n142), .Q(n138) );
  OAI222 U17 ( .A(n143), .B(n144), .C(n145), .D(n378), .Q(n137) );
  OAI222 U18 ( .A(n139), .B(n133), .C(n141), .D(n147), .Q(n146) );
  OAI222 U20 ( .A(n148), .B(n278), .C(n136), .D(n374), .Q(N793) );
  OAI222 U24 ( .A(n153), .B(n140), .C(n154), .D(n142), .Q(n150) );
  OAI222 U25 ( .A(n153), .B(n133), .C(n154), .D(n147), .Q(n149) );
  OAI212 U34 ( .A(n143), .B(n144), .C(n140), .Q(n134) );
  OAI212 U38 ( .A(n278), .B(n144), .C(n166), .Q(N791) );
  OAI212 U111 ( .A(n254), .B(n188), .C(n189), .Q(N1085) );
  OAI222 U129 ( .A(n294), .B(n319), .C(n206), .D(n207), .Q(N1079) );
  OAI212 U130 ( .A(n203), .B(n209), .C(n210), .Q(N1078) );
  OAI212 U131 ( .A(n211), .B(n212), .C(n203), .Q(n210) );
  OAI222 U132 ( .A(n213), .B(n214), .C(n215), .D(n216), .Q(n212) );
  OAI222 U133 ( .A(n323), .B(n209), .C(n217), .D(n218), .Q(n211) );
  OAI222 U136 ( .A(n203), .B(n344), .C(n219), .D(n319), .Q(N1077) );
  OAI222 U139 ( .A(n224), .B(n214), .C(n225), .D(n216), .Q(n222) );
  OAI222 U140 ( .A(n224), .B(n207), .C(n225), .D(n226), .Q(n220) );
  OAI212 U149 ( .A(n217), .B(n218), .C(n214), .Q(n208) );
  OAI212 U155 ( .A(n385), .B(n384), .C(n130), .Q(n237) );
  OAI212 U165 ( .A(n206), .B(n188), .C(n189), .Q(N1072) );
  ADD22 \add_236/U1_1_1  ( .A(n272), .B(j[0]), .CO(\add_236/carry [2]), .S(
        N974) );
  ADD22 \add_236/U1_1_2  ( .A(j[2]), .B(\add_236/carry [2]), .CO(
        \add_236/carry [3]), .S(N975) );
  ADD22 \add_236/U1_1_3  ( .A(n251), .B(\add_236/carry [3]), .CO(
        \add_236/carry [4]), .S(N976) );
  ADD22 \add_236/U1_1_4  ( .A(j[4]), .B(\add_236/carry [4]), .CO(
        \add_236/carry [5]), .S(N977) );
  ADD22 \add_236/U1_1_5  ( .A(j[5]), .B(\add_236/carry [5]), .CO(
        \add_236/carry [6]), .S(N978) );
  ADD22 \add_236/U1_1_6  ( .A(j[6]), .B(\add_236/carry [6]), .CO(
        \add_236/carry [7]), .S(N979) );
  ADD22 \add_236/U1_1_7  ( .A(j[7]), .B(\add_236/carry [7]), .CO(
        \add_236/carry [8]), .S(N980) );
  ADD22 \add_236/U1_1_8  ( .A(j[8]), .B(\add_236/carry [8]), .CO(
        \add_236/carry [9]), .S(N981) );
  ADD22 \add_236/U1_1_9  ( .A(j[9]), .B(\add_236/carry [9]), .CO(
        \add_236/carry [10]), .S(N982) );
  ADD22 \add_236/U1_1_10  ( .A(j[10]), .B(\add_236/carry [10]), .CO(
        \add_236/carry [11]), .S(N983) );
  ADD22 \add_236/U1_1_11  ( .A(j[11]), .B(\add_236/carry [11]), .CO(
        \add_236/carry [12]), .S(N984) );
  ADD22 \add_236/U1_1_12  ( .A(j[12]), .B(\add_236/carry [12]), .CO(
        \add_236/carry [13]), .S(N985) );
  ADD22 \add_236/U1_1_13  ( .A(j[13]), .B(\add_236/carry [13]), .CO(
        \add_236/carry [14]), .S(N986) );
  ADD22 \add_236/U1_1_14  ( .A(j[14]), .B(\add_236/carry [14]), .CO(
        \add_236/carry [15]), .S(N987) );
  ADD22 \add_236/U1_1_15  ( .A(j[15]), .B(\add_236/carry [15]), .CO(
        \add_236/carry [16]), .S(N988) );
  ADD22 \add_236/U1_1_16  ( .A(j[16]), .B(\add_236/carry [16]), .CO(
        \add_236/carry [17]), .S(N989) );
  ADD22 \add_236/U1_1_17  ( .A(j[17]), .B(\add_236/carry [17]), .CO(
        \add_236/carry [18]), .S(N990) );
  ADD22 \add_236/U1_1_18  ( .A(j[18]), .B(\add_236/carry [18]), .CO(
        \add_236/carry [19]), .S(N991) );
  ADD22 \add_173/U1_1_1  ( .A(n270), .B(n271), .CO(\add_173/carry [2]), .S(
        N692) );
  ADD22 \add_173/U1_1_2  ( .A(i[2]), .B(\add_173/carry [2]), .CO(
        \add_173/carry [3]), .S(N693) );
  ADD22 \add_173/U1_1_3  ( .A(n269), .B(\add_173/carry [3]), .CO(
        \add_173/carry [4]), .S(N694) );
  ADD22 \add_173/U1_1_4  ( .A(i[4]), .B(\add_173/carry [4]), .CO(
        \add_173/carry [5]), .S(N695) );
  ADD22 \add_173/U1_1_5  ( .A(i[5]), .B(\add_173/carry [5]), .CO(
        \add_173/carry [6]), .S(N696) );
  ADD22 \add_173/U1_1_6  ( .A(i[6]), .B(\add_173/carry [6]), .CO(
        \add_173/carry [7]), .S(N697) );
  ADD22 \add_173/U1_1_7  ( .A(i[7]), .B(\add_173/carry [7]), .CO(
        \add_173/carry [8]), .S(N698) );
  ADD22 \add_173/U1_1_8  ( .A(i[8]), .B(\add_173/carry [8]), .CO(
        \add_173/carry [9]), .S(N699) );
  ADD22 \add_173/U1_1_9  ( .A(i[9]), .B(\add_173/carry [9]), .CO(
        \add_173/carry [10]), .S(N700) );
  ADD22 \add_173/U1_1_10  ( .A(i[10]), .B(\add_173/carry [10]), .CO(
        \add_173/carry [11]), .S(N701) );
  ADD22 \add_173/U1_1_11  ( .A(i[11]), .B(\add_173/carry [11]), .CO(
        \add_173/carry [12]), .S(N702) );
  ADD22 \add_173/U1_1_12  ( .A(i[12]), .B(\add_173/carry [12]), .CO(
        \add_173/carry [13]), .S(N703) );
  ADD22 \add_173/U1_1_13  ( .A(i[13]), .B(\add_173/carry [13]), .CO(
        \add_173/carry [14]), .S(N704) );
  ADD22 \add_173/U1_1_14  ( .A(i[14]), .B(\add_173/carry [14]), .CO(
        \add_173/carry [15]), .S(N705) );
  ADD22 \add_173/U1_1_15  ( .A(i[15]), .B(\add_173/carry [15]), .CO(
        \add_173/carry [16]), .S(N706) );
  ADD22 \add_173/U1_1_16  ( .A(i[16]), .B(\add_173/carry [16]), .CO(
        \add_173/carry [17]), .S(N707) );
  ADD22 \add_173/U1_1_17  ( .A(i[17]), .B(\add_173/carry [17]), .CO(
        \add_173/carry [18]), .S(N708) );
  ADD22 \add_173/U1_1_18  ( .A(i[18]), .B(\add_173/carry [18]), .CO(
        \add_173/carry [19]), .S(N709) );
  ADD22 \add_78/U1_1_1  ( .A(c[1]), .B(c[0]), .CO(\add_78/carry [2]), .S(N459)
         );
  ADD22 \add_78/U1_1_2  ( .A(c[2]), .B(\add_78/carry [2]), .CO(
        \add_78/carry [3]), .S(N460) );
  ADD22 \add_78/U1_1_3  ( .A(c[3]), .B(\add_78/carry [3]), .CO(
        \add_78/carry [4]), .S(N461) );
  ADD22 \add_78/U1_1_4  ( .A(c[4]), .B(\add_78/carry [4]), .CO(
        \add_78/carry [5]), .S(N462) );
  ADD22 \add_78/U1_1_5  ( .A(c[5]), .B(\add_78/carry [5]), .CO(
        \add_78/carry [6]), .S(N463) );
  ADD22 \add_78/U1_1_6  ( .A(c[6]), .B(\add_78/carry [6]), .CO(
        \add_78/carry [7]), .S(N464) );
  ADD22 \add_78/U1_1_7  ( .A(c[7]), .B(\add_78/carry [7]), .CO(
        \add_78/carry [8]), .S(N465) );
  ADD22 \add_78/U1_1_8  ( .A(c[8]), .B(\add_78/carry [8]), .CO(
        \add_78/carry [9]), .S(N466) );
  ADD22 \add_78/U1_1_9  ( .A(c[9]), .B(\add_78/carry [9]), .CO(
        \add_78/carry [10]), .S(N467) );
  ADD22 \add_78/U1_1_10  ( .A(c[10]), .B(\add_78/carry [10]), .CO(
        \add_78/carry [11]), .S(N468) );
  ADD22 \add_78/U1_1_11  ( .A(c[11]), .B(\add_78/carry [11]), .CO(
        \add_78/carry [12]), .S(N469) );
  ADD22 \add_78/U1_1_12  ( .A(c[12]), .B(\add_78/carry [12]), .CO(
        \add_78/carry [13]), .S(N470) );
  ADD22 \add_78/U1_1_13  ( .A(c[13]), .B(\add_78/carry [13]), .CO(
        \add_78/carry [14]), .S(N471) );
  ADD22 \add_78/U1_1_14  ( .A(c[14]), .B(\add_78/carry [14]), .CO(
        \add_78/carry [15]), .S(N472) );
  ADD22 \add_78/U1_1_15  ( .A(c[15]), .B(\add_78/carry [15]), .CO(
        \add_78/carry [16]), .S(N473) );
  ADD22 \add_78/U1_1_16  ( .A(c[16]), .B(\add_78/carry [16]), .CO(
        \add_78/carry [17]), .S(N474) );
  ADD22 \add_78/U1_1_17  ( .A(c[17]), .B(\add_78/carry [17]), .CO(
        \add_78/carry [18]), .S(N475) );
  ADD22 \add_78/U1_1_18  ( .A(c[18]), .B(\add_78/carry [18]), .CO(
        \add_78/carry [19]), .S(N476) );
  DF3 \c_reg[0]  ( .D(N503), .C(clk), .Q(c[0]), .QN(n261) );
  DF3 \c_reg[1]  ( .D(N504), .C(clk), .Q(c[1]) );
  DF3 \c_reg[2]  ( .D(N505), .C(clk), .Q(c[2]) );
  DF3 \c_reg[3]  ( .D(N506), .C(clk), .Q(c[3]) );
  DF3 \c_reg[4]  ( .D(N507), .C(clk), .Q(c[4]) );
  DF3 \c_reg[5]  ( .D(N508), .C(clk), .Q(c[5]) );
  DF3 \c_reg[6]  ( .D(N509), .C(clk), .Q(c[6]) );
  DF3 \c_reg[7]  ( .D(N510), .C(clk), .Q(c[7]) );
  DF3 \c_reg[8]  ( .D(N511), .C(clk), .Q(c[8]) );
  DF3 \c_reg[9]  ( .D(N512), .C(clk), .Q(c[9]) );
  DF3 \c_reg[10]  ( .D(N513), .C(clk), .Q(c[10]) );
  DF3 \c_reg[11]  ( .D(N514), .C(clk), .Q(c[11]) );
  DF3 \c_reg[12]  ( .D(N515), .C(clk), .Q(c[12]) );
  DF3 \c_reg[13]  ( .D(N516), .C(clk), .Q(c[13]) );
  DF3 \c_reg[14]  ( .D(N517), .C(clk), .Q(c[14]) );
  DF3 \c_reg[15]  ( .D(N518), .C(clk), .Q(c[15]) );
  DF3 \c_reg[16]  ( .D(N519), .C(clk), .Q(c[16]) );
  DF3 \c_reg[17]  ( .D(N520), .C(clk), .Q(c[17]) );
  DF3 \c_reg[18]  ( .D(N521), .C(clk), .Q(c[18]) );
  DF3 \c_reg[19]  ( .D(N522), .C(clk), .Q(c[19]) );
  DF3 clk_10M_reg ( .D(n314), .C(clk), .Q(clk_10M) );
  DF3 \stateQ_reg[0]  ( .D(N501), .C(clk), .Q(\stateQ[0] ), .QN(n254) );
  DF3 \stateI_reg[0]  ( .D(N499), .C(clk), .Q(\stateI[0] ), .QN(n257) );
  DFE1 \next_stateQ_reg[0]  ( .D(N1098), .E(n316), .C(clk), .QN(n265) );
  DFE1 \next_stateI_reg[0]  ( .D(N1092), .E(n317), .C(clk), .QN(n264) );
  DFE1 sin_was_positiveQ_reg ( .D(n291), .E(n287), .C(clk), .Q(
        sin_was_positiveQ) );
  DFE1 sin_was_positiveI_reg ( .D(N564), .E(N563), .C(clk), .Q(
        sin_was_positiveI) );
  DFE1 old_i_data_reg ( .D(N1081), .E(N1080), .C(clk), .Q(old_i_data) );
  DFE1 my_clk_10M_reg ( .D(clk_10M), .E(reset), .C(clk), .Q(my_clk_10M), .QN(
        n250) );
  DFE1 isPositiveI_reg ( .D(N790), .E(n286), .C(clk), .Q(isPositiveI), .QN(
        n259) );
  DFE1 is9_reg ( .D(N1085), .E(N1084), .C(clk), .Q(is9) );
  DFE1 \j_reg[16]  ( .D(N1067), .E(N1050), .C(clk), .Q(j[16]) );
  DFE1 \i_reg[16]  ( .D(N784), .E(N767), .C(clk), .Q(i[16]) );
  DFE1 \j_reg[15]  ( .D(N1066), .E(n277), .C(clk), .Q(j[15]) );
  DFE1 \i_reg[15]  ( .D(N783), .E(n284), .C(clk), .Q(i[15]) );
  DFE1 \j_reg[17]  ( .D(N1068), .E(n277), .C(clk), .Q(j[17]) );
  DFE1 \i_reg[17]  ( .D(N785), .E(n284), .C(clk), .Q(i[17]) );
  DFE1 \j_reg[18]  ( .D(N1069), .E(N1050), .C(clk), .Q(j[18]) );
  DFE1 \i_reg[18]  ( .D(N786), .E(N767), .C(clk), .Q(i[18]) );
  DFE1 \j_reg[19]  ( .D(N1070), .E(n277), .C(clk), .Q(j[19]) );
  DFE1 \i_reg[19]  ( .D(N787), .E(n284), .C(clk), .Q(i[19]) );
  DFE1 isPositiveQ_reg ( .D(n293), .E(N1073), .C(clk), .Q(isPositiveQ), .QN(
        n260) );
  DFE1 IorQ_reg ( .D(N1083), .E(n285), .C(clk), .Q(IorQ), .QN(n263) );
  DFE1 \j_reg[12]  ( .D(N1063), .E(N1050), .C(clk), .Q(j[12]) );
  DFE1 \i_reg[12]  ( .D(N780), .E(N767), .C(clk), .Q(i[12]) );
  DFE1 \j_reg[14]  ( .D(N1065), .E(N1050), .C(clk), .Q(j[14]) );
  DFE1 \i_reg[14]  ( .D(N782), .E(N767), .C(clk), .Q(i[14]) );
  DFE1 \j_reg[13]  ( .D(N1064), .E(n277), .C(clk), .Q(j[13]) );
  DFE1 \i_reg[13]  ( .D(N781), .E(n284), .C(clk), .Q(i[13]) );
  DFE1 \j_reg[10]  ( .D(N1061), .E(N1050), .C(clk), .Q(j[10]) );
  DFE1 \j_reg[11]  ( .D(N1062), .E(n277), .C(clk), .Q(j[11]) );
  DFE1 \i_reg[10]  ( .D(N778), .E(N767), .C(clk), .Q(i[10]) );
  DFE1 \i_reg[11]  ( .D(N779), .E(n284), .C(clk), .Q(i[11]) );
  DFE1 \j_reg[9]  ( .D(N1060), .E(n277), .C(clk), .Q(j[9]) );
  DFE1 \i_reg[9]  ( .D(N777), .E(n284), .C(clk), .Q(i[9]) );
  DFE1 \j_reg[7]  ( .D(N1058), .E(n277), .C(clk), .Q(j[7]) );
  DFE1 \j_reg[8]  ( .D(N1059), .E(N1050), .C(clk), .Q(j[8]) );
  DFE1 \i_reg[7]  ( .D(N775), .E(n284), .C(clk), .Q(i[7]) );
  DFE1 \i_reg[8]  ( .D(N776), .E(N767), .C(clk), .Q(i[8]) );
  DFE1 \j_reg[4]  ( .D(N1055), .E(N1050), .C(clk), .Q(j[4]) );
  DFE1 \j_reg[5]  ( .D(N1056), .E(n277), .C(clk), .Q(j[5]) );
  DFE1 \i_reg[4]  ( .D(N772), .E(N767), .C(clk), .Q(i[4]) );
  DFE1 \i_reg[5]  ( .D(N773), .E(n284), .C(clk), .Q(i[5]) );
  DFE1 \j_reg[6]  ( .D(N1057), .E(N1050), .C(clk), .Q(j[6]) );
  DFE1 \i_reg[6]  ( .D(N774), .E(N767), .C(clk), .Q(i[6]) );
  DFE1 \j_reg[1]  ( .D(N1052), .E(n277), .C(clk), .Q(j[1]) );
  DFE1 \i_reg[1]  ( .D(N769), .E(n284), .C(clk), .Q(i[1]) );
  DFE1 \i_reg[3]  ( .D(N771), .E(n284), .C(clk), .Q(i[3]), .QN(n256) );
  DFE1 \j_reg[3]  ( .D(N1054), .E(n277), .C(clk), .Q(n251), .QN(n262) );
  DFE1 \i_reg[2]  ( .D(N770), .E(N767), .C(clk), .Q(i[2]), .QN(n258) );
  DFE1 \j_reg[2]  ( .D(N1053), .E(N1050), .C(clk), .Q(j[2]), .QN(n255) );
  DFE1 \j_reg[0]  ( .D(N1051), .E(N1050), .C(clk), .Q(j[0]), .QN(n253) );
  DFE1 \i_reg[0]  ( .D(N768), .E(N767), .C(clk), .Q(i[0]), .QN(n252) );
  DFE1 \o_sinQ_reg[0]  ( .D(N1076), .E(N1075), .C(clk), .Q(o_sinQ[0]) );
  DFE1 \o_sinI_reg[0]  ( .D(N792), .E(N791), .C(clk), .Q(o_sinI[0]) );
  DFE1 \o_sinI_reg[1]  ( .D(N793), .E(N791), .C(clk), .Q(o_sinI[1]) );
  DFE1 \o_sinI_reg[2]  ( .D(N794), .E(N791), .C(clk), .Q(o_sinI[2]) );
  DFE1 \o_sinI_reg[3]  ( .D(N795), .E(N791), .C(clk), .Q(o_sinI[3]) );
  DFE1 \o_sinQ_reg[1]  ( .D(N1077), .E(N1075), .C(clk), .Q(o_sinQ[1]) );
  DFE1 \o_sinQ_reg[2]  ( .D(N1078), .E(N1075), .C(clk), .Q(o_sinQ[2]) );
  DFE1 \o_sinQ_reg[3]  ( .D(N1079), .E(N1075), .C(clk), .Q(o_sinQ[3]) );
  DFE1 o_ready_reg ( .D(N1072), .E(N1071), .C(clk), .Q(o_ready) );
  NOR21 U335 ( .A(n281), .B(n266), .Q(N787) );
  NOR21 U336 ( .A(n274), .B(n267), .Q(N1070) );
  NOR21 U337 ( .A(n173), .B(n268), .Q(N522) );
  NAND22 U338 ( .A(n187), .B(n136), .Q(n188) );
  INV3 U339 ( .A(n206), .Q(n318) );
  NAND22 U340 ( .A(n320), .B(n323), .Q(n218) );
  NAND22 U341 ( .A(n351), .B(n145), .Q(n144) );
  INV3 U342 ( .A(n167), .Q(n351) );
  NOR21 U343 ( .A(n221), .B(n319), .Q(n206) );
  INV3 U344 ( .A(n203), .Q(n319) );
  AOI221 U345 ( .A(n347), .B(n385), .C(n346), .D(n384), .Q(n209) );
  INV3 U346 ( .A(n213), .Q(n347) );
  NAND41 U347 ( .A(n318), .B(n189), .C(n188), .D(n170), .Q(N1071) );
  NAND22 U348 ( .A(n203), .B(n184), .Q(n189) );
  NAND22 U349 ( .A(n274), .B(n131), .Q(N1050) );
  NAND22 U350 ( .A(n273), .B(n131), .Q(n277) );
  NAND22 U351 ( .A(n281), .B(n289), .Q(N767) );
  NAND22 U352 ( .A(n280), .B(n289), .Q(n284) );
  NOR21 U353 ( .A(n262), .B(n204), .Q(n184) );
  INV3 U354 ( .A(n145), .Q(n354) );
  NOR21 U355 ( .A(n204), .B(n251), .Q(n201) );
  NOR21 U356 ( .A(n205), .B(n256), .Q(n187) );
  INV3 U357 ( .A(n221), .Q(n323) );
  NOR21 U358 ( .A(n274), .B(n341), .Q(N1054) );
  INV3 U359 ( .A(N976), .Q(n341) );
  NOR21 U360 ( .A(n281), .B(n371), .Q(N771) );
  INV3 U361 ( .A(N694), .Q(n371) );
  NOR21 U362 ( .A(n276), .B(n343), .Q(N1052) );
  INV3 U363 ( .A(N974), .Q(n343) );
  NOR21 U364 ( .A(n283), .B(n373), .Q(N769) );
  INV3 U365 ( .A(N692), .Q(n373) );
  INV3 U366 ( .A(n170), .Q(n286) );
  INV3 U367 ( .A(n131), .Q(n287) );
  NOR21 U368 ( .A(n173), .B(n297), .Q(N520) );
  INV3 U369 ( .A(N475), .Q(n297) );
  NOR21 U370 ( .A(n276), .B(n327), .Q(N1068) );
  INV3 U371 ( .A(N990), .Q(n327) );
  NOR21 U372 ( .A(n275), .B(n328), .Q(N1067) );
  INV3 U373 ( .A(N989), .Q(n328) );
  NOR21 U374 ( .A(n283), .B(n357), .Q(N785) );
  INV3 U375 ( .A(N708), .Q(n357) );
  NOR21 U376 ( .A(n282), .B(n358), .Q(N784) );
  INV3 U377 ( .A(N707), .Q(n358) );
  NOR21 U378 ( .A(n280), .B(n356), .Q(N786) );
  INV3 U379 ( .A(N709), .Q(n356) );
  NOR21 U380 ( .A(n273), .B(n326), .Q(N1069) );
  INV3 U381 ( .A(N991), .Q(n326) );
  NOR21 U382 ( .A(n279), .B(n296), .Q(N521) );
  INV3 U383 ( .A(N476), .Q(n296) );
  NOR21 U384 ( .A(n279), .B(n298), .Q(N519) );
  INV3 U385 ( .A(N474), .Q(n298) );
  NOR21 U386 ( .A(n279), .B(n300), .Q(N517) );
  INV3 U387 ( .A(N472), .Q(n300) );
  NOR21 U388 ( .A(n274), .B(n331), .Q(N1064) );
  INV3 U389 ( .A(N986), .Q(n331) );
  NOR21 U390 ( .A(n281), .B(n361), .Q(N781) );
  INV3 U391 ( .A(N704), .Q(n361) );
  NOR21 U392 ( .A(n276), .B(n329), .Q(N1066) );
  INV3 U393 ( .A(N988), .Q(n329) );
  NOR21 U394 ( .A(n275), .B(n330), .Q(N1065) );
  INV3 U395 ( .A(N987), .Q(n330) );
  NOR21 U396 ( .A(n283), .B(n359), .Q(N783) );
  INV3 U397 ( .A(N706), .Q(n359) );
  NOR21 U398 ( .A(n282), .B(n360), .Q(N782) );
  INV3 U399 ( .A(N705), .Q(n360) );
  NOR21 U400 ( .A(n173), .B(n299), .Q(N518) );
  INV3 U401 ( .A(N473), .Q(n299) );
  NOR21 U402 ( .A(n173), .B(n301), .Q(N516) );
  INV3 U403 ( .A(N471), .Q(n301) );
  NOR21 U404 ( .A(n281), .B(n363), .Q(N779) );
  INV3 U405 ( .A(N702), .Q(n363) );
  NOR21 U406 ( .A(n274), .B(n333), .Q(N1062) );
  INV3 U407 ( .A(N984), .Q(n333) );
  NOR21 U408 ( .A(n280), .B(n362), .Q(N780) );
  INV3 U409 ( .A(N703), .Q(n362) );
  NOR21 U410 ( .A(n273), .B(n332), .Q(N1063) );
  INV3 U411 ( .A(N985), .Q(n332) );
  NOR21 U412 ( .A(n279), .B(n302), .Q(N515) );
  INV3 U413 ( .A(N470), .Q(n302) );
  NOR21 U414 ( .A(n173), .B(n305), .Q(N512) );
  INV3 U415 ( .A(N467), .Q(n305) );
  NOR21 U416 ( .A(n275), .B(n336), .Q(N1059) );
  INV3 U417 ( .A(N981), .Q(n336) );
  NOR21 U418 ( .A(n282), .B(n366), .Q(N776) );
  INV3 U419 ( .A(N699), .Q(n366) );
  NOR21 U420 ( .A(n280), .B(n364), .Q(N778) );
  INV3 U421 ( .A(N701), .Q(n364) );
  NOR21 U422 ( .A(n283), .B(n365), .Q(N777) );
  INV3 U423 ( .A(N700), .Q(n365) );
  NOR21 U424 ( .A(n273), .B(n334), .Q(N1061) );
  INV3 U425 ( .A(N983), .Q(n334) );
  NOR21 U426 ( .A(n276), .B(n335), .Q(N1060) );
  INV3 U427 ( .A(N982), .Q(n335) );
  NOR21 U428 ( .A(n173), .B(n303), .Q(N514) );
  INV3 U429 ( .A(N469), .Q(n303) );
  NOR21 U430 ( .A(n279), .B(n304), .Q(N513) );
  INV3 U431 ( .A(N468), .Q(n304) );
  AOI211 U432 ( .A(n136), .B(n167), .C(n168), .Q(n166) );
  AOI211 U433 ( .A(n147), .B(n133), .C(n169), .Q(n168) );
  NAND22 U434 ( .A(N652), .B(n259), .Q(n140) );
  INV3 U435 ( .A(n220), .Q(n344) );
  AOI2111 U436 ( .A(n220), .B(n221), .C(n222), .D(n223), .Q(n219) );
  OAI311 U437 ( .A(n250), .B(n159), .C(n257), .D(n161), .Q(N792) );
  AOI221 U438 ( .A(n383), .B(n162), .C(n382), .D(n162), .Q(n161) );
  AOI221 U439 ( .A(n163), .B(n162), .C(n162), .D(n134), .Q(n159) );
  INV3 U440 ( .A(n147), .Q(n382) );
  NOR21 U441 ( .A(n137), .B(n138), .Q(n135) );
  NAND22 U442 ( .A(n142), .B(n140), .Q(n167) );
  NOR21 U443 ( .A(n217), .B(n218), .Q(n223) );
  NOR21 U444 ( .A(n279), .B(n306), .Q(N511) );
  INV3 U445 ( .A(N466), .Q(n306) );
  NOR21 U446 ( .A(n173), .B(n307), .Q(N510) );
  INV3 U447 ( .A(N465), .Q(n307) );
  INV3 U448 ( .A(n238), .Q(n320) );
  NAND22 U449 ( .A(n216), .B(n214), .Q(n238) );
  NAND22 U450 ( .A(n142), .B(n144), .Q(n163) );
  NAND22 U451 ( .A(n216), .B(n218), .Q(n235) );
  NOR21 U452 ( .A(n274), .B(n339), .Q(N1056) );
  INV3 U453 ( .A(N978), .Q(n339) );
  NOR21 U454 ( .A(n281), .B(n369), .Q(N773) );
  INV3 U455 ( .A(N696), .Q(n369) );
  NOR21 U456 ( .A(n276), .B(n337), .Q(N1058) );
  INV3 U457 ( .A(N980), .Q(n337) );
  NOR21 U458 ( .A(n275), .B(n338), .Q(N1057) );
  INV3 U459 ( .A(N979), .Q(n338) );
  NOR21 U460 ( .A(n283), .B(n367), .Q(N775) );
  INV3 U461 ( .A(N698), .Q(n367) );
  NOR21 U462 ( .A(n282), .B(n368), .Q(N774) );
  INV3 U463 ( .A(N697), .Q(n368) );
  NOR21 U464 ( .A(n279), .B(n308), .Q(N509) );
  INV3 U465 ( .A(N464), .Q(n308) );
  NOR21 U466 ( .A(n254), .B(n250), .Q(n203) );
  OAI2111 U467 ( .A(n320), .B(n319), .C(n318), .D(n237), .Q(N1075) );
  NAND31 U468 ( .A(n353), .B(n141), .C(n271), .Q(n205) );
  INV3 U469 ( .A(n197), .Q(n353) );
  NAND31 U470 ( .A(n324), .B(n215), .C(j[0]), .Q(n204) );
  NAND31 U471 ( .A(n252), .B(n256), .C(n141), .Q(n158) );
  AOI211 U472 ( .A(n145), .B(n136), .C(n288), .Q(n170) );
  AOI2111 U473 ( .A(n252), .B(n269), .C(n155), .D(n375), .Q(n154) );
  AOI211 U474 ( .A(n271), .B(n270), .C(n258), .Q(n155) );
  INV3 U475 ( .A(n156), .Q(n375) );
  AOI311 U476 ( .A(n271), .B(n258), .C(n270), .D(n157), .Q(n156) );
  AOI2111 U477 ( .A(n253), .B(n251), .C(n227), .D(n345), .Q(n225) );
  AOI211 U478 ( .A(j[0]), .B(n272), .C(n255), .Q(n227) );
  INV3 U479 ( .A(n228), .Q(n345) );
  AOI311 U480 ( .A(j[0]), .B(n255), .C(n272), .D(n229), .Q(n228) );
  INV3 U481 ( .A(n146), .Q(n378) );
  NOR21 U482 ( .A(n158), .B(n197), .Q(n145) );
  AOI2111 U483 ( .A(n271), .B(n269), .C(n376), .D(n270), .Q(n153) );
  INV3 U484 ( .A(n158), .Q(n376) );
  NAND22 U485 ( .A(n230), .B(n324), .Q(n221) );
  AOI2111 U486 ( .A(j[0]), .B(n251), .C(n230), .D(n272), .Q(n224) );
  NOR31 U487 ( .A(n258), .B(n197), .C(n377), .Q(n193) );
  INV3 U488 ( .A(n198), .Q(n377) );
  NOR31 U489 ( .A(n271), .B(n269), .C(n270), .Q(n198) );
  INV3 U490 ( .A(n208), .Q(n294) );
  NOR21 U491 ( .A(n354), .B(n278), .Q(n132) );
  INV3 U492 ( .A(n134), .Q(n295) );
  INV3 U493 ( .A(n149), .Q(n374) );
  AOI2111 U494 ( .A(n149), .B(n354), .C(n150), .D(n151), .Q(n148) );
  NOR31 U495 ( .A(j[0]), .B(n251), .C(n346), .Q(n230) );
  NOR21 U496 ( .A(n215), .B(n251), .Q(n213) );
  NOR21 U497 ( .A(n205), .B(n269), .Q(n200) );
  NOR31 U498 ( .A(n164), .B(n354), .C(n278), .Q(N790) );
  NOR21 U499 ( .A(n141), .B(n269), .Q(n139) );
  NOR31 U500 ( .A(n252), .B(n269), .C(n270), .Q(n157) );
  BUF2 U501 ( .A(n249), .Q(n273) );
  BUF2 U502 ( .A(n249), .Q(n274) );
  BUF2 U503 ( .A(n171), .Q(n280) );
  BUF2 U504 ( .A(n171), .Q(n281) );
  NOR31 U505 ( .A(n253), .B(n251), .C(n272), .Q(n229) );
  NOR21 U506 ( .A(n173), .B(n309), .Q(N508) );
  INV3 U507 ( .A(N463), .Q(n309) );
  NOR21 U508 ( .A(n279), .B(n310), .Q(N507) );
  INV3 U509 ( .A(N462), .Q(n310) );
  NOR21 U510 ( .A(n173), .B(n311), .Q(N506) );
  INV3 U511 ( .A(N461), .Q(n311) );
  NOR21 U512 ( .A(n279), .B(n312), .Q(N505) );
  INV3 U513 ( .A(N460), .Q(n312) );
  NOR21 U514 ( .A(n173), .B(n313), .Q(N504) );
  INV3 U515 ( .A(N459), .Q(n313) );
  BUF2 U516 ( .A(n249), .Q(n276) );
  BUF2 U517 ( .A(n249), .Q(n275) );
  BUF2 U518 ( .A(n171), .Q(n283) );
  BUF2 U519 ( .A(n171), .Q(n282) );
  INV3 U520 ( .A(n226), .Q(n384) );
  INV3 U521 ( .A(n207), .Q(n385) );
  NOR21 U522 ( .A(n143), .B(n144), .Q(n151) );
  INV3 U523 ( .A(n215), .Q(n346) );
  INV3 U524 ( .A(n136), .Q(n278) );
  NOR21 U525 ( .A(n250), .B(n257), .Q(n136) );
  NOR21 U526 ( .A(n273), .B(n340), .Q(N1055) );
  INV3 U527 ( .A(N977), .Q(n340) );
  NOR21 U528 ( .A(n273), .B(n342), .Q(N1053) );
  INV3 U529 ( .A(N975), .Q(n342) );
  NOR21 U530 ( .A(n280), .B(n370), .Q(N772) );
  INV3 U531 ( .A(N695), .Q(n370) );
  NOR21 U532 ( .A(n280), .B(n372), .Q(N770) );
  INV3 U533 ( .A(N693), .Q(n372) );
  INV3 U534 ( .A(n194), .Q(n285) );
  AOI2111 U535 ( .A(n136), .B(n193), .C(n195), .D(n288), .Q(n194) );
  NOR21 U536 ( .A(n191), .B(n319), .Q(n195) );
  INV3 U537 ( .A(n239), .Q(n293) );
  NAND22 U538 ( .A(n217), .B(n206), .Q(n239) );
  NOR21 U539 ( .A(n288), .B(n130), .Q(n131) );
  INV3 U540 ( .A(N563), .Q(n289) );
  NOR21 U541 ( .A(n259), .B(n169), .Q(N564) );
  INV3 U542 ( .A(n128), .Q(n314) );
  INV3 U543 ( .A(n133), .Q(n383) );
  BUF2 U544 ( .A(i[0]), .Q(n271) );
  XNR21 U545 ( .A(\add_173/carry [19]), .B(i[19]), .Q(n266) );
  XNR21 U546 ( .A(\add_236/carry [19]), .B(j[19]), .Q(n267) );
  BUF2 U547 ( .A(i[3]), .Q(n269) );
  BUF2 U548 ( .A(i[1]), .Q(n270) );
  BUF2 U549 ( .A(j[1]), .Q(n272) );
  XNR21 U550 ( .A(\add_78/carry [19]), .B(c[19]), .Q(n268) );
  NAND41 U551 ( .A(n403), .B(n402), .C(n401), .D(n400), .Q(N934) );
  NOR31 U552 ( .A(j[11]), .B(j[13]), .C(j[12]), .Q(n402) );
  NOR21 U553 ( .A(j[10]), .B(j[0]), .Q(n403) );
  NOR40 U554 ( .A(j[16]), .B(n350), .C(j[15]), .D(j[14]), .Q(n401) );
  NAND41 U555 ( .A(n394), .B(n393), .C(n392), .D(n391), .Q(N652) );
  NOR31 U556 ( .A(i[11]), .B(i[13]), .C(i[12]), .Q(n393) );
  NOR21 U557 ( .A(i[10]), .B(n271), .Q(n394) );
  NOR40 U558 ( .A(i[16]), .B(n381), .C(i[15]), .D(i[14]), .Q(n392) );
  NAND22 U559 ( .A(N934), .B(isPositiveQ), .Q(n216) );
  NAND22 U560 ( .A(N652), .B(isPositiveI), .Q(n142) );
  NOR40 U561 ( .A(n399), .B(n348), .C(n272), .D(j[19]), .Q(n400) );
  NAND22 U562 ( .A(n397), .B(n396), .Q(n399) );
  INV3 U563 ( .A(n398), .Q(n348) );
  NOR21 U564 ( .A(j[6]), .B(j[5]), .Q(n397) );
  NOR40 U565 ( .A(n390), .B(n379), .C(n270), .D(i[19]), .Q(n391) );
  NAND22 U566 ( .A(n388), .B(n387), .Q(n390) );
  INV3 U567 ( .A(n389), .Q(n379) );
  NOR21 U568 ( .A(i[6]), .B(i[5]), .Q(n388) );
  NAND22 U569 ( .A(N934), .B(n260), .Q(n214) );
  OAI311 U570 ( .A(n254), .B(n232), .C(n250), .D(n233), .Q(N1076) );
  AOI221 U571 ( .A(n385), .B(n234), .C(n384), .D(n234), .Q(n233) );
  AOI221 U572 ( .A(n235), .B(n234), .C(n234), .D(n208), .Q(n232) );
  OAI2111 U573 ( .A(j[0]), .B(j[2]), .C(n272), .D(n236), .Q(n234) );
  NOR31 U574 ( .A(j[2]), .B(j[4]), .C(n251), .Q(n398) );
  NOR31 U575 ( .A(i[2]), .B(i[4]), .C(n269), .Q(n389) );
  NOR31 U576 ( .A(j[7]), .B(j[9]), .C(j[8]), .Q(n396) );
  NOR31 U577 ( .A(i[7]), .B(i[9]), .C(i[8]), .Q(n387) );
  OAI2111 U578 ( .A(n271), .B(i[2]), .C(n270), .D(n165), .Q(n162) );
  AOI211 U579 ( .A(n271), .B(i[2]), .C(n269), .Q(n165) );
  NAND22 U580 ( .A(reset), .B(n128), .Q(n173) );
  NAND22 U581 ( .A(reset), .B(n128), .Q(n279) );
  NAND41 U582 ( .A(n174), .B(n175), .C(n176), .D(n177), .Q(n128) );
  NOR21 U583 ( .A(c[14]), .B(c[13]), .Q(n174) );
  NOR31 U584 ( .A(c[15]), .B(c[17]), .C(c[16]), .Q(n175) );
  NOR40 U585 ( .A(n182), .B(c[10]), .C(c[12]), .D(c[11]), .Q(n176) );
  XOR21 U586 ( .A(sin_was_positiveQ), .B(n152), .Q(n217) );
  NAND41 U587 ( .A(n240), .B(n241), .C(n242), .D(n243), .Q(n197) );
  NOR40 U588 ( .A(i[9]), .B(i[8]), .C(i[7]), .D(i[6]), .Q(n243) );
  NOR40 U589 ( .A(i[5]), .B(i[4]), .C(i[19]), .D(i[18]), .Q(n242) );
  NOR40 U590 ( .A(i[17]), .B(i[16]), .C(i[15]), .D(i[14]), .Q(n241) );
  XNR21 U591 ( .A(old_i_data), .B(i_data), .Q(n152) );
  NAND31 U592 ( .A(n257), .B(n290), .C(IorQ), .Q(n169) );
  INV3 U593 ( .A(i_empty), .Q(n290) );
  NOR21 U594 ( .A(i[2]), .B(n270), .Q(n141) );
  XNR21 U595 ( .A(sin_was_positiveI), .B(n152), .Q(n164) );
  NAND22 U596 ( .A(isPositiveI), .B(is9), .Q(n147) );
  NAND31 U597 ( .A(j[2]), .B(n324), .C(n196), .Q(n191) );
  NOR31 U598 ( .A(j[0]), .B(n251), .C(n272), .Q(n196) );
  NAND22 U599 ( .A(is9), .B(n147), .Q(n133) );
  NOR40 U600 ( .A(j[13]), .B(j[12]), .C(j[11]), .D(j[10]), .Q(n245) );
  NOR40 U601 ( .A(i[13]), .B(i[12]), .C(i[11]), .D(i[10]), .Q(n240) );
  NOR40 U602 ( .A(i[12]), .B(i[11]), .C(i[10]), .D(n355), .Q(n409) );
  INV3 U603 ( .A(n404), .Q(n355) );
  OAI311 U604 ( .A(n271), .B(i[2]), .C(n270), .D(n269), .Q(n404) );
  NOR40 U605 ( .A(j[12]), .B(j[11]), .C(j[10]), .D(n325), .Q(n416) );
  INV3 U606 ( .A(n411), .Q(n325) );
  OAI311 U607 ( .A(j[0]), .B(j[2]), .C(n272), .D(n251), .Q(n411) );
  NOR21 U608 ( .A(j[2]), .B(n272), .Q(n215) );
  XOR21 U609 ( .A(sin_was_positiveI), .B(n152), .Q(n143) );
  NOR40 U610 ( .A(i[16]), .B(i[15]), .C(i[14]), .D(i[13]), .Q(n408) );
  NOR40 U611 ( .A(j[16]), .B(j[15]), .C(j[14]), .D(j[13]), .Q(n415) );
  NOR40 U612 ( .A(j[17]), .B(j[16]), .C(j[15]), .D(j[14]), .Q(n246) );
  NAND41 U613 ( .A(n189), .B(n188), .C(\stateQ[0] ), .D(n190), .Q(N1084) );
  NOR21 U614 ( .A(n257), .B(n288), .Q(n190) );
  NOR40 U615 ( .A(i[7]), .B(n380), .C(i[6]), .D(i[5]), .Q(n406) );
  INV3 U616 ( .A(n405), .Q(n380) );
  NOR21 U617 ( .A(i[9]), .B(i[8]), .Q(n405) );
  NOR40 U618 ( .A(j[7]), .B(n349), .C(j[6]), .D(j[5]), .Q(n413) );
  INV3 U619 ( .A(n412), .Q(n349) );
  NOR21 U620 ( .A(j[9]), .B(j[8]), .Q(n412) );
  NAND22 U621 ( .A(is9), .B(isPositiveQ), .Q(n226) );
  NOR40 U622 ( .A(n178), .B(n315), .C(c[19]), .D(c[18]), .Q(n177) );
  INV3 U623 ( .A(n179), .Q(n315) );
  NAND22 U624 ( .A(n180), .B(n181), .Q(n178) );
  NOR31 U625 ( .A(c[1]), .B(c[4]), .C(c[3]), .Q(n179) );
  NAND22 U626 ( .A(is9), .B(n226), .Q(n207) );
  OAI311 U627 ( .A(n322), .B(n292), .C(n319), .D(n199), .Q(N1081) );
  INV3 U628 ( .A(i_data), .Q(n292) );
  INV3 U629 ( .A(n201), .Q(n322) );
  NAND31 U630 ( .A(i_data), .B(n136), .C(n200), .Q(n199) );
  AOI211 U631 ( .A(j[0]), .B(j[2]), .C(n251), .Q(n236) );
  OAI311 U632 ( .A(n191), .B(IorQ), .C(n319), .D(n192), .Q(N1083) );
  NAND31 U633 ( .A(n136), .B(n263), .C(n193), .Q(n192) );
  NOR31 U634 ( .A(c[7]), .B(c[9]), .C(c[8]), .Q(n181) );
  NAND22 U635 ( .A(n321), .B(n203), .Q(n249) );
  INV3 U636 ( .A(n417), .Q(n321) );
  NAND41 U637 ( .A(n416), .B(n415), .C(n414), .D(n413), .Q(n417) );
  NOR40 U638 ( .A(j[4]), .B(j[19]), .C(j[18]), .D(j[17]), .Q(n414) );
  NAND22 U639 ( .A(n352), .B(n136), .Q(n171) );
  INV3 U640 ( .A(n410), .Q(n352) );
  NAND41 U641 ( .A(n409), .B(n408), .C(n407), .D(n406), .Q(n410) );
  NOR40 U642 ( .A(i[4]), .B(i[19]), .C(i[18]), .D(i[17]), .Q(n407) );
  NOR21 U643 ( .A(n279), .B(c[0]), .Q(N503) );
  INV3 U644 ( .A(n244), .Q(n324) );
  NAND41 U645 ( .A(n245), .B(n246), .C(n247), .D(n248), .Q(n244) );
  NOR40 U646 ( .A(j[9]), .B(j[8]), .C(j[7]), .D(j[6]), .Q(n248) );
  NOR40 U647 ( .A(j[5]), .B(j[4]), .C(j[19]), .D(j[18]), .Q(n247) );
  NAND22 U648 ( .A(c[2]), .B(n261), .Q(n182) );
  NAND22 U649 ( .A(reset), .B(n318), .Q(N1073) );
  NAND22 U650 ( .A(n202), .B(reset), .Q(N1080) );
  AOI221 U651 ( .A(n200), .B(n136), .C(n201), .D(n203), .Q(n202) );
  NOR21 U652 ( .A(n275), .B(j[0]), .Q(N1051) );
  NOR21 U653 ( .A(n282), .B(n271), .Q(N768) );
  INV3 U654 ( .A(n395), .Q(n350) );
  NOR21 U655 ( .A(j[18]), .B(j[17]), .Q(n395) );
  INV3 U656 ( .A(n386), .Q(n381) );
  NOR21 U657 ( .A(i[18]), .B(i[17]), .Q(n386) );
  INV3 U658 ( .A(n186), .Q(n317) );
  INV3 U659 ( .A(n183), .Q(n316) );
  NOR31 U660 ( .A(IorQ), .B(i_empty), .C(\stateQ[0] ), .Q(n130) );
  NOR31 U661 ( .A(IorQ), .B(\stateQ[0] ), .C(i_empty), .Q(N1098) );
  NAND22 U662 ( .A(reset), .B(n169), .Q(N563) );
  NOR31 U663 ( .A(n263), .B(\stateI[0] ), .C(i_empty), .Q(N1092) );
  NOR21 U664 ( .A(c[6]), .B(c[5]), .Q(n180) );
  INV3 U665 ( .A(n129), .Q(n291) );
  NAND22 U666 ( .A(n130), .B(isPositiveQ), .Q(n129) );
  NOR21 U667 ( .A(n264), .B(n288), .Q(N499) );
  NOR21 U668 ( .A(n265), .B(n288), .Q(N501) );
  INV3 U669 ( .A(reset), .Q(n288) );
  OAI222 U670 ( .A(n184), .B(n254), .C(my_clk_10M), .D(n254), .Q(n183) );
  OAI222 U671 ( .A(n187), .B(n257), .C(my_clk_10M), .D(n257), .Q(n186) );
endmodule

