
module outFIFO ( inClock, inReset, inReadEnable, inWriteEnable, inData, 
        outWriteCount, outReadCount, outReadError, outWriteError, outFull, 
        outEmpty, outAlmostEmpty, outAlmostFull, outDone, outData );
  output [7:0] outWriteCount;
  output [6:0] outReadCount;
  output [3:0] outData;
  input inClock, inReset, inReadEnable, inWriteEnable, inData;
  output outReadError, outWriteError, outFull, outEmpty, outAlmostEmpty,
         outAlmostFull, outDone;
  wire   N39, N40, N41, N42, N43, N44, N45, sig_fsm_start_R, sig_fsm_start_W,
         N47, N48, N49, N50, sigEnableCounter, N120, N121, N122, N123, N124,
         N125, N126, N128, N129, N130, N131, N132, N136, N137, N138, N139,
         N140, N141, N143, N144, N145, N146, N147, N148, N149, N150, N159,
         N160, N161, N162, N163, N164, N165, N183, N191, N192, N198, N201,
         \FIFO[127][3] , \FIFO[127][2] , \FIFO[127][1] , \FIFO[127][0] ,
         \FIFO[126][3] , \FIFO[126][2] , \FIFO[126][1] , \FIFO[126][0] ,
         \FIFO[125][3] , \FIFO[125][2] , \FIFO[125][1] , \FIFO[125][0] ,
         \FIFO[124][3] , \FIFO[124][2] , \FIFO[124][1] , \FIFO[124][0] ,
         \FIFO[123][3] , \FIFO[123][2] , \FIFO[123][1] , \FIFO[123][0] ,
         \FIFO[122][3] , \FIFO[122][2] , \FIFO[122][1] , \FIFO[122][0] ,
         \FIFO[121][3] , \FIFO[121][2] , \FIFO[121][1] , \FIFO[121][0] ,
         \FIFO[120][3] , \FIFO[120][2] , \FIFO[120][1] , \FIFO[120][0] ,
         \FIFO[119][3] , \FIFO[119][2] , \FIFO[119][1] , \FIFO[119][0] ,
         \FIFO[118][3] , \FIFO[118][2] , \FIFO[118][1] , \FIFO[118][0] ,
         \FIFO[117][3] , \FIFO[117][2] , \FIFO[117][1] , \FIFO[117][0] ,
         \FIFO[116][3] , \FIFO[116][2] , \FIFO[116][1] , \FIFO[116][0] ,
         \FIFO[115][3] , \FIFO[115][2] , \FIFO[115][1] , \FIFO[115][0] ,
         \FIFO[114][3] , \FIFO[114][2] , \FIFO[114][1] , \FIFO[114][0] ,
         \FIFO[113][3] , \FIFO[113][2] , \FIFO[113][1] , \FIFO[113][0] ,
         \FIFO[112][3] , \FIFO[112][2] , \FIFO[112][1] , \FIFO[112][0] ,
         \FIFO[111][3] , \FIFO[111][2] , \FIFO[111][1] , \FIFO[111][0] ,
         \FIFO[110][3] , \FIFO[110][2] , \FIFO[110][1] , \FIFO[110][0] ,
         \FIFO[109][3] , \FIFO[109][2] , \FIFO[109][1] , \FIFO[109][0] ,
         \FIFO[108][3] , \FIFO[108][2] , \FIFO[108][1] , \FIFO[108][0] ,
         \FIFO[107][3] , \FIFO[107][2] , \FIFO[107][1] , \FIFO[107][0] ,
         \FIFO[106][3] , \FIFO[106][2] , \FIFO[106][1] , \FIFO[106][0] ,
         \FIFO[105][3] , \FIFO[105][2] , \FIFO[105][1] , \FIFO[105][0] ,
         \FIFO[104][3] , \FIFO[104][2] , \FIFO[104][1] , \FIFO[104][0] ,
         \FIFO[103][3] , \FIFO[103][2] , \FIFO[103][1] , \FIFO[103][0] ,
         \FIFO[102][3] , \FIFO[102][2] , \FIFO[102][1] , \FIFO[102][0] ,
         \FIFO[101][3] , \FIFO[101][2] , \FIFO[101][1] , \FIFO[101][0] ,
         \FIFO[100][3] , \FIFO[100][2] , \FIFO[100][1] , \FIFO[100][0] ,
         \FIFO[99][3] , \FIFO[99][2] , \FIFO[99][1] , \FIFO[99][0] ,
         \FIFO[98][3] , \FIFO[98][2] , \FIFO[98][1] , \FIFO[98][0] ,
         \FIFO[97][3] , \FIFO[97][2] , \FIFO[97][1] , \FIFO[97][0] ,
         \FIFO[96][3] , \FIFO[96][2] , \FIFO[96][1] , \FIFO[96][0] ,
         \FIFO[95][3] , \FIFO[95][2] , \FIFO[95][1] , \FIFO[95][0] ,
         \FIFO[94][3] , \FIFO[94][2] , \FIFO[94][1] , \FIFO[94][0] ,
         \FIFO[93][3] , \FIFO[93][2] , \FIFO[93][1] , \FIFO[93][0] ,
         \FIFO[92][3] , \FIFO[92][2] , \FIFO[92][1] , \FIFO[92][0] ,
         \FIFO[91][3] , \FIFO[91][2] , \FIFO[91][1] , \FIFO[91][0] ,
         \FIFO[90][3] , \FIFO[90][2] , \FIFO[90][1] , \FIFO[90][0] ,
         \FIFO[89][3] , \FIFO[89][2] , \FIFO[89][1] , \FIFO[89][0] ,
         \FIFO[88][3] , \FIFO[88][2] , \FIFO[88][1] , \FIFO[88][0] ,
         \FIFO[87][3] , \FIFO[87][2] , \FIFO[87][1] , \FIFO[87][0] ,
         \FIFO[86][3] , \FIFO[86][2] , \FIFO[86][1] , \FIFO[86][0] ,
         \FIFO[85][3] , \FIFO[85][2] , \FIFO[85][1] , \FIFO[85][0] ,
         \FIFO[84][3] , \FIFO[84][2] , \FIFO[84][1] , \FIFO[84][0] ,
         \FIFO[83][3] , \FIFO[83][2] , \FIFO[83][1] , \FIFO[83][0] ,
         \FIFO[82][3] , \FIFO[82][2] , \FIFO[82][1] , \FIFO[82][0] ,
         \FIFO[81][3] , \FIFO[81][2] , \FIFO[81][1] , \FIFO[81][0] ,
         \FIFO[80][3] , \FIFO[80][2] , \FIFO[80][1] , \FIFO[80][0] ,
         \FIFO[79][3] , \FIFO[79][2] , \FIFO[79][1] , \FIFO[79][0] ,
         \FIFO[78][3] , \FIFO[78][2] , \FIFO[78][1] , \FIFO[78][0] ,
         \FIFO[77][3] , \FIFO[77][2] , \FIFO[77][1] , \FIFO[77][0] ,
         \FIFO[76][3] , \FIFO[76][2] , \FIFO[76][1] , \FIFO[76][0] ,
         \FIFO[75][3] , \FIFO[75][2] , \FIFO[75][1] , \FIFO[75][0] ,
         \FIFO[74][3] , \FIFO[74][2] , \FIFO[74][1] , \FIFO[74][0] ,
         \FIFO[73][3] , \FIFO[73][2] , \FIFO[73][1] , \FIFO[73][0] ,
         \FIFO[72][3] , \FIFO[72][2] , \FIFO[72][1] , \FIFO[72][0] ,
         \FIFO[71][3] , \FIFO[71][2] , \FIFO[71][1] , \FIFO[71][0] ,
         \FIFO[70][3] , \FIFO[70][2] , \FIFO[70][1] , \FIFO[70][0] ,
         \FIFO[69][3] , \FIFO[69][2] , \FIFO[69][1] , \FIFO[69][0] ,
         \FIFO[68][3] , \FIFO[68][2] , \FIFO[68][1] , \FIFO[68][0] ,
         \FIFO[67][3] , \FIFO[67][2] , \FIFO[67][1] , \FIFO[67][0] ,
         \FIFO[66][3] , \FIFO[66][2] , \FIFO[66][1] , \FIFO[66][0] ,
         \FIFO[65][3] , \FIFO[65][2] , \FIFO[65][1] , \FIFO[65][0] ,
         \FIFO[64][3] , \FIFO[64][2] , \FIFO[64][1] , \FIFO[64][0] ,
         \FIFO[63][3] , \FIFO[63][2] , \FIFO[63][1] , \FIFO[63][0] ,
         \FIFO[62][3] , \FIFO[62][2] , \FIFO[62][1] , \FIFO[62][0] ,
         \FIFO[61][3] , \FIFO[61][2] , \FIFO[61][1] , \FIFO[61][0] ,
         \FIFO[60][3] , \FIFO[60][2] , \FIFO[60][1] , \FIFO[60][0] ,
         \FIFO[59][3] , \FIFO[59][2] , \FIFO[59][1] , \FIFO[59][0] ,
         \FIFO[58][3] , \FIFO[58][2] , \FIFO[58][1] , \FIFO[58][0] ,
         \FIFO[57][3] , \FIFO[57][2] , \FIFO[57][1] , \FIFO[57][0] ,
         \FIFO[56][3] , \FIFO[56][2] , \FIFO[56][1] , \FIFO[56][0] ,
         \FIFO[55][3] , \FIFO[55][2] , \FIFO[55][1] , \FIFO[55][0] ,
         \FIFO[54][3] , \FIFO[54][2] , \FIFO[54][1] , \FIFO[54][0] ,
         \FIFO[53][3] , \FIFO[53][2] , \FIFO[53][1] , \FIFO[53][0] ,
         \FIFO[52][3] , \FIFO[52][2] , \FIFO[52][1] , \FIFO[52][0] ,
         \FIFO[51][3] , \FIFO[51][2] , \FIFO[51][1] , \FIFO[51][0] ,
         \FIFO[50][3] , \FIFO[50][2] , \FIFO[50][1] , \FIFO[50][0] ,
         \FIFO[49][3] , \FIFO[49][2] , \FIFO[49][1] , \FIFO[49][0] ,
         \FIFO[48][3] , \FIFO[48][2] , \FIFO[48][1] , \FIFO[48][0] ,
         \FIFO[47][3] , \FIFO[47][2] , \FIFO[47][1] , \FIFO[47][0] ,
         \FIFO[46][3] , \FIFO[46][2] , \FIFO[46][1] , \FIFO[46][0] ,
         \FIFO[45][3] , \FIFO[45][2] , \FIFO[45][1] , \FIFO[45][0] ,
         \FIFO[44][3] , \FIFO[44][2] , \FIFO[44][1] , \FIFO[44][0] ,
         \FIFO[43][3] , \FIFO[43][2] , \FIFO[43][1] , \FIFO[43][0] ,
         \FIFO[42][3] , \FIFO[42][2] , \FIFO[42][1] , \FIFO[42][0] ,
         \FIFO[41][3] , \FIFO[41][2] , \FIFO[41][1] , \FIFO[41][0] ,
         \FIFO[40][3] , \FIFO[40][2] , \FIFO[40][1] , \FIFO[40][0] ,
         \FIFO[39][3] , \FIFO[39][2] , \FIFO[39][1] , \FIFO[39][0] ,
         \FIFO[38][3] , \FIFO[38][2] , \FIFO[38][1] , \FIFO[38][0] ,
         \FIFO[37][3] , \FIFO[37][2] , \FIFO[37][1] , \FIFO[37][0] ,
         \FIFO[36][3] , \FIFO[36][2] , \FIFO[36][1] , \FIFO[36][0] ,
         \FIFO[35][3] , \FIFO[35][2] , \FIFO[35][1] , \FIFO[35][0] ,
         \FIFO[34][3] , \FIFO[34][2] , \FIFO[34][1] , \FIFO[34][0] ,
         \FIFO[33][3] , \FIFO[33][2] , \FIFO[33][1] , \FIFO[33][0] ,
         \FIFO[32][3] , \FIFO[32][2] , \FIFO[32][1] , \FIFO[32][0] ,
         \FIFO[31][3] , \FIFO[31][2] , \FIFO[31][1] , \FIFO[31][0] ,
         \FIFO[30][3] , \FIFO[30][2] , \FIFO[30][1] , \FIFO[30][0] ,
         \FIFO[29][3] , \FIFO[29][2] , \FIFO[29][1] , \FIFO[29][0] ,
         \FIFO[28][3] , \FIFO[28][2] , \FIFO[28][1] , \FIFO[28][0] ,
         \FIFO[27][3] , \FIFO[27][2] , \FIFO[27][1] , \FIFO[27][0] ,
         \FIFO[26][3] , \FIFO[26][2] , \FIFO[26][1] , \FIFO[26][0] ,
         \FIFO[25][3] , \FIFO[25][2] , \FIFO[25][1] , \FIFO[25][0] ,
         \FIFO[24][3] , \FIFO[24][2] , \FIFO[24][1] , \FIFO[24][0] ,
         \FIFO[23][3] , \FIFO[23][2] , \FIFO[23][1] , \FIFO[23][0] ,
         \FIFO[22][3] , \FIFO[22][2] , \FIFO[22][1] , \FIFO[22][0] ,
         \FIFO[21][3] , \FIFO[21][2] , \FIFO[21][1] , \FIFO[21][0] ,
         \FIFO[20][3] , \FIFO[20][2] , \FIFO[20][1] , \FIFO[20][0] ,
         \FIFO[19][3] , \FIFO[19][2] , \FIFO[19][1] , \FIFO[19][0] ,
         \FIFO[18][3] , \FIFO[18][2] , \FIFO[18][1] , \FIFO[18][0] ,
         \FIFO[17][3] , \FIFO[17][2] , \FIFO[17][1] , \FIFO[17][0] ,
         \FIFO[16][3] , \FIFO[16][2] , \FIFO[16][1] , \FIFO[16][0] ,
         \FIFO[15][3] , \FIFO[15][2] , \FIFO[15][1] , \FIFO[15][0] ,
         \FIFO[14][3] , \FIFO[14][2] , \FIFO[14][1] , \FIFO[14][0] ,
         \FIFO[13][3] , \FIFO[13][2] , \FIFO[13][1] , \FIFO[13][0] ,
         \FIFO[12][3] , \FIFO[12][2] , \FIFO[12][1] , \FIFO[12][0] ,
         \FIFO[11][3] , \FIFO[11][2] , \FIFO[11][1] , \FIFO[11][0] ,
         \FIFO[10][3] , \FIFO[10][2] , \FIFO[10][1] , \FIFO[10][0] ,
         \FIFO[9][3] , \FIFO[9][2] , \FIFO[9][1] , \FIFO[9][0] , \FIFO[8][3] ,
         \FIFO[8][2] , \FIFO[8][1] , \FIFO[8][0] , \FIFO[7][3] , \FIFO[7][2] ,
         \FIFO[7][1] , \FIFO[7][0] , \FIFO[6][3] , \FIFO[6][2] , \FIFO[6][1] ,
         \FIFO[6][0] , \FIFO[5][3] , \FIFO[5][2] , \FIFO[5][1] , \FIFO[5][0] ,
         \FIFO[4][3] , \FIFO[4][2] , \FIFO[4][1] , \FIFO[4][0] , \FIFO[3][3] ,
         \FIFO[3][2] , \FIFO[3][1] , \FIFO[3][0] , \FIFO[2][3] , \FIFO[2][2] ,
         \FIFO[2][1] , \FIFO[2][0] , \FIFO[1][3] , \FIFO[1][2] , \FIFO[1][1] ,
         \FIFO[1][0] , \FIFO[0][3] , \FIFO[0][2] , \FIFO[0][1] , \FIFO[0][0] ,
         N206, N207, N208, N209, N213, N216, N217, N218, N219, N220, N222,
         N223, N224, N225, N226, N227, N228, N918, N1269, N1270, N1276, N1277,
         N1285, N1286, N1287, N1291, N1292, N1293, N1294, N1295, N1296, N1297,
         N1298, N1299, N1300, N1301, N1302, N1303, N1304, N1305, N1306, N1307,
         N1308, N1309, N1310, N1311, N1312, N1313, N1314, N1315, N1316, N1317,
         N1318, N1319, N1320, N1321, N1322, N1323, N1324, N1325, N1326, N1327,
         N1328, N1329, N1330, N1331, N1332, N1333, N1334, N1335, N1336, N1337,
         N1338, N1339, N1340, N1341, N1342, N1343, N1344, N1345, N1346, N1347,
         N1348, N1349, N1350, N1351, N1352, N1353, N1354, N1355, N1356, N1357,
         N1358, N1359, N1360, N1361, N1362, N1363, N1364, N1365, N1366, N1367,
         N1368, N1369, N1370, N1371, N1372, N1373, N1374, N1375, N1376, N1377,
         N1378, N1379, N1380, N1381, N1382, N1383, N1384, N1385, N1386, N1387,
         N1388, N1389, N1390, N1391, N1392, N1393, N1394, N1395, N1396, N1397,
         N1398, N1399, N1400, N1401, N1402, N1403, N1404, N1405, N1406, N1407,
         N1408, N1409, N1410, N1411, N1412, N1413, N1414, N1415, N1416, N1417,
         N1418, N1419, N1420, N1421, N1422, N1423, N1424, N1425, N1426, N1427,
         N1428, N1429, N1430, N1431, N1432, N1433, N1434, N1435, N1436, N1437,
         N1438, N1439, N1440, N1441, N1442, N1443, N1444, N1445, N1446, N1447,
         N1448, N1449, N1450, N1451, N1452, N1453, N1454, N1455, N1456, N1457,
         N1458, N1459, N1460, N1461, N1462, N1463, N1464, N1465, N1466, N1467,
         N1468, N1469, N1470, N1471, N1472, N1473, N1474, N1475, N1476, N1477,
         N1478, N1479, N1480, N1481, N1482, N1483, N1484, N1485, N1486, N1487,
         N1488, N1489, N1490, N1491, N1492, N1493, N1494, N1495, N1496, N1497,
         N1498, N1499, N1500, N1501, N1502, N1503, N1504, N1505, N1506, N1507,
         N1508, N1509, N1510, N1511, N1512, N1513, N1514, N1515, N1516, N1517,
         N1518, N1519, N1520, N1521, N1522, N1523, N1524, N1525, N1526, N1527,
         N1528, N1529, N1530, N1531, N1532, N1533, N1534, N1535, N1536, N1537,
         N1538, N1539, N1540, N1541, N1542, N1543, N1544, N1545, N1546, N1547,
         N1548, N1549, N1550, N1551, N1552, N1553, N1554, N1555, N1556, N1557,
         N1558, N1559, N1560, N1561, N1562, N1563, N1564, N1565, N1566, N1567,
         N1568, N1569, N1570, N1571, N1572, N1573, N1574, N1575, N1576, N1577,
         N1578, N1579, N1580, N1581, N1582, N1583, N1584, N1585, N1586, N1587,
         N1588, N1589, N1590, N1591, N1592, N1593, N1594, N1595, N1596, N1597,
         N1598, N1599, N1600, N1601, N1602, N1603, N1604, N1605, N1606, N1607,
         N1608, N1609, N1610, N1611, N1612, N1613, N1614, N1615, N1616, N1617,
         N1618, N1619, N1620, N1621, N1622, N1623, N1624, N1625, N1626, N1627,
         N1628, N1629, N1630, N1631, N1632, N1633, N1634, N1635, N1636, N1637,
         N1638, N1639, N1640, N1641, N1642, N1643, N1644, N1645, N1646, N1647,
         N1648, N1649, N1650, N1651, N1652, N1653, N1654, N1655, N1656, N1657,
         N1658, N1659, N1660, N1661, N1662, N1663, N1664, N1665, N1666, N1667,
         N1668, N1669, N1670, N1671, N1672, N1673, N1674, N1675, N1676, N1677,
         N1678, N1679, N1680, N1681, N1682, N1683, N1684, N1685, N1686, N1687,
         N1688, N1689, N1690, N1691, N1692, N1693, N1694, N1695, N1696, N1697,
         N1698, N1699, N1700, N1701, N1702, N1703, N1704, N1705, N1706, N1707,
         N1708, N1709, N1710, N1711, N1712, N1713, N1714, N1715, N1716, N1717,
         N1718, N1719, N1720, N1721, N1722, N1723, N1724, N1725, N1726, N1727,
         N1728, N1729, N1730, N1731, N1732, N1733, N1734, N1735, N1736, N1737,
         N1738, N1739, N1740, N1741, N1742, N1743, N1744, N1745, N1746, N1747,
         N1748, N1749, N1750, N1751, N1752, N1753, N1754, N1755, N1756, N1757,
         N1758, N1759, N1760, N1761, N1762, N1763, N1764, N1765, N1766, N1767,
         N1768, N1769, N1770, N1771, N1772, N1773, N1774, N1775, N1776, N1777,
         N1778, N1779, N1780, N1781, N1782, N1783, N1784, N1785, N1786, N1787,
         N1788, N1789, N1790, N1791, N1792, N1793, N1794, N1795, N1796, N1797,
         N1798, N1799, N1800, N1801, N1802, N1804, N1806, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
         n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234,
         n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245,
         n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
         n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
         n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
         n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289,
         n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, \os1/sigQout2 ,
         \os1/sigQout1 , \os1/dff1/n2 , \os2/sigQout2 , \os2/sigQout1 , n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912;
  wire   [3:0] currentState;
  wire   [6:0] i_FIFO;
  wire   [1:0] k_FIFO;
  wire   [6:2] \add_360/carry ;
  wire   [6:2] \add_260/carry ;
  wire   [6:2] \add_256/carry ;
  wire   [7:2] \add_255/carry ;
  wire   [8:0] \r98/carry ;
  assign outFull = N1269;
  assign outEmpty = N1270;
  assign outAlmostEmpty = N1285;

  OAI212 U12 ( .A(n104), .B(n808), .C(n105), .Q(N49) );
  OAI222 U16 ( .A(N1269), .B(n107), .C(n868), .D(n108), .Q(n106) );
  OAI212 U17 ( .A(n109), .B(n808), .C(n831), .Q(N48) );
  OAI212 U23 ( .A(n115), .B(n808), .C(n105), .Q(N47) );
  OAI212 U40 ( .A(n546), .B(n118), .C(n772), .Q(N201) );
  OAI212 U46 ( .A(n661), .B(n631), .C(n798), .Q(N1802) );
  OAI212 U47 ( .A(n124), .B(n126), .C(n789), .Q(N1801) );
  OAI212 U48 ( .A(n124), .B(n127), .C(n790), .Q(N1800) );
  OAI212 U49 ( .A(n124), .B(n128), .C(n790), .Q(N1799) );
  OAI212 U50 ( .A(n632), .B(n659), .C(n790), .Q(N1798) );
  OAI212 U51 ( .A(n126), .B(n659), .C(n790), .Q(N1797) );
  OAI212 U52 ( .A(n127), .B(n659), .C(n790), .Q(N1796) );
  OAI212 U53 ( .A(n128), .B(n659), .C(n790), .Q(N1795) );
  OAI212 U54 ( .A(n632), .B(n657), .C(n790), .Q(N1794) );
  OAI212 U55 ( .A(n126), .B(n657), .C(n790), .Q(N1793) );
  OAI212 U56 ( .A(n127), .B(n657), .C(n790), .Q(N1792) );
  OAI212 U57 ( .A(n128), .B(n657), .C(n790), .Q(N1791) );
  OAI212 U58 ( .A(n632), .B(n655), .C(n790), .Q(N1790) );
  OAI212 U59 ( .A(n126), .B(n655), .C(n791), .Q(N1789) );
  OAI212 U60 ( .A(n127), .B(n655), .C(n791), .Q(N1788) );
  OAI212 U61 ( .A(n128), .B(n655), .C(n791), .Q(N1787) );
  OAI212 U62 ( .A(n632), .B(n653), .C(n791), .Q(N1786) );
  OAI212 U63 ( .A(n126), .B(n653), .C(n791), .Q(N1785) );
  OAI212 U64 ( .A(n127), .B(n653), .C(n791), .Q(N1784) );
  OAI212 U65 ( .A(n128), .B(n653), .C(n791), .Q(N1783) );
  OAI212 U66 ( .A(n632), .B(n651), .C(n791), .Q(N1782) );
  OAI212 U67 ( .A(n126), .B(n651), .C(n791), .Q(N1781) );
  OAI212 U68 ( .A(n127), .B(n651), .C(n791), .Q(N1780) );
  OAI212 U69 ( .A(n128), .B(n651), .C(n791), .Q(N1779) );
  OAI212 U70 ( .A(n632), .B(n649), .C(n792), .Q(N1778) );
  OAI212 U71 ( .A(n126), .B(n649), .C(n792), .Q(N1777) );
  OAI212 U72 ( .A(n127), .B(n649), .C(n792), .Q(N1776) );
  OAI212 U73 ( .A(n128), .B(n649), .C(n792), .Q(N1775) );
  OAI212 U74 ( .A(n632), .B(n647), .C(n792), .Q(N1774) );
  OAI212 U75 ( .A(n126), .B(n647), .C(n792), .Q(N1773) );
  OAI212 U76 ( .A(n127), .B(n647), .C(n792), .Q(N1772) );
  OAI212 U77 ( .A(n128), .B(n647), .C(n792), .Q(N1771) );
  OAI212 U78 ( .A(n632), .B(n645), .C(n792), .Q(N1770) );
  OAI212 U79 ( .A(n126), .B(n645), .C(n792), .Q(N1769) );
  OAI212 U80 ( .A(n127), .B(n645), .C(n792), .Q(N1768) );
  OAI212 U81 ( .A(n128), .B(n645), .C(n793), .Q(N1767) );
  OAI212 U82 ( .A(n631), .B(n643), .C(n793), .Q(N1766) );
  OAI212 U83 ( .A(n126), .B(n643), .C(n793), .Q(N1765) );
  OAI212 U84 ( .A(n127), .B(n643), .C(n793), .Q(N1764) );
  OAI212 U85 ( .A(n128), .B(n643), .C(n793), .Q(N1763) );
  OAI212 U86 ( .A(n631), .B(n641), .C(n793), .Q(N1762) );
  OAI212 U87 ( .A(n126), .B(n641), .C(n793), .Q(N1761) );
  OAI212 U88 ( .A(n127), .B(n641), .C(n793), .Q(N1760) );
  OAI212 U89 ( .A(n128), .B(n641), .C(n793), .Q(N1759) );
  OAI212 U90 ( .A(n631), .B(n595), .C(n793), .Q(N1758) );
  OAI212 U91 ( .A(n126), .B(n139), .C(n793), .Q(N1757) );
  OAI212 U92 ( .A(n127), .B(n595), .C(n794), .Q(N1756) );
  OAI212 U93 ( .A(n128), .B(n139), .C(n794), .Q(N1755) );
  OAI212 U94 ( .A(n631), .B(n594), .C(n794), .Q(N1754) );
  OAI212 U95 ( .A(n126), .B(n140), .C(n794), .Q(N1753) );
  OAI212 U96 ( .A(n127), .B(n594), .C(n794), .Q(N1752) );
  OAI212 U97 ( .A(n128), .B(n140), .C(n794), .Q(N1751) );
  OAI212 U98 ( .A(n631), .B(n593), .C(n794), .Q(N1750) );
  OAI212 U99 ( .A(n126), .B(n141), .C(n794), .Q(N1749) );
  OAI212 U100 ( .A(n127), .B(n593), .C(n794), .Q(N1748) );
  OAI212 U101 ( .A(n128), .B(n141), .C(n794), .Q(N1747) );
  OAI212 U102 ( .A(n631), .B(n142), .C(n794), .Q(N1746) );
  OAI212 U103 ( .A(n126), .B(n592), .C(n795), .Q(N1745) );
  OAI212 U104 ( .A(n127), .B(n591), .C(n795), .Q(N1744) );
  OAI212 U105 ( .A(n128), .B(n142), .C(n795), .Q(N1743) );
  OAI212 U106 ( .A(n631), .B(n143), .C(n795), .Q(N1742) );
  OAI212 U108 ( .A(n126), .B(n586), .C(n795), .Q(N1741) );
  OAI212 U110 ( .A(n127), .B(n585), .C(n795), .Q(N1740) );
  OAI212 U113 ( .A(n128), .B(n143), .C(n795), .Q(N1739) );
  OAI212 U116 ( .A(n124), .B(n630), .C(n795), .Q(N1738) );
  OAI212 U117 ( .A(n124), .B(n628), .C(n795), .Q(N1737) );
  OAI212 U118 ( .A(n124), .B(n626), .C(n795), .Q(N1736) );
  OAI212 U119 ( .A(n124), .B(n624), .C(n795), .Q(N1735) );
  OAI212 U120 ( .A(n659), .B(n630), .C(n796), .Q(N1734) );
  OAI212 U121 ( .A(n659), .B(n628), .C(n796), .Q(N1733) );
  OAI212 U122 ( .A(n659), .B(n626), .C(n796), .Q(N1732) );
  OAI212 U123 ( .A(n659), .B(n624), .C(n796), .Q(N1731) );
  OAI212 U124 ( .A(n657), .B(n630), .C(n796), .Q(N1730) );
  OAI212 U126 ( .A(n657), .B(n628), .C(n796), .Q(N1729) );
  OAI212 U127 ( .A(n657), .B(n626), .C(n796), .Q(N1728) );
  OAI212 U128 ( .A(n657), .B(n624), .C(n796), .Q(N1727) );
  OAI212 U129 ( .A(n655), .B(n630), .C(n796), .Q(N1726) );
  OAI212 U130 ( .A(n655), .B(n628), .C(n796), .Q(N1725) );
  OAI212 U131 ( .A(n655), .B(n626), .C(n796), .Q(N1724) );
  OAI212 U132 ( .A(n655), .B(n624), .C(n797), .Q(N1723) );
  OAI212 U133 ( .A(n653), .B(n630), .C(n797), .Q(N1722) );
  OAI212 U134 ( .A(n653), .B(n628), .C(n797), .Q(N1721) );
  OAI212 U135 ( .A(n653), .B(n626), .C(n797), .Q(N1720) );
  OAI212 U137 ( .A(n653), .B(n624), .C(n797), .Q(N1719) );
  OAI212 U138 ( .A(n651), .B(n630), .C(n797), .Q(N1718) );
  OAI212 U139 ( .A(n651), .B(n628), .C(n797), .Q(N1717) );
  OAI212 U140 ( .A(n651), .B(n626), .C(n797), .Q(N1716) );
  OAI212 U141 ( .A(n651), .B(n624), .C(n797), .Q(N1715) );
  OAI212 U142 ( .A(n649), .B(n630), .C(n797), .Q(N1714) );
  OAI212 U143 ( .A(n649), .B(n628), .C(n797), .Q(N1713) );
  OAI212 U144 ( .A(n649), .B(n626), .C(n798), .Q(N1712) );
  OAI212 U145 ( .A(n649), .B(n624), .C(n798), .Q(N1711) );
  OAI212 U146 ( .A(n647), .B(n630), .C(n798), .Q(N1710) );
  OAI212 U148 ( .A(n647), .B(n628), .C(n798), .Q(N1709) );
  OAI212 U149 ( .A(n647), .B(n626), .C(n798), .Q(N1708) );
  OAI212 U150 ( .A(n647), .B(n624), .C(n798), .Q(N1707) );
  OAI212 U151 ( .A(n645), .B(n629), .C(n798), .Q(N1706) );
  OAI212 U152 ( .A(n645), .B(n627), .C(n798), .Q(N1705) );
  OAI212 U153 ( .A(n645), .B(n625), .C(n798), .Q(N1704) );
  OAI212 U154 ( .A(n645), .B(n623), .C(n798), .Q(N1703) );
  OAI212 U155 ( .A(n643), .B(n629), .C(n799), .Q(N1702) );
  OAI212 U156 ( .A(n643), .B(n627), .C(n799), .Q(N1701) );
  OAI212 U157 ( .A(n643), .B(n625), .C(n799), .Q(N1700) );
  OAI212 U159 ( .A(n643), .B(n623), .C(n799), .Q(N1699) );
  OAI212 U160 ( .A(n641), .B(n629), .C(n799), .Q(N1698) );
  OAI212 U161 ( .A(n641), .B(n627), .C(n799), .Q(N1697) );
  OAI212 U162 ( .A(n641), .B(n625), .C(n799), .Q(N1696) );
  OAI212 U163 ( .A(n641), .B(n623), .C(n799), .Q(N1695) );
  OAI212 U164 ( .A(n595), .B(n629), .C(n799), .Q(N1694) );
  OAI212 U165 ( .A(n139), .B(n627), .C(n799), .Q(N1693) );
  OAI212 U166 ( .A(n595), .B(n625), .C(n799), .Q(N1692) );
  OAI212 U167 ( .A(n139), .B(n623), .C(n800), .Q(N1691) );
  OAI212 U168 ( .A(n594), .B(n629), .C(n800), .Q(N1690) );
  OAI212 U170 ( .A(n140), .B(n627), .C(n800), .Q(N1689) );
  OAI212 U171 ( .A(n594), .B(n625), .C(n800), .Q(N1688) );
  OAI212 U172 ( .A(n140), .B(n623), .C(n800), .Q(N1687) );
  OAI212 U173 ( .A(n593), .B(n629), .C(n800), .Q(N1686) );
  OAI212 U174 ( .A(n141), .B(n627), .C(n800), .Q(N1685) );
  OAI212 U175 ( .A(n593), .B(n625), .C(n800), .Q(N1684) );
  OAI212 U176 ( .A(n141), .B(n623), .C(n800), .Q(N1683) );
  OAI212 U177 ( .A(n592), .B(n629), .C(n800), .Q(N1682) );
  OAI212 U178 ( .A(n591), .B(n627), .C(n800), .Q(N1681) );
  OAI212 U179 ( .A(n142), .B(n625), .C(n801), .Q(N1680) );
  OAI212 U181 ( .A(n592), .B(n623), .C(n801), .Q(N1679) );
  OAI212 U182 ( .A(n586), .B(n629), .C(n801), .Q(N1678) );
  OAI212 U184 ( .A(n585), .B(n627), .C(n801), .Q(N1677) );
  OAI212 U186 ( .A(n143), .B(n625), .C(n801), .Q(N1676) );
  OAI212 U188 ( .A(n586), .B(n623), .C(n801), .Q(N1675) );
  OAI212 U191 ( .A(n124), .B(n622), .C(n801), .Q(N1674) );
  OAI212 U192 ( .A(n124), .B(n619), .C(n801), .Q(N1673) );
  OAI212 U193 ( .A(n661), .B(n617), .C(n801), .Q(N1672) );
  OAI212 U194 ( .A(n661), .B(n615), .C(n801), .Q(N1671) );
  OAI212 U195 ( .A(n659), .B(n622), .C(n801), .Q(N1670) );
  OAI212 U197 ( .A(n659), .B(n620), .C(n802), .Q(N1669) );
  OAI212 U198 ( .A(n659), .B(n617), .C(n802), .Q(N1668) );
  OAI212 U199 ( .A(n659), .B(n615), .C(n802), .Q(N1667) );
  OAI212 U200 ( .A(n657), .B(n622), .C(n802), .Q(N1666) );
  OAI212 U201 ( .A(n657), .B(n619), .C(n802), .Q(N1665) );
  OAI212 U202 ( .A(n657), .B(n617), .C(n802), .Q(N1664) );
  OAI212 U203 ( .A(n657), .B(n615), .C(n802), .Q(N1663) );
  OAI212 U204 ( .A(n655), .B(n622), .C(n802), .Q(N1662) );
  OAI212 U205 ( .A(n655), .B(n620), .C(n802), .Q(N1661) );
  OAI212 U206 ( .A(n655), .B(n617), .C(n802), .Q(N1660) );
  OAI212 U207 ( .A(n655), .B(n615), .C(n802), .Q(N1659) );
  OAI212 U208 ( .A(n653), .B(n622), .C(n803), .Q(N1658) );
  OAI212 U209 ( .A(n653), .B(n619), .C(n803), .Q(N1657) );
  OAI212 U210 ( .A(n653), .B(n617), .C(n803), .Q(N1656) );
  OAI212 U211 ( .A(n653), .B(n615), .C(n803), .Q(N1655) );
  OAI212 U212 ( .A(n651), .B(n622), .C(n803), .Q(N1654) );
  OAI212 U213 ( .A(n651), .B(n620), .C(n803), .Q(N1653) );
  OAI212 U214 ( .A(n651), .B(n617), .C(n803), .Q(N1652) );
  OAI212 U215 ( .A(n651), .B(n615), .C(n803), .Q(N1651) );
  OAI212 U216 ( .A(n649), .B(n622), .C(n803), .Q(N1650) );
  OAI212 U218 ( .A(n649), .B(n619), .C(n803), .Q(N1649) );
  OAI212 U219 ( .A(n649), .B(n617), .C(n803), .Q(N1648) );
  OAI212 U220 ( .A(n649), .B(n615), .C(n804), .Q(N1647) );
  OAI212 U221 ( .A(n647), .B(n622), .C(n804), .Q(N1646) );
  OAI212 U222 ( .A(n647), .B(n620), .C(n804), .Q(N1645) );
  OAI212 U223 ( .A(n647), .B(n617), .C(n804), .Q(N1644) );
  OAI212 U224 ( .A(n647), .B(n615), .C(n804), .Q(N1643) );
  OAI212 U225 ( .A(n645), .B(n621), .C(n804), .Q(N1642) );
  OAI212 U226 ( .A(n645), .B(n619), .C(n804), .Q(N1641) );
  OAI212 U227 ( .A(n645), .B(n616), .C(n804), .Q(N1640) );
  OAI212 U229 ( .A(n645), .B(n614), .C(n804), .Q(N1639) );
  OAI212 U230 ( .A(n643), .B(n621), .C(n804), .Q(N1638) );
  OAI212 U231 ( .A(n643), .B(n620), .C(n804), .Q(N1637) );
  OAI212 U232 ( .A(n643), .B(n616), .C(n805), .Q(N1636) );
  OAI212 U233 ( .A(n643), .B(n614), .C(n805), .Q(N1635) );
  OAI212 U234 ( .A(n641), .B(n621), .C(n805), .Q(N1634) );
  OAI212 U235 ( .A(n641), .B(n618), .C(n805), .Q(N1633) );
  OAI212 U236 ( .A(n641), .B(n616), .C(n805), .Q(N1632) );
  OAI212 U237 ( .A(n641), .B(n614), .C(n805), .Q(N1631) );
  OAI212 U238 ( .A(n595), .B(n621), .C(n805), .Q(N1630) );
  OAI212 U240 ( .A(n139), .B(n618), .C(n805), .Q(N1629) );
  OAI212 U241 ( .A(n595), .B(n616), .C(n805), .Q(N1628) );
  OAI212 U242 ( .A(n139), .B(n614), .C(n805), .Q(N1627) );
  OAI212 U243 ( .A(n594), .B(n621), .C(n805), .Q(N1626) );
  OAI212 U244 ( .A(n140), .B(n618), .C(n806), .Q(N1625) );
  OAI212 U245 ( .A(n594), .B(n616), .C(n806), .Q(N1624) );
  OAI212 U246 ( .A(n140), .B(n614), .C(n806), .Q(N1623) );
  OAI212 U247 ( .A(n593), .B(n621), .C(n806), .Q(N1622) );
  OAI212 U248 ( .A(n141), .B(n618), .C(n806), .Q(N1621) );
  OAI212 U249 ( .A(n593), .B(n616), .C(n806), .Q(N1620) );
  OAI212 U251 ( .A(n141), .B(n614), .C(n806), .Q(N1619) );
  OAI212 U252 ( .A(n591), .B(n621), .C(n806), .Q(N1618) );
  OAI212 U253 ( .A(n142), .B(n618), .C(n782), .Q(N1617) );
  OAI212 U254 ( .A(n592), .B(n616), .C(n782), .Q(N1616) );
  OAI212 U255 ( .A(n591), .B(n614), .C(n781), .Q(N1615) );
  OAI212 U256 ( .A(n585), .B(n621), .C(n781), .Q(N1614) );
  OAI212 U258 ( .A(n143), .B(n618), .C(n781), .Q(N1613) );
  OAI212 U260 ( .A(n586), .B(n616), .C(n781), .Q(N1612) );
  OAI212 U262 ( .A(n585), .B(n614), .C(n781), .Q(N1611) );
  OAI212 U265 ( .A(n661), .B(n613), .C(n781), .Q(N1610) );
  OAI212 U267 ( .A(n661), .B(n610), .C(n781), .Q(N1609) );
  OAI212 U268 ( .A(n661), .B(n607), .C(n781), .Q(N1608) );
  OAI212 U269 ( .A(n661), .B(n605), .C(n781), .Q(N1607) );
  OAI212 U270 ( .A(n659), .B(n613), .C(n781), .Q(N1606) );
  OAI212 U271 ( .A(n129), .B(n611), .C(n781), .Q(N1605) );
  OAI212 U272 ( .A(n129), .B(n608), .C(n780), .Q(N1604) );
  OAI212 U273 ( .A(n129), .B(n605), .C(n780), .Q(N1603) );
  OAI212 U274 ( .A(n657), .B(n613), .C(n780), .Q(N1602) );
  OAI212 U275 ( .A(n130), .B(n610), .C(n780), .Q(N1601) );
  OAI212 U276 ( .A(n130), .B(n607), .C(n780), .Q(N1600) );
  OAI212 U278 ( .A(n130), .B(n605), .C(n780), .Q(N1599) );
  OAI212 U279 ( .A(n655), .B(n613), .C(n780), .Q(N1598) );
  OAI212 U280 ( .A(n131), .B(n611), .C(n780), .Q(N1597) );
  OAI212 U281 ( .A(n131), .B(n608), .C(n780), .Q(N1596) );
  OAI212 U282 ( .A(n131), .B(n605), .C(n780), .Q(N1595) );
  OAI212 U283 ( .A(n653), .B(n613), .C(n780), .Q(N1594) );
  OAI212 U284 ( .A(n132), .B(n610), .C(n779), .Q(N1593) );
  OAI212 U285 ( .A(n132), .B(n607), .C(n779), .Q(N1592) );
  OAI212 U286 ( .A(n132), .B(n605), .C(n779), .Q(N1591) );
  OAI212 U287 ( .A(n651), .B(n613), .C(n779), .Q(N1590) );
  OAI212 U289 ( .A(n133), .B(n611), .C(n779), .Q(N1589) );
  OAI212 U290 ( .A(n133), .B(n608), .C(n779), .Q(N1588) );
  OAI212 U291 ( .A(n133), .B(n605), .C(n779), .Q(N1587) );
  OAI212 U292 ( .A(n649), .B(n613), .C(n779), .Q(N1586) );
  OAI212 U293 ( .A(n134), .B(n610), .C(n779), .Q(N1585) );
  OAI212 U294 ( .A(n134), .B(n607), .C(n779), .Q(N1584) );
  OAI212 U295 ( .A(n134), .B(n605), .C(n779), .Q(N1583) );
  OAI212 U296 ( .A(n647), .B(n613), .C(n778), .Q(N1582) );
  OAI212 U297 ( .A(n135), .B(n611), .C(n778), .Q(N1581) );
  OAI212 U298 ( .A(n135), .B(n608), .C(n778), .Q(N1580) );
  OAI212 U300 ( .A(n135), .B(n605), .C(n778), .Q(N1579) );
  OAI212 U301 ( .A(n645), .B(n612), .C(n778), .Q(N1578) );
  OAI212 U302 ( .A(n136), .B(n610), .C(n778), .Q(N1577) );
  OAI212 U303 ( .A(n136), .B(n607), .C(n778), .Q(N1576) );
  OAI212 U304 ( .A(n136), .B(n604), .C(n778), .Q(N1575) );
  OAI212 U305 ( .A(n643), .B(n612), .C(n778), .Q(N1574) );
  OAI212 U306 ( .A(n137), .B(n611), .C(n778), .Q(N1573) );
  OAI212 U307 ( .A(n137), .B(n608), .C(n777), .Q(N1572) );
  OAI212 U308 ( .A(n137), .B(n604), .C(n777), .Q(N1571) );
  OAI212 U309 ( .A(n641), .B(n612), .C(n777), .Q(N1570) );
  OAI212 U311 ( .A(n138), .B(n609), .C(n777), .Q(N1569) );
  OAI212 U312 ( .A(n138), .B(n606), .C(n777), .Q(N1568) );
  OAI212 U313 ( .A(n138), .B(n604), .C(n777), .Q(N1567) );
  OAI212 U314 ( .A(n595), .B(n612), .C(n777), .Q(N1566) );
  OAI212 U315 ( .A(n139), .B(n609), .C(n777), .Q(N1565) );
  OAI212 U316 ( .A(n595), .B(n606), .C(n777), .Q(N1564) );
  OAI212 U317 ( .A(n139), .B(n604), .C(n777), .Q(N1563) );
  OAI212 U318 ( .A(n594), .B(n612), .C(n777), .Q(N1562) );
  OAI212 U319 ( .A(n140), .B(n609), .C(n776), .Q(N1561) );
  OAI212 U320 ( .A(n594), .B(n606), .C(n776), .Q(N1560) );
  OAI212 U322 ( .A(n140), .B(n604), .C(n776), .Q(N1559) );
  OAI212 U323 ( .A(n593), .B(n612), .C(n776), .Q(N1558) );
  OAI212 U324 ( .A(n141), .B(n609), .C(n776), .Q(N1557) );
  OAI212 U325 ( .A(n593), .B(n606), .C(n776), .Q(N1556) );
  OAI212 U326 ( .A(n141), .B(n604), .C(n776), .Q(N1555) );
  OAI212 U327 ( .A(n142), .B(n612), .C(n776), .Q(N1554) );
  OAI212 U328 ( .A(n592), .B(n609), .C(n776), .Q(N1553) );
  OAI212 U329 ( .A(n591), .B(n606), .C(n776), .Q(N1552) );
  OAI212 U330 ( .A(n142), .B(n604), .C(n776), .Q(N1551) );
  OAI212 U331 ( .A(n143), .B(n612), .C(n775), .Q(N1550) );
  OAI212 U334 ( .A(n586), .B(n609), .C(n775), .Q(N1549) );
  OAI212 U336 ( .A(n585), .B(n606), .C(n775), .Q(N1548) );
  OAI212 U338 ( .A(n143), .B(n604), .C(n775), .Q(N1547) );
  OAI212 U341 ( .A(n661), .B(n603), .C(n775), .Q(N1546) );
  OAI212 U342 ( .A(n661), .B(n178), .C(n775), .Q(N1545) );
  OAI212 U343 ( .A(n661), .B(n179), .C(n775), .Q(N1544) );
  OAI212 U344 ( .A(n661), .B(n180), .C(n775), .Q(N1543) );
  OAI212 U345 ( .A(n129), .B(n603), .C(n775), .Q(N1542) );
  OAI212 U346 ( .A(n129), .B(n178), .C(n775), .Q(N1541) );
  OAI212 U347 ( .A(n129), .B(n179), .C(n774), .Q(N1540) );
  OAI212 U349 ( .A(n129), .B(n180), .C(n775), .Q(N1539) );
  OAI212 U350 ( .A(n130), .B(n603), .C(n774), .Q(N1538) );
  OAI212 U351 ( .A(n130), .B(n178), .C(n774), .Q(N1537) );
  OAI212 U352 ( .A(n130), .B(n179), .C(n774), .Q(N1536) );
  OAI212 U353 ( .A(n130), .B(n180), .C(n774), .Q(N1535) );
  OAI212 U354 ( .A(n131), .B(n603), .C(n774), .Q(N1534) );
  OAI212 U355 ( .A(n131), .B(n178), .C(n778), .Q(N1533) );
  OAI212 U356 ( .A(n131), .B(n179), .C(n782), .Q(N1532) );
  OAI212 U357 ( .A(n131), .B(n180), .C(n782), .Q(N1531) );
  OAI212 U358 ( .A(n132), .B(n603), .C(n782), .Q(N1530) );
  OAI212 U360 ( .A(n132), .B(n178), .C(n782), .Q(N1529) );
  OAI212 U361 ( .A(n132), .B(n179), .C(n782), .Q(N1528) );
  OAI212 U362 ( .A(n132), .B(n180), .C(n782), .Q(N1527) );
  OAI212 U363 ( .A(n133), .B(n603), .C(n782), .Q(N1526) );
  OAI212 U364 ( .A(n133), .B(n178), .C(n782), .Q(N1525) );
  OAI212 U365 ( .A(n133), .B(n179), .C(n789), .Q(N1524) );
  OAI212 U366 ( .A(n133), .B(n180), .C(n782), .Q(N1523) );
  OAI212 U367 ( .A(n134), .B(n603), .C(n783), .Q(N1522) );
  OAI212 U368 ( .A(n134), .B(n178), .C(n783), .Q(N1521) );
  OAI212 U369 ( .A(n134), .B(n179), .C(n783), .Q(N1520) );
  OAI212 U371 ( .A(n134), .B(n180), .C(n783), .Q(N1519) );
  OAI212 U372 ( .A(n135), .B(n603), .C(n783), .Q(N1518) );
  OAI212 U373 ( .A(n135), .B(n178), .C(n783), .Q(N1517) );
  OAI212 U374 ( .A(n135), .B(n179), .C(n783), .Q(N1516) );
  OAI212 U375 ( .A(n135), .B(n180), .C(n783), .Q(N1515) );
  OAI212 U376 ( .A(n136), .B(n602), .C(n783), .Q(N1514) );
  OAI212 U377 ( .A(n136), .B(n178), .C(n783), .Q(N1513) );
  OAI212 U378 ( .A(n136), .B(n179), .C(n783), .Q(N1512) );
  OAI212 U379 ( .A(n136), .B(n180), .C(n784), .Q(N1511) );
  OAI212 U380 ( .A(n137), .B(n602), .C(n784), .Q(N1510) );
  OAI212 U381 ( .A(n137), .B(n178), .C(n784), .Q(N1509) );
  OAI212 U382 ( .A(n137), .B(n179), .C(n784), .Q(N1508) );
  OAI212 U383 ( .A(n137), .B(n180), .C(n784), .Q(N1507) );
  OAI212 U384 ( .A(n138), .B(n602), .C(n784), .Q(N1506) );
  OAI212 U385 ( .A(n138), .B(n178), .C(n784), .Q(N1505) );
  OAI212 U386 ( .A(n138), .B(n179), .C(n784), .Q(N1504) );
  OAI212 U387 ( .A(n138), .B(n180), .C(n784), .Q(N1503) );
  OAI212 U390 ( .A(n595), .B(n602), .C(n784), .Q(N1502) );
  OAI212 U391 ( .A(n139), .B(n178), .C(n784), .Q(N1501) );
  OAI212 U394 ( .A(n595), .B(n179), .C(n785), .Q(N1500) );
  OAI212 U399 ( .A(n594), .B(n602), .C(n785), .Q(N1498) );
  OAI212 U406 ( .A(n593), .B(n602), .C(n785), .Q(N1494) );
  OAI212 U413 ( .A(n592), .B(n602), .C(n785), .Q(N1490) );
  OAI212 U420 ( .A(n586), .B(n602), .C(n785), .Q(N1486) );
  OAI212 U432 ( .A(n661), .B(n601), .C(n785), .Q(N1482) );
  OAI212 U439 ( .A(n129), .B(n601), .C(n785), .Q(N1478) );
  OAI212 U446 ( .A(n130), .B(n601), .C(n785), .Q(N1474) );
  OAI212 U453 ( .A(n131), .B(n601), .C(n785), .Q(N1470) );
  OAI212 U460 ( .A(n132), .B(n601), .C(n785), .Q(N1466) );
  OAI212 U467 ( .A(n133), .B(n601), .C(n785), .Q(N1462) );
  OAI212 U474 ( .A(n134), .B(n601), .C(n786), .Q(N1458) );
  OAI212 U481 ( .A(n135), .B(n601), .C(n786), .Q(N1454) );
  OAI212 U488 ( .A(n136), .B(n600), .C(n786), .Q(N1450) );
  OAI212 U495 ( .A(n137), .B(n600), .C(n786), .Q(N1446) );
  OAI212 U502 ( .A(n138), .B(n600), .C(n786), .Q(N1442) );
  OAI212 U509 ( .A(n139), .B(n600), .C(n786), .Q(N1438) );
  OAI212 U516 ( .A(n140), .B(n600), .C(n786), .Q(N1434) );
  OAI212 U523 ( .A(n141), .B(n600), .C(n786), .Q(N1430) );
  OAI212 U530 ( .A(n591), .B(n600), .C(n786), .Q(N1426) );
  OAI212 U537 ( .A(n585), .B(n600), .C(n786), .Q(N1422) );
  OAI212 U549 ( .A(n661), .B(n597), .C(n786), .Q(N1418) );
  OAI212 U556 ( .A(n659), .B(n597), .C(n787), .Q(N1414) );
  OAI212 U563 ( .A(n130), .B(n597), .C(n787), .Q(N1410) );
  OAI212 U570 ( .A(n655), .B(n597), .C(n787), .Q(N1406) );
  OAI212 U577 ( .A(n132), .B(n597), .C(n787), .Q(N1402) );
  OAI212 U584 ( .A(n133), .B(n597), .C(n787), .Q(N1398) );
  OAI212 U591 ( .A(n134), .B(n597), .C(n787), .Q(N1394) );
  OAI212 U598 ( .A(n135), .B(n597), .C(n787), .Q(N1390) );
  OAI212 U605 ( .A(n136), .B(n596), .C(n787), .Q(N1386) );
  OAI212 U612 ( .A(n137), .B(n596), .C(n787), .Q(N1382) );
  OAI212 U619 ( .A(n138), .B(n596), .C(n787), .Q(N1378) );
  OAI212 U626 ( .A(n595), .B(n596), .C(n787), .Q(N1374) );
  OAI212 U633 ( .A(n594), .B(n596), .C(n788), .Q(N1370) );
  OAI212 U640 ( .A(n593), .B(n596), .C(n788), .Q(N1366) );
  OAI212 U647 ( .A(n592), .B(n596), .C(n788), .Q(N1362) );
  OAI212 U654 ( .A(n586), .B(n596), .C(n788), .Q(N1358) );
  OAI212 U666 ( .A(n661), .B(n590), .C(n788), .Q(N1354) );
  OAI212 U674 ( .A(n659), .B(n590), .C(n788), .Q(N1350) );
  OAI212 U682 ( .A(n657), .B(n590), .C(n788), .Q(N1346) );
  OAI212 U690 ( .A(n655), .B(n590), .C(n788), .Q(N1342) );
  OAI212 U699 ( .A(n653), .B(n590), .C(n788), .Q(N1338) );
  OAI212 U707 ( .A(n651), .B(n590), .C(n788), .Q(N1334) );
  OAI212 U715 ( .A(n649), .B(n590), .C(n788), .Q(N1330) );
  OAI212 U723 ( .A(n647), .B(n590), .C(n789), .Q(N1326) );
  OAI212 U732 ( .A(n645), .B(n589), .C(n789), .Q(N1322) );
  OAI212 U740 ( .A(n643), .B(n589), .C(n789), .Q(N1318) );
  OAI212 U748 ( .A(n641), .B(n589), .C(n789), .Q(N1314) );
  OAI212 U756 ( .A(n595), .B(n589), .C(n789), .Q(N1310) );
  OAI212 U765 ( .A(n594), .B(n589), .C(n789), .Q(N1306) );
  OAI212 U774 ( .A(n593), .B(n589), .C(n789), .Q(N1302) );
  OAI212 U783 ( .A(n591), .B(n589), .C(n789), .Q(N1298) );
  OAI212 U792 ( .A(n585), .B(n589), .C(n789), .Q(N1294) );
  ADD22 \add_360/U1_1_1  ( .A(n582), .B(n824), .CO(\add_360/carry [2]), .S(
        N216) );
  ADD22 \add_360/U1_1_2  ( .A(n581), .B(\add_360/carry [2]), .CO(
        \add_360/carry [3]), .S(N217) );
  ADD22 \add_360/U1_1_3  ( .A(n814), .B(\add_360/carry [3]), .CO(
        \add_360/carry [4]), .S(N218) );
  ADD22 \add_360/U1_1_4  ( .A(n580), .B(\add_360/carry [4]), .CO(
        \add_360/carry [5]), .S(N219) );
  ADD22 \add_360/U1_1_5  ( .A(n579), .B(\add_360/carry [5]), .CO(
        \add_360/carry [6]), .S(N220) );
  ADD22 \add_260/U1_1_1  ( .A(outReadCount[1]), .B(outReadCount[0]), .CO(
        \add_260/carry [2]), .S(N136) );
  ADD22 \add_260/U1_1_2  ( .A(outReadCount[2]), .B(\add_260/carry [2]), .CO(
        \add_260/carry [3]), .S(N137) );
  ADD22 \add_260/U1_1_3  ( .A(outReadCount[3]), .B(\add_260/carry [3]), .CO(
        \add_260/carry [4]), .S(N138) );
  ADD22 \add_260/U1_1_4  ( .A(outReadCount[4]), .B(\add_260/carry [4]), .CO(
        \add_260/carry [5]), .S(N139) );
  ADD22 \add_260/U1_1_5  ( .A(outReadCount[5]), .B(\add_260/carry [5]), .CO(
        \add_260/carry [6]), .S(N140) );
  ADD22 \add_256/U1_1_1  ( .A(i_FIFO[1]), .B(i_FIFO[0]), .CO(
        \add_256/carry [2]), .S(N128) );
  ADD22 \add_256/U1_1_2  ( .A(i_FIFO[2]), .B(\add_256/carry [2]), .CO(
        \add_256/carry [3]), .S(N129) );
  ADD22 \add_256/U1_1_3  ( .A(i_FIFO[3]), .B(\add_256/carry [3]), .CO(
        \add_256/carry [4]), .S(N130) );
  ADD22 \add_256/U1_1_4  ( .A(i_FIFO[4]), .B(\add_256/carry [4]), .CO(
        \add_256/carry [5]), .S(N131) );
  ADD22 \add_256/U1_1_5  ( .A(i_FIFO[5]), .B(\add_256/carry [5]), .CO(
        \add_256/carry [6]), .S(N132) );
  ADD22 \add_255/U1_1_1  ( .A(outWriteCount[1]), .B(outWriteCount[0]), .CO(
        \add_255/carry [2]), .S(N120) );
  ADD22 \add_255/U1_1_2  ( .A(outWriteCount[2]), .B(\add_255/carry [2]), .CO(
        \add_255/carry [3]), .S(N121) );
  ADD22 \add_255/U1_1_3  ( .A(outWriteCount[3]), .B(\add_255/carry [3]), .CO(
        \add_255/carry [4]), .S(N122) );
  ADD22 \add_255/U1_1_4  ( .A(outWriteCount[4]), .B(\add_255/carry [4]), .CO(
        \add_255/carry [5]), .S(N123) );
  ADD22 \add_255/U1_1_5  ( .A(outWriteCount[5]), .B(\add_255/carry [5]), .CO(
        \add_255/carry [6]), .S(N124) );
  ADD22 \add_255/U1_1_6  ( .A(outWriteCount[6]), .B(\add_255/carry [6]), .CO(
        \add_255/carry [7]), .S(N125) );
  ADD32 \r98/U2_1  ( .A(outWriteCount[1]), .B(n549), .CI(\r98/carry [1]), .CO(
        \r98/carry [2]), .S(N144) );
  ADD32 \r98/U2_2  ( .A(outWriteCount[2]), .B(n551), .CI(\r98/carry [2]), .CO(
        \r98/carry [3]), .S(N145) );
  ADD32 \r98/U2_3  ( .A(outWriteCount[3]), .B(n555), .CI(\r98/carry [3]), .CO(
        \r98/carry [4]), .S(N146) );
  ADD32 \r98/U2_4  ( .A(outWriteCount[4]), .B(n554), .CI(\r98/carry [4]), .CO(
        \r98/carry [5]), .S(N147) );
  ADD32 \r98/U2_5  ( .A(outWriteCount[5]), .B(n570), .CI(\r98/carry [5]), .CO(
        \r98/carry [6]), .S(N148) );
  ADD32 \r98/U2_6  ( .A(outWriteCount[6]), .B(n567), .CI(\r98/carry [6]), .CO(
        \r98/carry [7]), .S(N149) );
  DF3 sigEnableCounter_reg ( .D(N198), .C(inClock), .Q(sigEnableCounter), .QN(
        n572) );
  DF3 \currentState_reg[2]  ( .D(N49), .C(inClock), .Q(currentState[2]), .QN(
        n558) );
  DF3 \currentState_reg[0]  ( .D(N47), .C(inClock), .Q(currentState[0]), .QN(
        n548) );
  DF3 \currentState_reg[1]  ( .D(N48), .C(inClock), .Q(currentState[1]), .QN(
        n546) );
  DF3 \currentState_reg[3]  ( .D(N50), .C(inClock), .Q(currentState[3]), .QN(
        n575) );
  DF3 \os1/dff1/s_qout_reg  ( .D(n850), .C(inClock), .Q(\os1/sigQout1 ), .QN(
        n573) );
  DF3 \os2/dff2/s_qout_reg  ( .D(n849), .C(inClock), .Q(\os2/sigQout2 ) );
  DF3 \os2/dff1/s_qout_reg  ( .D(n848), .C(inClock), .Q(\os2/sigQout1 ), .QN(
        n574) );
  DF3 \os1/dff2/s_qout_reg  ( .D(n847), .C(inClock), .Q(\os1/sigQout2 ) );
  DFE1 \FIFO_reg[110][3]  ( .D(n682), .E(N1359), .C(inClock), .Q(
        \FIFO[110][3] ) );
  DFE1 \FIFO_reg[110][2]  ( .D(n682), .E(N1360), .C(inClock), .Q(
        \FIFO[110][2] ) );
  DFE1 \FIFO_reg[110][1]  ( .D(n682), .E(N1361), .C(inClock), .Q(
        \FIFO[110][1] ) );
  DFE1 \FIFO_reg[110][0]  ( .D(n682), .E(N1362), .C(inClock), .Q(
        \FIFO[110][0] ) );
  DFE1 \FIFO_reg[106][3]  ( .D(n684), .E(N1375), .C(inClock), .Q(
        \FIFO[106][3] ) );
  DFE1 \FIFO_reg[106][2]  ( .D(n684), .E(N1376), .C(inClock), .Q(
        \FIFO[106][2] ) );
  DFE1 \FIFO_reg[106][1]  ( .D(n684), .E(N1377), .C(inClock), .Q(
        \FIFO[106][1] ) );
  DFE1 \FIFO_reg[106][0]  ( .D(n684), .E(N1378), .C(inClock), .Q(
        \FIFO[106][0] ) );
  DFE1 \FIFO_reg[102][3]  ( .D(n686), .E(N1391), .C(inClock), .Q(
        \FIFO[102][3] ) );
  DFE1 \FIFO_reg[102][2]  ( .D(n686), .E(N1392), .C(inClock), .Q(
        \FIFO[102][2] ) );
  DFE1 \FIFO_reg[102][1]  ( .D(n686), .E(N1393), .C(inClock), .Q(
        \FIFO[102][1] ) );
  DFE1 \FIFO_reg[102][0]  ( .D(n686), .E(N1394), .C(inClock), .Q(
        \FIFO[102][0] ) );
  DFE1 \FIFO_reg[94][3]  ( .D(n690), .E(N1423), .C(inClock), .Q(\FIFO[94][3] )
         );
  DFE1 \FIFO_reg[94][2]  ( .D(n690), .E(N1424), .C(inClock), .Q(\FIFO[94][2] )
         );
  DFE1 \FIFO_reg[94][1]  ( .D(n690), .E(N1425), .C(inClock), .Q(\FIFO[94][1] )
         );
  DFE1 \FIFO_reg[94][0]  ( .D(n690), .E(N1426), .C(inClock), .Q(\FIFO[94][0] )
         );
  DFE1 \FIFO_reg[90][3]  ( .D(n692), .E(N1439), .C(inClock), .Q(\FIFO[90][3] )
         );
  DFE1 \FIFO_reg[90][2]  ( .D(n692), .E(N1440), .C(inClock), .Q(\FIFO[90][2] )
         );
  DFE1 \FIFO_reg[90][1]  ( .D(n692), .E(N1441), .C(inClock), .Q(\FIFO[90][1] )
         );
  DFE1 \FIFO_reg[90][0]  ( .D(n692), .E(N1442), .C(inClock), .Q(\FIFO[90][0] )
         );
  DFE1 \FIFO_reg[86][3]  ( .D(n694), .E(N1455), .C(inClock), .Q(\FIFO[86][3] )
         );
  DFE1 \FIFO_reg[86][2]  ( .D(n694), .E(N1456), .C(inClock), .Q(\FIFO[86][2] )
         );
  DFE1 \FIFO_reg[86][1]  ( .D(n694), .E(N1457), .C(inClock), .Q(\FIFO[86][1] )
         );
  DFE1 \FIFO_reg[86][0]  ( .D(n694), .E(N1458), .C(inClock), .Q(\FIFO[86][0] )
         );
  DFE1 \FIFO_reg[82][3]  ( .D(n696), .E(N1471), .C(inClock), .Q(\FIFO[82][3] )
         );
  DFE1 \FIFO_reg[82][2]  ( .D(n696), .E(N1472), .C(inClock), .Q(\FIFO[82][2] )
         );
  DFE1 \FIFO_reg[82][1]  ( .D(n696), .E(N1473), .C(inClock), .Q(\FIFO[82][1] )
         );
  DFE1 \FIFO_reg[82][0]  ( .D(n696), .E(N1474), .C(inClock), .Q(\FIFO[82][0] )
         );
  DFE1 \FIFO_reg[78][3]  ( .D(n698), .E(N1487), .C(inClock), .Q(\FIFO[78][3] )
         );
  DFE1 \FIFO_reg[78][2]  ( .D(n698), .E(N1488), .C(inClock), .Q(\FIFO[78][2] )
         );
  DFE1 \FIFO_reg[78][1]  ( .D(n698), .E(N1489), .C(inClock), .Q(\FIFO[78][1] )
         );
  DFE1 \FIFO_reg[78][0]  ( .D(n698), .E(N1490), .C(inClock), .Q(\FIFO[78][0] )
         );
  DFE1 \FIFO_reg[74][3]  ( .D(n700), .E(N1503), .C(inClock), .Q(\FIFO[74][3] )
         );
  DFE1 \FIFO_reg[74][2]  ( .D(n700), .E(N1504), .C(inClock), .Q(\FIFO[74][2] )
         );
  DFE1 \FIFO_reg[74][1]  ( .D(n700), .E(N1505), .C(inClock), .Q(\FIFO[74][1] )
         );
  DFE1 \FIFO_reg[74][0]  ( .D(n700), .E(N1506), .C(inClock), .Q(\FIFO[74][0] )
         );
  DFE1 \FIFO_reg[70][3]  ( .D(n702), .E(N1519), .C(inClock), .Q(\FIFO[70][3] )
         );
  DFE1 \FIFO_reg[70][2]  ( .D(n702), .E(N1520), .C(inClock), .Q(\FIFO[70][2] )
         );
  DFE1 \FIFO_reg[70][1]  ( .D(n702), .E(N1521), .C(inClock), .Q(\FIFO[70][1] )
         );
  DFE1 \FIFO_reg[70][0]  ( .D(n702), .E(N1522), .C(inClock), .Q(\FIFO[70][0] )
         );
  DFE1 \FIFO_reg[62][3]  ( .D(n706), .E(N1551), .C(inClock), .Q(\FIFO[62][3] )
         );
  DFE1 \FIFO_reg[62][2]  ( .D(n706), .E(N1552), .C(inClock), .Q(\FIFO[62][2] )
         );
  DFE1 \FIFO_reg[62][1]  ( .D(n706), .E(N1553), .C(inClock), .Q(\FIFO[62][1] )
         );
  DFE1 \FIFO_reg[62][0]  ( .D(n706), .E(N1554), .C(inClock), .Q(\FIFO[62][0] )
         );
  DFE1 \FIFO_reg[58][3]  ( .D(n708), .E(N1567), .C(inClock), .Q(\FIFO[58][3] )
         );
  DFE1 \FIFO_reg[58][2]  ( .D(n708), .E(N1568), .C(inClock), .Q(\FIFO[58][2] )
         );
  DFE1 \FIFO_reg[58][1]  ( .D(n708), .E(N1569), .C(inClock), .Q(\FIFO[58][1] )
         );
  DFE1 \FIFO_reg[58][0]  ( .D(n708), .E(N1570), .C(inClock), .Q(\FIFO[58][0] )
         );
  DFE1 \FIFO_reg[54][3]  ( .D(n710), .E(N1583), .C(inClock), .Q(\FIFO[54][3] )
         );
  DFE1 \FIFO_reg[54][2]  ( .D(n710), .E(N1584), .C(inClock), .Q(\FIFO[54][2] )
         );
  DFE1 \FIFO_reg[54][1]  ( .D(n710), .E(N1585), .C(inClock), .Q(\FIFO[54][1] )
         );
  DFE1 \FIFO_reg[54][0]  ( .D(n710), .E(N1586), .C(inClock), .Q(\FIFO[54][0] )
         );
  DFE1 \FIFO_reg[50][3]  ( .D(n712), .E(N1599), .C(inClock), .Q(\FIFO[50][3] )
         );
  DFE1 \FIFO_reg[50][2]  ( .D(n712), .E(N1600), .C(inClock), .Q(\FIFO[50][2] )
         );
  DFE1 \FIFO_reg[50][1]  ( .D(n712), .E(N1601), .C(inClock), .Q(\FIFO[50][1] )
         );
  DFE1 \FIFO_reg[50][0]  ( .D(n712), .E(N1602), .C(inClock), .Q(\FIFO[50][0] )
         );
  DFE1 \FIFO_reg[46][3]  ( .D(n714), .E(N1615), .C(inClock), .Q(\FIFO[46][3] )
         );
  DFE1 \FIFO_reg[46][2]  ( .D(n714), .E(N1616), .C(inClock), .Q(\FIFO[46][2] )
         );
  DFE1 \FIFO_reg[46][1]  ( .D(n714), .E(N1617), .C(inClock), .Q(\FIFO[46][1] )
         );
  DFE1 \FIFO_reg[46][0]  ( .D(n714), .E(N1618), .C(inClock), .Q(\FIFO[46][0] )
         );
  DFE1 \FIFO_reg[42][3]  ( .D(n716), .E(N1631), .C(inClock), .Q(\FIFO[42][3] )
         );
  DFE1 \FIFO_reg[42][2]  ( .D(n716), .E(N1632), .C(inClock), .Q(\FIFO[42][2] )
         );
  DFE1 \FIFO_reg[42][1]  ( .D(n716), .E(N1633), .C(inClock), .Q(\FIFO[42][1] )
         );
  DFE1 \FIFO_reg[42][0]  ( .D(n716), .E(N1634), .C(inClock), .Q(\FIFO[42][0] )
         );
  DFE1 \FIFO_reg[38][3]  ( .D(n718), .E(N1647), .C(inClock), .Q(\FIFO[38][3] )
         );
  DFE1 \FIFO_reg[38][2]  ( .D(n718), .E(N1648), .C(inClock), .Q(\FIFO[38][2] )
         );
  DFE1 \FIFO_reg[38][1]  ( .D(n718), .E(N1649), .C(inClock), .Q(\FIFO[38][1] )
         );
  DFE1 \FIFO_reg[38][0]  ( .D(n718), .E(N1650), .C(inClock), .Q(\FIFO[38][0] )
         );
  DFE1 \FIFO_reg[34][3]  ( .D(n720), .E(N1663), .C(inClock), .Q(\FIFO[34][3] )
         );
  DFE1 \FIFO_reg[34][2]  ( .D(n720), .E(N1664), .C(inClock), .Q(\FIFO[34][2] )
         );
  DFE1 \FIFO_reg[34][1]  ( .D(n720), .E(N1665), .C(inClock), .Q(\FIFO[34][1] )
         );
  DFE1 \FIFO_reg[34][0]  ( .D(n720), .E(N1666), .C(inClock), .Q(\FIFO[34][0] )
         );
  DFE1 \FIFO_reg[30][3]  ( .D(n722), .E(N1679), .C(inClock), .Q(\FIFO[30][3] )
         );
  DFE1 \FIFO_reg[30][2]  ( .D(n722), .E(N1680), .C(inClock), .Q(\FIFO[30][2] )
         );
  DFE1 \FIFO_reg[30][1]  ( .D(n722), .E(N1681), .C(inClock), .Q(\FIFO[30][1] )
         );
  DFE1 \FIFO_reg[30][0]  ( .D(n722), .E(N1682), .C(inClock), .Q(\FIFO[30][0] )
         );
  DFE1 \FIFO_reg[26][3]  ( .D(n724), .E(N1695), .C(inClock), .Q(\FIFO[26][3] )
         );
  DFE1 \FIFO_reg[26][2]  ( .D(n724), .E(N1696), .C(inClock), .Q(\FIFO[26][2] )
         );
  DFE1 \FIFO_reg[26][1]  ( .D(n724), .E(N1697), .C(inClock), .Q(\FIFO[26][1] )
         );
  DFE1 \FIFO_reg[26][0]  ( .D(n724), .E(N1698), .C(inClock), .Q(\FIFO[26][0] )
         );
  DFE1 \FIFO_reg[22][3]  ( .D(n726), .E(N1711), .C(inClock), .Q(\FIFO[22][3] )
         );
  DFE1 \FIFO_reg[22][2]  ( .D(n726), .E(N1712), .C(inClock), .Q(\FIFO[22][2] )
         );
  DFE1 \FIFO_reg[22][1]  ( .D(n726), .E(N1713), .C(inClock), .Q(\FIFO[22][1] )
         );
  DFE1 \FIFO_reg[22][0]  ( .D(n726), .E(N1714), .C(inClock), .Q(\FIFO[22][0] )
         );
  DFE1 \FIFO_reg[18][3]  ( .D(n728), .E(N1727), .C(inClock), .Q(\FIFO[18][3] )
         );
  DFE1 \FIFO_reg[18][2]  ( .D(n728), .E(N1728), .C(inClock), .Q(\FIFO[18][2] )
         );
  DFE1 \FIFO_reg[18][1]  ( .D(n728), .E(N1729), .C(inClock), .Q(\FIFO[18][1] )
         );
  DFE1 \FIFO_reg[18][0]  ( .D(n728), .E(N1730), .C(inClock), .Q(\FIFO[18][0] )
         );
  DFE1 \FIFO_reg[14][3]  ( .D(n730), .E(N1743), .C(inClock), .Q(\FIFO[14][3] )
         );
  DFE1 \FIFO_reg[14][2]  ( .D(n730), .E(N1744), .C(inClock), .Q(\FIFO[14][2] )
         );
  DFE1 \FIFO_reg[14][1]  ( .D(n730), .E(N1745), .C(inClock), .Q(\FIFO[14][1] )
         );
  DFE1 \FIFO_reg[14][0]  ( .D(n730), .E(N1746), .C(inClock), .Q(\FIFO[14][0] )
         );
  DFE1 \FIFO_reg[10][3]  ( .D(n732), .E(N1759), .C(inClock), .Q(\FIFO[10][3] )
         );
  DFE1 \FIFO_reg[10][2]  ( .D(n732), .E(N1760), .C(inClock), .Q(\FIFO[10][2] )
         );
  DFE1 \FIFO_reg[10][1]  ( .D(n732), .E(N1761), .C(inClock), .Q(\FIFO[10][1] )
         );
  DFE1 \FIFO_reg[10][0]  ( .D(n732), .E(N1762), .C(inClock), .Q(\FIFO[10][0] )
         );
  DFE1 \FIFO_reg[6][3]  ( .D(n734), .E(N1775), .C(inClock), .Q(\FIFO[6][3] )
         );
  DFE1 \FIFO_reg[6][2]  ( .D(n734), .E(N1776), .C(inClock), .Q(\FIFO[6][2] )
         );
  DFE1 \FIFO_reg[6][1]  ( .D(n734), .E(N1777), .C(inClock), .Q(\FIFO[6][1] )
         );
  DFE1 \FIFO_reg[6][0]  ( .D(n734), .E(N1778), .C(inClock), .Q(\FIFO[6][0] )
         );
  DFE1 \FIFO_reg[2][3]  ( .D(n736), .E(N1791), .C(inClock), .Q(\FIFO[2][3] )
         );
  DFE1 \FIFO_reg[2][2]  ( .D(n736), .E(N1792), .C(inClock), .Q(\FIFO[2][2] )
         );
  DFE1 \FIFO_reg[2][1]  ( .D(n736), .E(N1793), .C(inClock), .Q(\FIFO[2][1] )
         );
  DFE1 \FIFO_reg[2][0]  ( .D(n736), .E(N1794), .C(inClock), .Q(\FIFO[2][0] )
         );
  DFE1 \FIFO_reg[109][3]  ( .D(n683), .E(N1363), .C(inClock), .Q(
        \FIFO[109][3] ) );
  DFE1 \FIFO_reg[109][2]  ( .D(n683), .E(N1364), .C(inClock), .Q(
        \FIFO[109][2] ) );
  DFE1 \FIFO_reg[109][1]  ( .D(n683), .E(N1365), .C(inClock), .Q(
        \FIFO[109][1] ) );
  DFE1 \FIFO_reg[109][0]  ( .D(n683), .E(N1366), .C(inClock), .Q(
        \FIFO[109][0] ) );
  DFE1 \FIFO_reg[108][3]  ( .D(n683), .E(N1367), .C(inClock), .Q(
        \FIFO[108][3] ) );
  DFE1 \FIFO_reg[108][2]  ( .D(n683), .E(N1368), .C(inClock), .Q(
        \FIFO[108][2] ) );
  DFE1 \FIFO_reg[108][1]  ( .D(n683), .E(N1369), .C(inClock), .Q(
        \FIFO[108][1] ) );
  DFE1 \FIFO_reg[108][0]  ( .D(n683), .E(N1370), .C(inClock), .Q(
        \FIFO[108][0] ) );
  DFE1 \FIFO_reg[101][3]  ( .D(n687), .E(N1395), .C(inClock), .Q(
        \FIFO[101][3] ) );
  DFE1 \FIFO_reg[101][2]  ( .D(n687), .E(N1396), .C(inClock), .Q(
        \FIFO[101][2] ) );
  DFE1 \FIFO_reg[101][1]  ( .D(n687), .E(N1397), .C(inClock), .Q(
        \FIFO[101][1] ) );
  DFE1 \FIFO_reg[101][0]  ( .D(n687), .E(N1398), .C(inClock), .Q(
        \FIFO[101][0] ) );
  DFE1 \FIFO_reg[100][3]  ( .D(n687), .E(N1399), .C(inClock), .Q(
        \FIFO[100][3] ) );
  DFE1 \FIFO_reg[100][2]  ( .D(n687), .E(N1400), .C(inClock), .Q(
        \FIFO[100][2] ) );
  DFE1 \FIFO_reg[100][1]  ( .D(n687), .E(N1401), .C(inClock), .Q(
        \FIFO[100][1] ) );
  DFE1 \FIFO_reg[100][0]  ( .D(n687), .E(N1402), .C(inClock), .Q(
        \FIFO[100][0] ) );
  DFE1 \FIFO_reg[95][3]  ( .D(n690), .E(N1419), .C(inClock), .Q(\FIFO[95][3] )
         );
  DFE1 \FIFO_reg[95][2]  ( .D(n690), .E(N1420), .C(inClock), .Q(\FIFO[95][2] )
         );
  DFE1 \FIFO_reg[95][1]  ( .D(n690), .E(N1421), .C(inClock), .Q(\FIFO[95][1] )
         );
  DFE1 \FIFO_reg[95][0]  ( .D(n690), .E(N1422), .C(inClock), .Q(\FIFO[95][0] )
         );
  DFE1 \FIFO_reg[93][3]  ( .D(n691), .E(N1427), .C(inClock), .Q(\FIFO[93][3] )
         );
  DFE1 \FIFO_reg[93][2]  ( .D(n691), .E(N1428), .C(inClock), .Q(\FIFO[93][2] )
         );
  DFE1 \FIFO_reg[93][1]  ( .D(n691), .E(N1429), .C(inClock), .Q(\FIFO[93][1] )
         );
  DFE1 \FIFO_reg[93][0]  ( .D(n691), .E(N1430), .C(inClock), .Q(\FIFO[93][0] )
         );
  DFE1 \FIFO_reg[92][3]  ( .D(n691), .E(N1431), .C(inClock), .Q(\FIFO[92][3] )
         );
  DFE1 \FIFO_reg[92][2]  ( .D(n691), .E(N1432), .C(inClock), .Q(\FIFO[92][2] )
         );
  DFE1 \FIFO_reg[92][1]  ( .D(n691), .E(N1433), .C(inClock), .Q(\FIFO[92][1] )
         );
  DFE1 \FIFO_reg[92][0]  ( .D(n691), .E(N1434), .C(inClock), .Q(\FIFO[92][0] )
         );
  DFE1 \FIFO_reg[89][3]  ( .D(n693), .E(N1443), .C(inClock), .Q(\FIFO[89][3] )
         );
  DFE1 \FIFO_reg[89][2]  ( .D(n693), .E(N1444), .C(inClock), .Q(\FIFO[89][2] )
         );
  DFE1 \FIFO_reg[89][1]  ( .D(n693), .E(N1445), .C(inClock), .Q(\FIFO[89][1] )
         );
  DFE1 \FIFO_reg[89][0]  ( .D(n693), .E(N1446), .C(inClock), .Q(\FIFO[89][0] )
         );
  DFE1 \FIFO_reg[88][3]  ( .D(n693), .E(N1447), .C(inClock), .Q(\FIFO[88][3] )
         );
  DFE1 \FIFO_reg[88][2]  ( .D(n693), .E(N1448), .C(inClock), .Q(\FIFO[88][2] )
         );
  DFE1 \FIFO_reg[88][1]  ( .D(n693), .E(N1449), .C(inClock), .Q(\FIFO[88][1] )
         );
  DFE1 \FIFO_reg[88][0]  ( .D(n693), .E(N1450), .C(inClock), .Q(\FIFO[88][0] )
         );
  DFE1 \FIFO_reg[87][3]  ( .D(n694), .E(N1451), .C(inClock), .Q(\FIFO[87][3] )
         );
  DFE1 \FIFO_reg[87][2]  ( .D(n694), .E(N1452), .C(inClock), .Q(\FIFO[87][2] )
         );
  DFE1 \FIFO_reg[87][1]  ( .D(n694), .E(N1453), .C(inClock), .Q(\FIFO[87][1] )
         );
  DFE1 \FIFO_reg[87][0]  ( .D(n694), .E(N1454), .C(inClock), .Q(\FIFO[87][0] )
         );
  DFE1 \FIFO_reg[85][3]  ( .D(n695), .E(N1459), .C(inClock), .Q(\FIFO[85][3] )
         );
  DFE1 \FIFO_reg[85][2]  ( .D(n695), .E(N1460), .C(inClock), .Q(\FIFO[85][2] )
         );
  DFE1 \FIFO_reg[85][1]  ( .D(n695), .E(N1461), .C(inClock), .Q(\FIFO[85][1] )
         );
  DFE1 \FIFO_reg[85][0]  ( .D(n695), .E(N1462), .C(inClock), .Q(\FIFO[85][0] )
         );
  DFE1 \FIFO_reg[84][3]  ( .D(n695), .E(N1463), .C(inClock), .Q(\FIFO[84][3] )
         );
  DFE1 \FIFO_reg[84][2]  ( .D(n695), .E(N1464), .C(inClock), .Q(\FIFO[84][2] )
         );
  DFE1 \FIFO_reg[84][1]  ( .D(n695), .E(N1465), .C(inClock), .Q(\FIFO[84][1] )
         );
  DFE1 \FIFO_reg[84][0]  ( .D(n695), .E(N1466), .C(inClock), .Q(\FIFO[84][0] )
         );
  DFE1 \FIFO_reg[81][3]  ( .D(n697), .E(N1475), .C(inClock), .Q(\FIFO[81][3] )
         );
  DFE1 \FIFO_reg[81][2]  ( .D(n697), .E(N1476), .C(inClock), .Q(\FIFO[81][2] )
         );
  DFE1 \FIFO_reg[81][1]  ( .D(n697), .E(N1477), .C(inClock), .Q(\FIFO[81][1] )
         );
  DFE1 \FIFO_reg[81][0]  ( .D(n697), .E(N1478), .C(inClock), .Q(\FIFO[81][0] )
         );
  DFE1 \FIFO_reg[80][3]  ( .D(n697), .E(N1479), .C(inClock), .Q(\FIFO[80][3] )
         );
  DFE1 \FIFO_reg[80][2]  ( .D(n697), .E(N1480), .C(inClock), .Q(\FIFO[80][2] )
         );
  DFE1 \FIFO_reg[80][1]  ( .D(n697), .E(N1481), .C(inClock), .Q(\FIFO[80][1] )
         );
  DFE1 \FIFO_reg[80][0]  ( .D(n697), .E(N1482), .C(inClock), .Q(\FIFO[80][0] )
         );
  DFE1 \FIFO_reg[77][3]  ( .D(n699), .E(N1491), .C(inClock), .Q(\FIFO[77][3] )
         );
  DFE1 \FIFO_reg[77][2]  ( .D(n699), .E(N1492), .C(inClock), .Q(\FIFO[77][2] )
         );
  DFE1 \FIFO_reg[77][1]  ( .D(n699), .E(N1493), .C(inClock), .Q(\FIFO[77][1] )
         );
  DFE1 \FIFO_reg[77][0]  ( .D(n699), .E(N1494), .C(inClock), .Q(\FIFO[77][0] )
         );
  DFE1 \FIFO_reg[76][3]  ( .D(n699), .E(N1495), .C(inClock), .Q(\FIFO[76][3] )
         );
  DFE1 \FIFO_reg[76][2]  ( .D(n699), .E(N1496), .C(inClock), .Q(\FIFO[76][2] )
         );
  DFE1 \FIFO_reg[76][1]  ( .D(n699), .E(N1497), .C(inClock), .Q(\FIFO[76][1] )
         );
  DFE1 \FIFO_reg[76][0]  ( .D(n699), .E(N1498), .C(inClock), .Q(\FIFO[76][0] )
         );
  DFE1 \FIFO_reg[69][3]  ( .D(n703), .E(N1523), .C(inClock), .Q(\FIFO[69][3] )
         );
  DFE1 \FIFO_reg[69][2]  ( .D(n703), .E(N1524), .C(inClock), .Q(\FIFO[69][2] )
         );
  DFE1 \FIFO_reg[69][1]  ( .D(n703), .E(N1525), .C(inClock), .Q(\FIFO[69][1] )
         );
  DFE1 \FIFO_reg[69][0]  ( .D(n703), .E(N1526), .C(inClock), .Q(\FIFO[69][0] )
         );
  DFE1 \FIFO_reg[68][3]  ( .D(n703), .E(N1527), .C(inClock), .Q(\FIFO[68][3] )
         );
  DFE1 \FIFO_reg[68][2]  ( .D(n703), .E(N1528), .C(inClock), .Q(\FIFO[68][2] )
         );
  DFE1 \FIFO_reg[68][1]  ( .D(n703), .E(N1529), .C(inClock), .Q(\FIFO[68][1] )
         );
  DFE1 \FIFO_reg[68][0]  ( .D(n703), .E(N1530), .C(inClock), .Q(\FIFO[68][0] )
         );
  DFE1 \FIFO_reg[63][3]  ( .D(n706), .E(N1547), .C(inClock), .Q(\FIFO[63][3] )
         );
  DFE1 \FIFO_reg[63][2]  ( .D(n706), .E(N1548), .C(inClock), .Q(\FIFO[63][2] )
         );
  DFE1 \FIFO_reg[63][1]  ( .D(n706), .E(N1549), .C(inClock), .Q(\FIFO[63][1] )
         );
  DFE1 \FIFO_reg[63][0]  ( .D(n706), .E(N1550), .C(inClock), .Q(\FIFO[63][0] )
         );
  DFE1 \FIFO_reg[61][3]  ( .D(n707), .E(N1555), .C(inClock), .Q(\FIFO[61][3] )
         );
  DFE1 \FIFO_reg[61][2]  ( .D(n707), .E(N1556), .C(inClock), .Q(\FIFO[61][2] )
         );
  DFE1 \FIFO_reg[61][1]  ( .D(n707), .E(N1557), .C(inClock), .Q(\FIFO[61][1] )
         );
  DFE1 \FIFO_reg[61][0]  ( .D(n707), .E(N1558), .C(inClock), .Q(\FIFO[61][0] )
         );
  DFE1 \FIFO_reg[60][3]  ( .D(n707), .E(N1559), .C(inClock), .Q(\FIFO[60][3] )
         );
  DFE1 \FIFO_reg[60][2]  ( .D(n707), .E(N1560), .C(inClock), .Q(\FIFO[60][2] )
         );
  DFE1 \FIFO_reg[60][1]  ( .D(n707), .E(N1561), .C(inClock), .Q(\FIFO[60][1] )
         );
  DFE1 \FIFO_reg[60][0]  ( .D(n707), .E(N1562), .C(inClock), .Q(\FIFO[60][0] )
         );
  DFE1 \FIFO_reg[57][3]  ( .D(n709), .E(N1571), .C(inClock), .Q(\FIFO[57][3] )
         );
  DFE1 \FIFO_reg[57][2]  ( .D(n709), .E(N1572), .C(inClock), .Q(\FIFO[57][2] )
         );
  DFE1 \FIFO_reg[57][1]  ( .D(n709), .E(N1573), .C(inClock), .Q(\FIFO[57][1] )
         );
  DFE1 \FIFO_reg[57][0]  ( .D(n709), .E(N1574), .C(inClock), .Q(\FIFO[57][0] )
         );
  DFE1 \FIFO_reg[56][3]  ( .D(n709), .E(N1575), .C(inClock), .Q(\FIFO[56][3] )
         );
  DFE1 \FIFO_reg[56][2]  ( .D(n709), .E(N1576), .C(inClock), .Q(\FIFO[56][2] )
         );
  DFE1 \FIFO_reg[56][1]  ( .D(n709), .E(N1577), .C(inClock), .Q(\FIFO[56][1] )
         );
  DFE1 \FIFO_reg[56][0]  ( .D(n709), .E(N1578), .C(inClock), .Q(\FIFO[56][0] )
         );
  DFE1 \FIFO_reg[55][3]  ( .D(n710), .E(N1579), .C(inClock), .Q(\FIFO[55][3] )
         );
  DFE1 \FIFO_reg[55][2]  ( .D(n710), .E(N1580), .C(inClock), .Q(\FIFO[55][2] )
         );
  DFE1 \FIFO_reg[55][1]  ( .D(n710), .E(N1581), .C(inClock), .Q(\FIFO[55][1] )
         );
  DFE1 \FIFO_reg[55][0]  ( .D(n710), .E(N1582), .C(inClock), .Q(\FIFO[55][0] )
         );
  DFE1 \FIFO_reg[53][3]  ( .D(n711), .E(N1587), .C(inClock), .Q(\FIFO[53][3] )
         );
  DFE1 \FIFO_reg[53][2]  ( .D(n711), .E(N1588), .C(inClock), .Q(\FIFO[53][2] )
         );
  DFE1 \FIFO_reg[53][1]  ( .D(n711), .E(N1589), .C(inClock), .Q(\FIFO[53][1] )
         );
  DFE1 \FIFO_reg[53][0]  ( .D(n711), .E(N1590), .C(inClock), .Q(\FIFO[53][0] )
         );
  DFE1 \FIFO_reg[52][3]  ( .D(n711), .E(N1591), .C(inClock), .Q(\FIFO[52][3] )
         );
  DFE1 \FIFO_reg[52][2]  ( .D(n711), .E(N1592), .C(inClock), .Q(\FIFO[52][2] )
         );
  DFE1 \FIFO_reg[52][1]  ( .D(n711), .E(N1593), .C(inClock), .Q(\FIFO[52][1] )
         );
  DFE1 \FIFO_reg[52][0]  ( .D(n711), .E(N1594), .C(inClock), .Q(\FIFO[52][0] )
         );
  DFE1 \FIFO_reg[49][3]  ( .D(n713), .E(N1603), .C(inClock), .Q(\FIFO[49][3] )
         );
  DFE1 \FIFO_reg[49][2]  ( .D(n713), .E(N1604), .C(inClock), .Q(\FIFO[49][2] )
         );
  DFE1 \FIFO_reg[49][1]  ( .D(n713), .E(N1605), .C(inClock), .Q(\FIFO[49][1] )
         );
  DFE1 \FIFO_reg[49][0]  ( .D(n713), .E(N1606), .C(inClock), .Q(\FIFO[49][0] )
         );
  DFE1 \FIFO_reg[48][3]  ( .D(n713), .E(N1607), .C(inClock), .Q(\FIFO[48][3] )
         );
  DFE1 \FIFO_reg[48][2]  ( .D(n713), .E(N1608), .C(inClock), .Q(\FIFO[48][2] )
         );
  DFE1 \FIFO_reg[48][1]  ( .D(n713), .E(N1609), .C(inClock), .Q(\FIFO[48][1] )
         );
  DFE1 \FIFO_reg[48][0]  ( .D(n713), .E(N1610), .C(inClock), .Q(\FIFO[48][0] )
         );
  DFE1 \FIFO_reg[47][3]  ( .D(n714), .E(N1611), .C(inClock), .Q(\FIFO[47][3] )
         );
  DFE1 \FIFO_reg[47][2]  ( .D(n714), .E(N1612), .C(inClock), .Q(\FIFO[47][2] )
         );
  DFE1 \FIFO_reg[47][1]  ( .D(n714), .E(N1613), .C(inClock), .Q(\FIFO[47][1] )
         );
  DFE1 \FIFO_reg[47][0]  ( .D(n714), .E(N1614), .C(inClock), .Q(\FIFO[47][0] )
         );
  DFE1 \FIFO_reg[45][3]  ( .D(n715), .E(N1619), .C(inClock), .Q(\FIFO[45][3] )
         );
  DFE1 \FIFO_reg[45][2]  ( .D(n715), .E(N1620), .C(inClock), .Q(\FIFO[45][2] )
         );
  DFE1 \FIFO_reg[45][1]  ( .D(n715), .E(N1621), .C(inClock), .Q(\FIFO[45][1] )
         );
  DFE1 \FIFO_reg[45][0]  ( .D(n715), .E(N1622), .C(inClock), .Q(\FIFO[45][0] )
         );
  DFE1 \FIFO_reg[44][3]  ( .D(n715), .E(N1623), .C(inClock), .Q(\FIFO[44][3] )
         );
  DFE1 \FIFO_reg[44][2]  ( .D(n715), .E(N1624), .C(inClock), .Q(\FIFO[44][2] )
         );
  DFE1 \FIFO_reg[44][1]  ( .D(n715), .E(N1625), .C(inClock), .Q(\FIFO[44][1] )
         );
  DFE1 \FIFO_reg[44][0]  ( .D(n715), .E(N1626), .C(inClock), .Q(\FIFO[44][0] )
         );
  DFE1 \FIFO_reg[43][3]  ( .D(n716), .E(N1627), .C(inClock), .Q(\FIFO[43][3] )
         );
  DFE1 \FIFO_reg[43][2]  ( .D(n716), .E(N1628), .C(inClock), .Q(\FIFO[43][2] )
         );
  DFE1 \FIFO_reg[43][1]  ( .D(n716), .E(N1629), .C(inClock), .Q(\FIFO[43][1] )
         );
  DFE1 \FIFO_reg[43][0]  ( .D(n716), .E(N1630), .C(inClock), .Q(\FIFO[43][0] )
         );
  DFE1 \FIFO_reg[41][3]  ( .D(n717), .E(N1635), .C(inClock), .Q(\FIFO[41][3] )
         );
  DFE1 \FIFO_reg[41][2]  ( .D(n717), .E(N1636), .C(inClock), .Q(\FIFO[41][2] )
         );
  DFE1 \FIFO_reg[41][1]  ( .D(n717), .E(N1637), .C(inClock), .Q(\FIFO[41][1] )
         );
  DFE1 \FIFO_reg[41][0]  ( .D(n717), .E(N1638), .C(inClock), .Q(\FIFO[41][0] )
         );
  DFE1 \FIFO_reg[40][3]  ( .D(n717), .E(N1639), .C(inClock), .Q(\FIFO[40][3] )
         );
  DFE1 \FIFO_reg[40][2]  ( .D(n717), .E(N1640), .C(inClock), .Q(\FIFO[40][2] )
         );
  DFE1 \FIFO_reg[40][1]  ( .D(n717), .E(N1641), .C(inClock), .Q(\FIFO[40][1] )
         );
  DFE1 \FIFO_reg[40][0]  ( .D(n717), .E(N1642), .C(inClock), .Q(\FIFO[40][0] )
         );
  DFE1 \FIFO_reg[39][3]  ( .D(n718), .E(N1643), .C(inClock), .Q(\FIFO[39][3] )
         );
  DFE1 \FIFO_reg[39][2]  ( .D(n718), .E(N1644), .C(inClock), .Q(\FIFO[39][2] )
         );
  DFE1 \FIFO_reg[39][1]  ( .D(n718), .E(N1645), .C(inClock), .Q(\FIFO[39][1] )
         );
  DFE1 \FIFO_reg[39][0]  ( .D(n718), .E(N1646), .C(inClock), .Q(\FIFO[39][0] )
         );
  DFE1 \FIFO_reg[37][3]  ( .D(n719), .E(N1651), .C(inClock), .Q(\FIFO[37][3] )
         );
  DFE1 \FIFO_reg[37][2]  ( .D(n719), .E(N1652), .C(inClock), .Q(\FIFO[37][2] )
         );
  DFE1 \FIFO_reg[37][1]  ( .D(n719), .E(N1653), .C(inClock), .Q(\FIFO[37][1] )
         );
  DFE1 \FIFO_reg[37][0]  ( .D(n719), .E(N1654), .C(inClock), .Q(\FIFO[37][0] )
         );
  DFE1 \FIFO_reg[36][3]  ( .D(n719), .E(N1655), .C(inClock), .Q(\FIFO[36][3] )
         );
  DFE1 \FIFO_reg[36][2]  ( .D(n719), .E(N1656), .C(inClock), .Q(\FIFO[36][2] )
         );
  DFE1 \FIFO_reg[36][1]  ( .D(n719), .E(N1657), .C(inClock), .Q(\FIFO[36][1] )
         );
  DFE1 \FIFO_reg[36][0]  ( .D(n719), .E(N1658), .C(inClock), .Q(\FIFO[36][0] )
         );
  DFE1 \FIFO_reg[35][3]  ( .D(n720), .E(N1659), .C(inClock), .Q(\FIFO[35][3] )
         );
  DFE1 \FIFO_reg[35][2]  ( .D(n720), .E(N1660), .C(inClock), .Q(\FIFO[35][2] )
         );
  DFE1 \FIFO_reg[35][1]  ( .D(n720), .E(N1661), .C(inClock), .Q(\FIFO[35][1] )
         );
  DFE1 \FIFO_reg[35][0]  ( .D(n720), .E(N1662), .C(inClock), .Q(\FIFO[35][0] )
         );
  DFE1 \FIFO_reg[33][3]  ( .D(n721), .E(N1667), .C(inClock), .Q(\FIFO[33][3] )
         );
  DFE1 \FIFO_reg[33][2]  ( .D(n721), .E(N1668), .C(inClock), .Q(\FIFO[33][2] )
         );
  DFE1 \FIFO_reg[33][1]  ( .D(n721), .E(N1669), .C(inClock), .Q(\FIFO[33][1] )
         );
  DFE1 \FIFO_reg[33][0]  ( .D(n721), .E(N1670), .C(inClock), .Q(\FIFO[33][0] )
         );
  DFE1 \FIFO_reg[32][3]  ( .D(n721), .E(N1671), .C(inClock), .Q(\FIFO[32][3] )
         );
  DFE1 \FIFO_reg[32][2]  ( .D(n721), .E(N1672), .C(inClock), .Q(\FIFO[32][2] )
         );
  DFE1 \FIFO_reg[32][1]  ( .D(n721), .E(N1673), .C(inClock), .Q(\FIFO[32][1] )
         );
  DFE1 \FIFO_reg[32][0]  ( .D(n721), .E(N1674), .C(inClock), .Q(\FIFO[32][0] )
         );
  DFE1 \FIFO_reg[31][3]  ( .D(n722), .E(N1675), .C(inClock), .Q(\FIFO[31][3] )
         );
  DFE1 \FIFO_reg[31][2]  ( .D(n722), .E(N1676), .C(inClock), .Q(\FIFO[31][2] )
         );
  DFE1 \FIFO_reg[31][1]  ( .D(n722), .E(N1677), .C(inClock), .Q(\FIFO[31][1] )
         );
  DFE1 \FIFO_reg[31][0]  ( .D(n722), .E(N1678), .C(inClock), .Q(\FIFO[31][0] )
         );
  DFE1 \FIFO_reg[29][3]  ( .D(n723), .E(N1683), .C(inClock), .Q(\FIFO[29][3] )
         );
  DFE1 \FIFO_reg[29][2]  ( .D(n723), .E(N1684), .C(inClock), .Q(\FIFO[29][2] )
         );
  DFE1 \FIFO_reg[29][1]  ( .D(n723), .E(N1685), .C(inClock), .Q(\FIFO[29][1] )
         );
  DFE1 \FIFO_reg[29][0]  ( .D(n723), .E(N1686), .C(inClock), .Q(\FIFO[29][0] )
         );
  DFE1 \FIFO_reg[28][3]  ( .D(n723), .E(N1687), .C(inClock), .Q(\FIFO[28][3] )
         );
  DFE1 \FIFO_reg[28][2]  ( .D(n723), .E(N1688), .C(inClock), .Q(\FIFO[28][2] )
         );
  DFE1 \FIFO_reg[28][1]  ( .D(n723), .E(N1689), .C(inClock), .Q(\FIFO[28][1] )
         );
  DFE1 \FIFO_reg[28][0]  ( .D(n723), .E(N1690), .C(inClock), .Q(\FIFO[28][0] )
         );
  DFE1 \FIFO_reg[27][3]  ( .D(n724), .E(N1691), .C(inClock), .Q(\FIFO[27][3] )
         );
  DFE1 \FIFO_reg[27][2]  ( .D(n724), .E(N1692), .C(inClock), .Q(\FIFO[27][2] )
         );
  DFE1 \FIFO_reg[27][1]  ( .D(n724), .E(N1693), .C(inClock), .Q(\FIFO[27][1] )
         );
  DFE1 \FIFO_reg[27][0]  ( .D(n724), .E(N1694), .C(inClock), .Q(\FIFO[27][0] )
         );
  DFE1 \FIFO_reg[25][3]  ( .D(n725), .E(N1699), .C(inClock), .Q(\FIFO[25][3] )
         );
  DFE1 \FIFO_reg[25][2]  ( .D(n725), .E(N1700), .C(inClock), .Q(\FIFO[25][2] )
         );
  DFE1 \FIFO_reg[25][1]  ( .D(n725), .E(N1701), .C(inClock), .Q(\FIFO[25][1] )
         );
  DFE1 \FIFO_reg[25][0]  ( .D(n725), .E(N1702), .C(inClock), .Q(\FIFO[25][0] )
         );
  DFE1 \FIFO_reg[24][3]  ( .D(n725), .E(N1703), .C(inClock), .Q(\FIFO[24][3] )
         );
  DFE1 \FIFO_reg[24][2]  ( .D(n725), .E(N1704), .C(inClock), .Q(\FIFO[24][2] )
         );
  DFE1 \FIFO_reg[24][1]  ( .D(n725), .E(N1705), .C(inClock), .Q(\FIFO[24][1] )
         );
  DFE1 \FIFO_reg[24][0]  ( .D(n725), .E(N1706), .C(inClock), .Q(\FIFO[24][0] )
         );
  DFE1 \FIFO_reg[23][3]  ( .D(n726), .E(N1707), .C(inClock), .Q(\FIFO[23][3] )
         );
  DFE1 \FIFO_reg[23][2]  ( .D(n726), .E(N1708), .C(inClock), .Q(\FIFO[23][2] )
         );
  DFE1 \FIFO_reg[23][1]  ( .D(n726), .E(N1709), .C(inClock), .Q(\FIFO[23][1] )
         );
  DFE1 \FIFO_reg[23][0]  ( .D(n726), .E(N1710), .C(inClock), .Q(\FIFO[23][0] )
         );
  DFE1 \FIFO_reg[21][3]  ( .D(n727), .E(N1715), .C(inClock), .Q(\FIFO[21][3] )
         );
  DFE1 \FIFO_reg[21][2]  ( .D(n727), .E(N1716), .C(inClock), .Q(\FIFO[21][2] )
         );
  DFE1 \FIFO_reg[21][1]  ( .D(n727), .E(N1717), .C(inClock), .Q(\FIFO[21][1] )
         );
  DFE1 \FIFO_reg[21][0]  ( .D(n727), .E(N1718), .C(inClock), .Q(\FIFO[21][0] )
         );
  DFE1 \FIFO_reg[20][3]  ( .D(n727), .E(N1719), .C(inClock), .Q(\FIFO[20][3] )
         );
  DFE1 \FIFO_reg[20][2]  ( .D(n727), .E(N1720), .C(inClock), .Q(\FIFO[20][2] )
         );
  DFE1 \FIFO_reg[20][1]  ( .D(n727), .E(N1721), .C(inClock), .Q(\FIFO[20][1] )
         );
  DFE1 \FIFO_reg[20][0]  ( .D(n727), .E(N1722), .C(inClock), .Q(\FIFO[20][0] )
         );
  DFE1 \FIFO_reg[19][3]  ( .D(n728), .E(N1723), .C(inClock), .Q(\FIFO[19][3] )
         );
  DFE1 \FIFO_reg[19][2]  ( .D(n728), .E(N1724), .C(inClock), .Q(\FIFO[19][2] )
         );
  DFE1 \FIFO_reg[19][1]  ( .D(n728), .E(N1725), .C(inClock), .Q(\FIFO[19][1] )
         );
  DFE1 \FIFO_reg[19][0]  ( .D(n728), .E(N1726), .C(inClock), .Q(\FIFO[19][0] )
         );
  DFE1 \FIFO_reg[17][3]  ( .D(n729), .E(N1731), .C(inClock), .Q(\FIFO[17][3] )
         );
  DFE1 \FIFO_reg[17][2]  ( .D(n729), .E(N1732), .C(inClock), .Q(\FIFO[17][2] )
         );
  DFE1 \FIFO_reg[17][1]  ( .D(n729), .E(N1733), .C(inClock), .Q(\FIFO[17][1] )
         );
  DFE1 \FIFO_reg[17][0]  ( .D(n729), .E(N1734), .C(inClock), .Q(\FIFO[17][0] )
         );
  DFE1 \FIFO_reg[16][3]  ( .D(n729), .E(N1735), .C(inClock), .Q(\FIFO[16][3] )
         );
  DFE1 \FIFO_reg[16][2]  ( .D(n729), .E(N1736), .C(inClock), .Q(\FIFO[16][2] )
         );
  DFE1 \FIFO_reg[16][1]  ( .D(n729), .E(N1737), .C(inClock), .Q(\FIFO[16][1] )
         );
  DFE1 \FIFO_reg[16][0]  ( .D(n729), .E(N1738), .C(inClock), .Q(\FIFO[16][0] )
         );
  DFE1 \FIFO_reg[15][3]  ( .D(n730), .E(N1739), .C(inClock), .Q(\FIFO[15][3] )
         );
  DFE1 \FIFO_reg[15][2]  ( .D(n730), .E(N1740), .C(inClock), .Q(\FIFO[15][2] )
         );
  DFE1 \FIFO_reg[15][1]  ( .D(n730), .E(N1741), .C(inClock), .Q(\FIFO[15][1] )
         );
  DFE1 \FIFO_reg[15][0]  ( .D(n730), .E(N1742), .C(inClock), .Q(\FIFO[15][0] )
         );
  DFE1 \FIFO_reg[13][3]  ( .D(n731), .E(N1747), .C(inClock), .Q(\FIFO[13][3] )
         );
  DFE1 \FIFO_reg[13][2]  ( .D(n731), .E(N1748), .C(inClock), .Q(\FIFO[13][2] )
         );
  DFE1 \FIFO_reg[13][1]  ( .D(n731), .E(N1749), .C(inClock), .Q(\FIFO[13][1] )
         );
  DFE1 \FIFO_reg[13][0]  ( .D(n731), .E(N1750), .C(inClock), .Q(\FIFO[13][0] )
         );
  DFE1 \FIFO_reg[12][3]  ( .D(n731), .E(N1751), .C(inClock), .Q(\FIFO[12][3] )
         );
  DFE1 \FIFO_reg[12][2]  ( .D(n731), .E(N1752), .C(inClock), .Q(\FIFO[12][2] )
         );
  DFE1 \FIFO_reg[12][1]  ( .D(n731), .E(N1753), .C(inClock), .Q(\FIFO[12][1] )
         );
  DFE1 \FIFO_reg[12][0]  ( .D(n731), .E(N1754), .C(inClock), .Q(\FIFO[12][0] )
         );
  DFE1 \FIFO_reg[11][3]  ( .D(n732), .E(N1755), .C(inClock), .Q(\FIFO[11][3] )
         );
  DFE1 \FIFO_reg[11][2]  ( .D(n732), .E(N1756), .C(inClock), .Q(\FIFO[11][2] )
         );
  DFE1 \FIFO_reg[11][1]  ( .D(n732), .E(N1757), .C(inClock), .Q(\FIFO[11][1] )
         );
  DFE1 \FIFO_reg[11][0]  ( .D(n732), .E(N1758), .C(inClock), .Q(\FIFO[11][0] )
         );
  DFE1 \FIFO_reg[9][3]  ( .D(n733), .E(N1763), .C(inClock), .Q(\FIFO[9][3] )
         );
  DFE1 \FIFO_reg[9][2]  ( .D(n733), .E(N1764), .C(inClock), .Q(\FIFO[9][2] )
         );
  DFE1 \FIFO_reg[9][1]  ( .D(n733), .E(N1765), .C(inClock), .Q(\FIFO[9][1] )
         );
  DFE1 \FIFO_reg[9][0]  ( .D(n733), .E(N1766), .C(inClock), .Q(\FIFO[9][0] )
         );
  DFE1 \FIFO_reg[8][3]  ( .D(n733), .E(N1767), .C(inClock), .Q(\FIFO[8][3] )
         );
  DFE1 \FIFO_reg[8][2]  ( .D(n733), .E(N1768), .C(inClock), .Q(\FIFO[8][2] )
         );
  DFE1 \FIFO_reg[8][1]  ( .D(n733), .E(N1769), .C(inClock), .Q(\FIFO[8][1] )
         );
  DFE1 \FIFO_reg[8][0]  ( .D(n733), .E(N1770), .C(inClock), .Q(\FIFO[8][0] )
         );
  DFE1 \FIFO_reg[7][3]  ( .D(n734), .E(N1771), .C(inClock), .Q(\FIFO[7][3] )
         );
  DFE1 \FIFO_reg[7][2]  ( .D(n734), .E(N1772), .C(inClock), .Q(\FIFO[7][2] )
         );
  DFE1 \FIFO_reg[7][1]  ( .D(n734), .E(N1773), .C(inClock), .Q(\FIFO[7][1] )
         );
  DFE1 \FIFO_reg[7][0]  ( .D(n734), .E(N1774), .C(inClock), .Q(\FIFO[7][0] )
         );
  DFE1 \FIFO_reg[5][3]  ( .D(n735), .E(N1779), .C(inClock), .Q(\FIFO[5][3] )
         );
  DFE1 \FIFO_reg[5][2]  ( .D(n735), .E(N1780), .C(inClock), .Q(\FIFO[5][2] )
         );
  DFE1 \FIFO_reg[5][1]  ( .D(n735), .E(N1781), .C(inClock), .Q(\FIFO[5][1] )
         );
  DFE1 \FIFO_reg[5][0]  ( .D(n735), .E(N1782), .C(inClock), .Q(\FIFO[5][0] )
         );
  DFE1 \FIFO_reg[4][3]  ( .D(n735), .E(N1783), .C(inClock), .Q(\FIFO[4][3] )
         );
  DFE1 \FIFO_reg[4][2]  ( .D(n735), .E(N1784), .C(inClock), .Q(\FIFO[4][2] )
         );
  DFE1 \FIFO_reg[4][1]  ( .D(n735), .E(N1785), .C(inClock), .Q(\FIFO[4][1] )
         );
  DFE1 \FIFO_reg[4][0]  ( .D(n735), .E(N1786), .C(inClock), .Q(\FIFO[4][0] )
         );
  DFE1 \FIFO_reg[3][3]  ( .D(n736), .E(N1787), .C(inClock), .Q(\FIFO[3][3] )
         );
  DFE1 \FIFO_reg[3][2]  ( .D(n736), .E(N1788), .C(inClock), .Q(\FIFO[3][2] )
         );
  DFE1 \FIFO_reg[3][1]  ( .D(n736), .E(N1789), .C(inClock), .Q(\FIFO[3][1] )
         );
  DFE1 \FIFO_reg[3][0]  ( .D(n736), .E(N1790), .C(inClock), .Q(\FIFO[3][0] )
         );
  DFE1 \FIFO_reg[1][3]  ( .D(n737), .E(N1795), .C(inClock), .Q(\FIFO[1][3] )
         );
  DFE1 \FIFO_reg[1][2]  ( .D(n737), .E(N1796), .C(inClock), .Q(\FIFO[1][2] )
         );
  DFE1 \FIFO_reg[1][1]  ( .D(n737), .E(N1797), .C(inClock), .Q(\FIFO[1][1] )
         );
  DFE1 \FIFO_reg[1][0]  ( .D(n737), .E(N1798), .C(inClock), .Q(\FIFO[1][0] )
         );
  DFE1 \FIFO_reg[0][3]  ( .D(n737), .E(N1799), .C(inClock), .Q(\FIFO[0][3] )
         );
  DFE1 \FIFO_reg[0][2]  ( .D(n737), .E(N1800), .C(inClock), .Q(\FIFO[0][2] )
         );
  DFE1 \FIFO_reg[0][1]  ( .D(n737), .E(N1801), .C(inClock), .Q(\FIFO[0][1] )
         );
  DFE1 \FIFO_reg[0][0]  ( .D(n737), .E(N1802), .C(inClock), .Q(\FIFO[0][0] )
         );
  DFE1 \j_FIFO_reg[5]  ( .D(N227), .E(N213), .C(inClock), .Q(N44) );
  DFE1 \j_FIFO_reg[6]  ( .D(N228), .E(N213), .C(inClock), .Q(N45) );
  DFE1 \FIFO_reg[126][3]  ( .D(n674), .E(N1295), .C(inClock), .Q(
        \FIFO[126][3] ) );
  DFE1 \FIFO_reg[126][2]  ( .D(n674), .E(N1296), .C(inClock), .Q(
        \FIFO[126][2] ) );
  DFE1 \FIFO_reg[126][1]  ( .D(n674), .E(N1297), .C(inClock), .Q(
        \FIFO[126][1] ) );
  DFE1 \FIFO_reg[126][0]  ( .D(n674), .E(N1298), .C(inClock), .Q(
        \FIFO[126][0] ) );
  DFE1 \FIFO_reg[122][3]  ( .D(n676), .E(N1311), .C(inClock), .Q(
        \FIFO[122][3] ) );
  DFE1 \FIFO_reg[122][2]  ( .D(n676), .E(N1312), .C(inClock), .Q(
        \FIFO[122][2] ) );
  DFE1 \FIFO_reg[122][1]  ( .D(n676), .E(N1313), .C(inClock), .Q(
        \FIFO[122][1] ) );
  DFE1 \FIFO_reg[122][0]  ( .D(n676), .E(N1314), .C(inClock), .Q(
        \FIFO[122][0] ) );
  DFE1 \FIFO_reg[118][3]  ( .D(n678), .E(N1327), .C(inClock), .Q(
        \FIFO[118][3] ) );
  DFE1 \FIFO_reg[118][2]  ( .D(n678), .E(N1328), .C(inClock), .Q(
        \FIFO[118][2] ) );
  DFE1 \FIFO_reg[118][1]  ( .D(n678), .E(N1329), .C(inClock), .Q(
        \FIFO[118][1] ) );
  DFE1 \FIFO_reg[118][0]  ( .D(n678), .E(N1330), .C(inClock), .Q(
        \FIFO[118][0] ) );
  DFE1 \FIFO_reg[114][3]  ( .D(n680), .E(N1343), .C(inClock), .Q(
        \FIFO[114][3] ) );
  DFE1 \FIFO_reg[114][2]  ( .D(n680), .E(N1344), .C(inClock), .Q(
        \FIFO[114][2] ) );
  DFE1 \FIFO_reg[114][1]  ( .D(n680), .E(N1345), .C(inClock), .Q(
        \FIFO[114][1] ) );
  DFE1 \FIFO_reg[114][0]  ( .D(n680), .E(N1346), .C(inClock), .Q(
        \FIFO[114][0] ) );
  DFE1 \FIFO_reg[98][3]  ( .D(n688), .E(N1407), .C(inClock), .Q(\FIFO[98][3] )
         );
  DFE1 \FIFO_reg[98][2]  ( .D(n688), .E(N1408), .C(inClock), .Q(\FIFO[98][2] )
         );
  DFE1 \FIFO_reg[98][1]  ( .D(n688), .E(N1409), .C(inClock), .Q(\FIFO[98][1] )
         );
  DFE1 \FIFO_reg[98][0]  ( .D(n688), .E(N1410), .C(inClock), .Q(\FIFO[98][0] )
         );
  DFE1 \FIFO_reg[66][3]  ( .D(n704), .E(N1535), .C(inClock), .Q(\FIFO[66][3] )
         );
  DFE1 \FIFO_reg[66][2]  ( .D(n704), .E(N1536), .C(inClock), .Q(\FIFO[66][2] )
         );
  DFE1 \FIFO_reg[66][1]  ( .D(n704), .E(N1537), .C(inClock), .Q(\FIFO[66][1] )
         );
  DFE1 \FIFO_reg[66][0]  ( .D(n704), .E(N1538), .C(inClock), .Q(\FIFO[66][0] )
         );
  DFE1 \FIFO_reg[127][3]  ( .D(n674), .E(N1291), .C(inClock), .Q(
        \FIFO[127][3] ) );
  DFE1 \FIFO_reg[127][2]  ( .D(n674), .E(N1292), .C(inClock), .Q(
        \FIFO[127][2] ) );
  DFE1 \FIFO_reg[127][1]  ( .D(n674), .E(N1293), .C(inClock), .Q(
        \FIFO[127][1] ) );
  DFE1 \FIFO_reg[127][0]  ( .D(n674), .E(N1294), .C(inClock), .Q(
        \FIFO[127][0] ) );
  DFE1 \FIFO_reg[125][3]  ( .D(n675), .E(N1299), .C(inClock), .Q(
        \FIFO[125][3] ) );
  DFE1 \FIFO_reg[125][2]  ( .D(n675), .E(N1300), .C(inClock), .Q(
        \FIFO[125][2] ) );
  DFE1 \FIFO_reg[125][1]  ( .D(n675), .E(N1301), .C(inClock), .Q(
        \FIFO[125][1] ) );
  DFE1 \FIFO_reg[125][0]  ( .D(n675), .E(N1302), .C(inClock), .Q(
        \FIFO[125][0] ) );
  DFE1 \FIFO_reg[124][3]  ( .D(n675), .E(N1303), .C(inClock), .Q(
        \FIFO[124][3] ) );
  DFE1 \FIFO_reg[124][2]  ( .D(n675), .E(N1304), .C(inClock), .Q(
        \FIFO[124][2] ) );
  DFE1 \FIFO_reg[124][1]  ( .D(n675), .E(N1305), .C(inClock), .Q(
        \FIFO[124][1] ) );
  DFE1 \FIFO_reg[124][0]  ( .D(n675), .E(N1306), .C(inClock), .Q(
        \FIFO[124][0] ) );
  DFE1 \FIFO_reg[123][3]  ( .D(n676), .E(N1307), .C(inClock), .Q(
        \FIFO[123][3] ) );
  DFE1 \FIFO_reg[123][2]  ( .D(n676), .E(N1308), .C(inClock), .Q(
        \FIFO[123][2] ) );
  DFE1 \FIFO_reg[123][1]  ( .D(n676), .E(N1309), .C(inClock), .Q(
        \FIFO[123][1] ) );
  DFE1 \FIFO_reg[123][0]  ( .D(n676), .E(N1310), .C(inClock), .Q(
        \FIFO[123][0] ) );
  DFE1 \FIFO_reg[121][3]  ( .D(n677), .E(N1315), .C(inClock), .Q(
        \FIFO[121][3] ) );
  DFE1 \FIFO_reg[121][2]  ( .D(n677), .E(N1316), .C(inClock), .Q(
        \FIFO[121][2] ) );
  DFE1 \FIFO_reg[121][1]  ( .D(n677), .E(N1317), .C(inClock), .Q(
        \FIFO[121][1] ) );
  DFE1 \FIFO_reg[121][0]  ( .D(n677), .E(N1318), .C(inClock), .Q(
        \FIFO[121][0] ) );
  DFE1 \FIFO_reg[120][3]  ( .D(n677), .E(N1319), .C(inClock), .Q(
        \FIFO[120][3] ) );
  DFE1 \FIFO_reg[120][2]  ( .D(n677), .E(N1320), .C(inClock), .Q(
        \FIFO[120][2] ) );
  DFE1 \FIFO_reg[120][1]  ( .D(n677), .E(N1321), .C(inClock), .Q(
        \FIFO[120][1] ) );
  DFE1 \FIFO_reg[120][0]  ( .D(n677), .E(N1322), .C(inClock), .Q(
        \FIFO[120][0] ) );
  DFE1 \FIFO_reg[119][3]  ( .D(n678), .E(N1323), .C(inClock), .Q(
        \FIFO[119][3] ) );
  DFE1 \FIFO_reg[119][2]  ( .D(n678), .E(N1324), .C(inClock), .Q(
        \FIFO[119][2] ) );
  DFE1 \FIFO_reg[119][1]  ( .D(n678), .E(N1325), .C(inClock), .Q(
        \FIFO[119][1] ) );
  DFE1 \FIFO_reg[119][0]  ( .D(n678), .E(N1326), .C(inClock), .Q(
        \FIFO[119][0] ) );
  DFE1 \FIFO_reg[117][3]  ( .D(n679), .E(N1331), .C(inClock), .Q(
        \FIFO[117][3] ) );
  DFE1 \FIFO_reg[117][2]  ( .D(n679), .E(N1332), .C(inClock), .Q(
        \FIFO[117][2] ) );
  DFE1 \FIFO_reg[117][1]  ( .D(n679), .E(N1333), .C(inClock), .Q(
        \FIFO[117][1] ) );
  DFE1 \FIFO_reg[117][0]  ( .D(n679), .E(N1334), .C(inClock), .Q(
        \FIFO[117][0] ) );
  DFE1 \FIFO_reg[116][3]  ( .D(n679), .E(N1335), .C(inClock), .Q(
        \FIFO[116][3] ) );
  DFE1 \FIFO_reg[116][2]  ( .D(n679), .E(N1336), .C(inClock), .Q(
        \FIFO[116][2] ) );
  DFE1 \FIFO_reg[116][1]  ( .D(n679), .E(N1337), .C(inClock), .Q(
        \FIFO[116][1] ) );
  DFE1 \FIFO_reg[116][0]  ( .D(n679), .E(N1338), .C(inClock), .Q(
        \FIFO[116][0] ) );
  DFE1 \FIFO_reg[115][3]  ( .D(n680), .E(N1339), .C(inClock), .Q(
        \FIFO[115][3] ) );
  DFE1 \FIFO_reg[115][2]  ( .D(n680), .E(N1340), .C(inClock), .Q(
        \FIFO[115][2] ) );
  DFE1 \FIFO_reg[115][1]  ( .D(n680), .E(N1341), .C(inClock), .Q(
        \FIFO[115][1] ) );
  DFE1 \FIFO_reg[115][0]  ( .D(n680), .E(N1342), .C(inClock), .Q(
        \FIFO[115][0] ) );
  DFE1 \FIFO_reg[113][3]  ( .D(n681), .E(N1347), .C(inClock), .Q(
        \FIFO[113][3] ) );
  DFE1 \FIFO_reg[113][2]  ( .D(n681), .E(N1348), .C(inClock), .Q(
        \FIFO[113][2] ) );
  DFE1 \FIFO_reg[113][1]  ( .D(n681), .E(N1349), .C(inClock), .Q(
        \FIFO[113][1] ) );
  DFE1 \FIFO_reg[113][0]  ( .D(n681), .E(N1350), .C(inClock), .Q(
        \FIFO[113][0] ) );
  DFE1 \FIFO_reg[112][3]  ( .D(n681), .E(N1351), .C(inClock), .Q(
        \FIFO[112][3] ) );
  DFE1 \FIFO_reg[112][2]  ( .D(n681), .E(N1352), .C(inClock), .Q(
        \FIFO[112][2] ) );
  DFE1 \FIFO_reg[112][1]  ( .D(n681), .E(N1353), .C(inClock), .Q(
        \FIFO[112][1] ) );
  DFE1 \FIFO_reg[112][0]  ( .D(n681), .E(N1354), .C(inClock), .Q(
        \FIFO[112][0] ) );
  DFE1 \FIFO_reg[111][3]  ( .D(n682), .E(N1355), .C(inClock), .Q(
        \FIFO[111][3] ) );
  DFE1 \FIFO_reg[111][2]  ( .D(n682), .E(N1356), .C(inClock), .Q(
        \FIFO[111][2] ) );
  DFE1 \FIFO_reg[111][1]  ( .D(n682), .E(N1357), .C(inClock), .Q(
        \FIFO[111][1] ) );
  DFE1 \FIFO_reg[111][0]  ( .D(n682), .E(N1358), .C(inClock), .Q(
        \FIFO[111][0] ) );
  DFE1 \FIFO_reg[107][3]  ( .D(n684), .E(N1371), .C(inClock), .Q(
        \FIFO[107][3] ) );
  DFE1 \FIFO_reg[107][2]  ( .D(n684), .E(N1372), .C(inClock), .Q(
        \FIFO[107][2] ) );
  DFE1 \FIFO_reg[107][1]  ( .D(n684), .E(N1373), .C(inClock), .Q(
        \FIFO[107][1] ) );
  DFE1 \FIFO_reg[107][0]  ( .D(n684), .E(N1374), .C(inClock), .Q(
        \FIFO[107][0] ) );
  DFE1 \FIFO_reg[105][3]  ( .D(n685), .E(N1379), .C(inClock), .Q(
        \FIFO[105][3] ) );
  DFE1 \FIFO_reg[105][2]  ( .D(n685), .E(N1380), .C(inClock), .Q(
        \FIFO[105][2] ) );
  DFE1 \FIFO_reg[105][1]  ( .D(n685), .E(N1381), .C(inClock), .Q(
        \FIFO[105][1] ) );
  DFE1 \FIFO_reg[105][0]  ( .D(n685), .E(N1382), .C(inClock), .Q(
        \FIFO[105][0] ) );
  DFE1 \FIFO_reg[104][3]  ( .D(n685), .E(N1383), .C(inClock), .Q(
        \FIFO[104][3] ) );
  DFE1 \FIFO_reg[104][2]  ( .D(n685), .E(N1384), .C(inClock), .Q(
        \FIFO[104][2] ) );
  DFE1 \FIFO_reg[104][1]  ( .D(n685), .E(N1385), .C(inClock), .Q(
        \FIFO[104][1] ) );
  DFE1 \FIFO_reg[104][0]  ( .D(n685), .E(N1386), .C(inClock), .Q(
        \FIFO[104][0] ) );
  DFE1 \FIFO_reg[103][3]  ( .D(n686), .E(N1387), .C(inClock), .Q(
        \FIFO[103][3] ) );
  DFE1 \FIFO_reg[103][2]  ( .D(n686), .E(N1388), .C(inClock), .Q(
        \FIFO[103][2] ) );
  DFE1 \FIFO_reg[103][1]  ( .D(n686), .E(N1389), .C(inClock), .Q(
        \FIFO[103][1] ) );
  DFE1 \FIFO_reg[103][0]  ( .D(n686), .E(N1390), .C(inClock), .Q(
        \FIFO[103][0] ) );
  DFE1 \FIFO_reg[99][3]  ( .D(n688), .E(N1403), .C(inClock), .Q(\FIFO[99][3] )
         );
  DFE1 \FIFO_reg[99][2]  ( .D(n688), .E(N1404), .C(inClock), .Q(\FIFO[99][2] )
         );
  DFE1 \FIFO_reg[99][1]  ( .D(n688), .E(N1405), .C(inClock), .Q(\FIFO[99][1] )
         );
  DFE1 \FIFO_reg[99][0]  ( .D(n688), .E(N1406), .C(inClock), .Q(\FIFO[99][0] )
         );
  DFE1 \FIFO_reg[97][3]  ( .D(n689), .E(N1411), .C(inClock), .Q(\FIFO[97][3] )
         );
  DFE1 \FIFO_reg[97][2]  ( .D(n689), .E(N1412), .C(inClock), .Q(\FIFO[97][2] )
         );
  DFE1 \FIFO_reg[97][1]  ( .D(n689), .E(N1413), .C(inClock), .Q(\FIFO[97][1] )
         );
  DFE1 \FIFO_reg[97][0]  ( .D(n689), .E(N1414), .C(inClock), .Q(\FIFO[97][0] )
         );
  DFE1 \FIFO_reg[96][3]  ( .D(n689), .E(N1415), .C(inClock), .Q(\FIFO[96][3] )
         );
  DFE1 \FIFO_reg[96][2]  ( .D(n689), .E(N1416), .C(inClock), .Q(\FIFO[96][2] )
         );
  DFE1 \FIFO_reg[96][1]  ( .D(n689), .E(N1417), .C(inClock), .Q(\FIFO[96][1] )
         );
  DFE1 \FIFO_reg[96][0]  ( .D(n689), .E(N1418), .C(inClock), .Q(\FIFO[96][0] )
         );
  DFE1 \FIFO_reg[91][3]  ( .D(n692), .E(N1435), .C(inClock), .Q(\FIFO[91][3] )
         );
  DFE1 \FIFO_reg[91][2]  ( .D(n692), .E(N1436), .C(inClock), .Q(\FIFO[91][2] )
         );
  DFE1 \FIFO_reg[91][1]  ( .D(n692), .E(N1437), .C(inClock), .Q(\FIFO[91][1] )
         );
  DFE1 \FIFO_reg[91][0]  ( .D(n692), .E(N1438), .C(inClock), .Q(\FIFO[91][0] )
         );
  DFE1 \FIFO_reg[83][3]  ( .D(n696), .E(N1467), .C(inClock), .Q(\FIFO[83][3] )
         );
  DFE1 \FIFO_reg[83][2]  ( .D(n696), .E(N1468), .C(inClock), .Q(\FIFO[83][2] )
         );
  DFE1 \FIFO_reg[83][1]  ( .D(n696), .E(N1469), .C(inClock), .Q(\FIFO[83][1] )
         );
  DFE1 \FIFO_reg[83][0]  ( .D(n696), .E(N1470), .C(inClock), .Q(\FIFO[83][0] )
         );
  DFE1 \FIFO_reg[79][3]  ( .D(n698), .E(N1483), .C(inClock), .Q(\FIFO[79][3] )
         );
  DFE1 \FIFO_reg[79][2]  ( .D(n698), .E(N1484), .C(inClock), .Q(\FIFO[79][2] )
         );
  DFE1 \FIFO_reg[79][1]  ( .D(n698), .E(N1485), .C(inClock), .Q(\FIFO[79][1] )
         );
  DFE1 \FIFO_reg[79][0]  ( .D(n698), .E(N1486), .C(inClock), .Q(\FIFO[79][0] )
         );
  DFE1 \FIFO_reg[75][3]  ( .D(n700), .E(N1499), .C(inClock), .Q(\FIFO[75][3] )
         );
  DFE1 \FIFO_reg[75][2]  ( .D(n700), .E(N1500), .C(inClock), .Q(\FIFO[75][2] )
         );
  DFE1 \FIFO_reg[75][1]  ( .D(n700), .E(N1501), .C(inClock), .Q(\FIFO[75][1] )
         );
  DFE1 \FIFO_reg[75][0]  ( .D(n700), .E(N1502), .C(inClock), .Q(\FIFO[75][0] )
         );
  DFE1 \FIFO_reg[73][3]  ( .D(n701), .E(N1507), .C(inClock), .Q(\FIFO[73][3] )
         );
  DFE1 \FIFO_reg[73][2]  ( .D(n701), .E(N1508), .C(inClock), .Q(\FIFO[73][2] )
         );
  DFE1 \FIFO_reg[73][1]  ( .D(n701), .E(N1509), .C(inClock), .Q(\FIFO[73][1] )
         );
  DFE1 \FIFO_reg[73][0]  ( .D(n701), .E(N1510), .C(inClock), .Q(\FIFO[73][0] )
         );
  DFE1 \FIFO_reg[72][3]  ( .D(n701), .E(N1511), .C(inClock), .Q(\FIFO[72][3] )
         );
  DFE1 \FIFO_reg[72][2]  ( .D(n701), .E(N1512), .C(inClock), .Q(\FIFO[72][2] )
         );
  DFE1 \FIFO_reg[72][1]  ( .D(n701), .E(N1513), .C(inClock), .Q(\FIFO[72][1] )
         );
  DFE1 \FIFO_reg[72][0]  ( .D(n701), .E(N1514), .C(inClock), .Q(\FIFO[72][0] )
         );
  DFE1 \FIFO_reg[71][3]  ( .D(n702), .E(N1515), .C(inClock), .Q(\FIFO[71][3] )
         );
  DFE1 \FIFO_reg[71][2]  ( .D(n702), .E(N1516), .C(inClock), .Q(\FIFO[71][2] )
         );
  DFE1 \FIFO_reg[71][1]  ( .D(n702), .E(N1517), .C(inClock), .Q(\FIFO[71][1] )
         );
  DFE1 \FIFO_reg[71][0]  ( .D(n702), .E(N1518), .C(inClock), .Q(\FIFO[71][0] )
         );
  DFE1 \FIFO_reg[67][3]  ( .D(n704), .E(N1531), .C(inClock), .Q(\FIFO[67][3] )
         );
  DFE1 \FIFO_reg[67][2]  ( .D(n704), .E(N1532), .C(inClock), .Q(\FIFO[67][2] )
         );
  DFE1 \FIFO_reg[67][1]  ( .D(n704), .E(N1533), .C(inClock), .Q(\FIFO[67][1] )
         );
  DFE1 \FIFO_reg[67][0]  ( .D(n704), .E(N1534), .C(inClock), .Q(\FIFO[67][0] )
         );
  DFE1 \FIFO_reg[65][3]  ( .D(n705), .E(N1539), .C(inClock), .Q(\FIFO[65][3] )
         );
  DFE1 \FIFO_reg[65][2]  ( .D(n705), .E(N1540), .C(inClock), .Q(\FIFO[65][2] )
         );
  DFE1 \FIFO_reg[65][1]  ( .D(n705), .E(N1541), .C(inClock), .Q(\FIFO[65][1] )
         );
  DFE1 \FIFO_reg[65][0]  ( .D(n705), .E(N1542), .C(inClock), .Q(\FIFO[65][0] )
         );
  DFE1 \FIFO_reg[64][3]  ( .D(n705), .E(N1543), .C(inClock), .Q(\FIFO[64][3] )
         );
  DFE1 \FIFO_reg[64][2]  ( .D(n705), .E(N1544), .C(inClock), .Q(\FIFO[64][2] )
         );
  DFE1 \FIFO_reg[64][1]  ( .D(n705), .E(N1545), .C(inClock), .Q(\FIFO[64][1] )
         );
  DFE1 \FIFO_reg[64][0]  ( .D(n705), .E(N1546), .C(inClock), .Q(\FIFO[64][0] )
         );
  DFE1 \FIFO_reg[59][3]  ( .D(n708), .E(N1563), .C(inClock), .Q(\FIFO[59][3] )
         );
  DFE1 \FIFO_reg[59][2]  ( .D(n708), .E(N1564), .C(inClock), .Q(\FIFO[59][2] )
         );
  DFE1 \FIFO_reg[59][1]  ( .D(n708), .E(N1565), .C(inClock), .Q(\FIFO[59][1] )
         );
  DFE1 \FIFO_reg[59][0]  ( .D(n708), .E(N1566), .C(inClock), .Q(\FIFO[59][0] )
         );
  DFE1 \FIFO_reg[51][3]  ( .D(n712), .E(N1595), .C(inClock), .Q(\FIFO[51][3] )
         );
  DFE1 \FIFO_reg[51][2]  ( .D(n712), .E(N1596), .C(inClock), .Q(\FIFO[51][2] )
         );
  DFE1 \FIFO_reg[51][1]  ( .D(n712), .E(N1597), .C(inClock), .Q(\FIFO[51][1] )
         );
  DFE1 \FIFO_reg[51][0]  ( .D(n712), .E(N1598), .C(inClock), .Q(\FIFO[51][0] )
         );
  DFE1 \i_FIFO_reg[6]  ( .D(N165), .E(n584), .C(inClock), .Q(i_FIFO[6]) );
  DFE1 \j_FIFO_reg[4]  ( .D(N226), .E(N213), .C(inClock), .Q(N43) );
  DFE1 \k_FIFO_reg[1]  ( .D(N192), .E(N183), .C(inClock), .Q(k_FIFO[1]), .QN(
        n569) );
  DFE1 \j_FIFO_reg[3]  ( .D(N225), .E(N213), .C(inClock), .Q(N42) );
  DFE1 \k_FIFO_reg[0]  ( .D(N191), .E(N183), .C(inClock), .Q(k_FIFO[0]), .QN(
        n547) );
  DFE1 \sigRDCOUNT_reg[6]  ( .D(n846), .E(N1287), .C(inClock), .Q(
        outReadCount[6]), .QN(n567) );
  DFE1 \i_FIFO_reg[2]  ( .D(N161), .E(n584), .C(inClock), .Q(i_FIFO[2]), .QN(
        n543) );
  DFE1 \i_FIFO_reg[3]  ( .D(N162), .E(n584), .C(inClock), .Q(i_FIFO[3]), .QN(
        n557) );
  DFE1 \sigWRCOUNT_reg[7]  ( .D(n839), .E(N1286), .C(inClock), .Q(
        outWriteCount[7]), .QN(n571) );
  DFE1 \sigWRCOUNT_reg[6]  ( .D(n838), .E(N1286), .C(inClock), .Q(
        outWriteCount[6]), .QN(n564) );
  DFE1 \i_FIFO_reg[4]  ( .D(N163), .E(n584), .C(inClock), .Q(i_FIFO[4]), .QN(
        n544) );
  DFE1 \i_FIFO_reg[5]  ( .D(N164), .E(n584), .C(inClock), .Q(i_FIFO[5]), .QN(
        n563) );
  DFE1 \j_FIFO_reg[1]  ( .D(N223), .E(N213), .C(inClock), .Q(N40) );
  DFE1 \j_FIFO_reg[2]  ( .D(N224), .E(N213), .C(inClock), .Q(N41), .QN(n545)
         );
  DFE1 \sigRDCOUNT_reg[4]  ( .D(n844), .E(N1287), .C(inClock), .Q(
        outReadCount[4]), .QN(n554) );
  DFE1 \sigRDCOUNT_reg[5]  ( .D(n845), .E(N1287), .C(inClock), .Q(
        outReadCount[5]), .QN(n570) );
  DFE1 \i_FIFO_reg[1]  ( .D(N160), .E(n584), .C(inClock), .Q(i_FIFO[1]), .QN(
        n556) );
  DFE1 \j_FIFO_reg[0]  ( .D(N222), .E(N213), .C(inClock), .Q(N39) );
  DFE1 \sigWRCOUNT_reg[5]  ( .D(n837), .E(N1286), .C(inClock), .Q(
        outWriteCount[5]), .QN(n566) );
  DFE1 \i_FIFO_reg[0]  ( .D(N159), .E(n584), .C(inClock), .Q(i_FIFO[0]), .QN(
        n542) );
  DFE1 \sigWRCOUNT_reg[4]  ( .D(n836), .E(N1286), .C(inClock), .Q(
        outWriteCount[4]), .QN(n568) );
  DFE1 \sigRDCOUNT_reg[1]  ( .D(n841), .E(N1287), .C(inClock), .Q(
        outReadCount[1]), .QN(n549) );
  DFE1 \sigRDCOUNT_reg[2]  ( .D(n842), .E(N1287), .C(inClock), .Q(
        outReadCount[2]), .QN(n551) );
  DFE1 \sigRDCOUNT_reg[3]  ( .D(n843), .E(N1287), .C(inClock), .Q(
        outReadCount[3]), .QN(n555) );
  DFE1 \sigWRCOUNT_reg[2]  ( .D(n834), .E(N1286), .C(inClock), .Q(
        outWriteCount[2]), .QN(n553) );
  DFE1 \sigWRCOUNT_reg[3]  ( .D(n835), .E(N1286), .C(inClock), .Q(
        outWriteCount[3]), .QN(n565) );
  DFE1 \sigWRCOUNT_reg[1]  ( .D(n833), .E(N1286), .C(inClock), .Q(
        outWriteCount[1]) );
  DFE1 \sigRDCOUNT_reg[0]  ( .D(n840), .E(N1287), .C(inClock), .Q(
        outReadCount[0]), .QN(n550) );
  DFE1 \sigWRCOUNT_reg[0]  ( .D(n832), .E(N1286), .C(inClock), .Q(
        outWriteCount[0]), .QN(n552) );
  IMUX40 U1080 ( .A(n535), .B(n525), .C(n530), .D(n520), .S0(n579), .S1(n580), 
        .Q(n540) );
  IMUX40 U1046 ( .A(n493), .B(n483), .C(n488), .D(n478), .S0(n579), .S1(n580), 
        .Q(n498) );
  IMUX40 U1012 ( .A(n451), .B(n441), .C(n446), .D(n436), .S0(n579), .S1(n580), 
        .Q(n456) );
  IMUX40 U978 ( .A(n409), .B(n399), .C(n404), .D(n394), .S0(n579), .S1(n580), 
        .Q(n414) );
  IMUX40 U951 ( .A(\FIFO[100][0] ), .B(\FIFO[101][0] ), .C(\FIFO[102][0] ), 
        .D(\FIFO[103][0] ), .S0(n829), .S1(n817), .Q(n382) );
  IMUX40 U947 ( .A(\FIFO[116][0] ), .B(\FIFO[117][0] ), .C(\FIFO[118][0] ), 
        .D(\FIFO[119][0] ), .S0(n828), .S1(n818), .Q(n377) );
  IMUX40 U1057 ( .A(\FIFO[84][3] ), .B(\FIFO[85][3] ), .C(\FIFO[86][3] ), .D(
        \FIFO[87][3] ), .S0(n826), .S1(n819), .Q(n513) );
  IMUX40 U1053 ( .A(\FIFO[100][3] ), .B(\FIFO[101][3] ), .C(\FIFO[102][3] ), 
        .D(\FIFO[103][3] ), .S0(n820), .S1(n819), .Q(n508) );
  IMUX40 U1061 ( .A(\FIFO[68][3] ), .B(\FIFO[69][3] ), .C(\FIFO[70][3] ), .D(
        \FIFO[71][3] ), .S0(n826), .S1(n819), .Q(n518) );
  IMUX40 U1023 ( .A(\FIFO[84][2] ), .B(\FIFO[85][2] ), .C(\FIFO[86][2] ), .D(
        \FIFO[87][2] ), .S0(n822), .S1(n816), .Q(n471) );
  IMUX40 U1019 ( .A(\FIFO[100][2] ), .B(\FIFO[101][2] ), .C(\FIFO[102][2] ), 
        .D(\FIFO[103][2] ), .S0(n822), .S1(n817), .Q(n466) );
  IMUX40 U1027 ( .A(\FIFO[68][2] ), .B(\FIFO[69][2] ), .C(\FIFO[70][2] ), .D(
        \FIFO[71][2] ), .S0(n830), .S1(n816), .Q(n476) );
  IMUX40 U989 ( .A(\FIFO[84][1] ), .B(\FIFO[85][1] ), .C(\FIFO[86][1] ), .D(
        \FIFO[87][1] ), .S0(n830), .S1(n816), .Q(n429) );
  IMUX40 U985 ( .A(\FIFO[100][1] ), .B(\FIFO[101][1] ), .C(\FIFO[102][1] ), 
        .D(\FIFO[103][1] ), .S0(n830), .S1(n815), .Q(n424) );
  IMUX40 U993 ( .A(\FIFO[68][1] ), .B(\FIFO[69][1] ), .C(\FIFO[70][1] ), .D(
        \FIFO[71][1] ), .S0(n829), .S1(n816), .Q(n434) );
  IMUX40 U955 ( .A(\FIFO[84][0] ), .B(\FIFO[85][0] ), .C(\FIFO[86][0] ), .D(
        \FIFO[87][0] ), .S0(n822), .S1(n819), .Q(n387) );
  IMUX40 U1075 ( .A(\FIFO[16][3] ), .B(\FIFO[17][3] ), .C(\FIFO[18][3] ), .D(
        \FIFO[19][3] ), .S0(n825), .S1(n818), .Q(n531) );
  IMUX40 U1073 ( .A(\FIFO[24][3] ), .B(\FIFO[25][3] ), .C(\FIFO[26][3] ), .D(
        \FIFO[27][3] ), .S0(n825), .S1(n817), .Q(n532) );
  IMUX40 U1074 ( .A(\FIFO[20][3] ), .B(\FIFO[21][3] ), .C(\FIFO[22][3] ), .D(
        \FIFO[23][3] ), .S0(n825), .S1(n815), .Q(n533) );
  IMUX40 U942 ( .A(n531), .B(n532), .C(n533), .D(n534), .S0(n813), .S1(n581), 
        .Q(n530) );
  IMUX40 U1041 ( .A(\FIFO[16][2] ), .B(\FIFO[17][2] ), .C(\FIFO[18][2] ), .D(
        \FIFO[19][2] ), .S0(n820), .S1(n818), .Q(n489) );
  IMUX40 U1039 ( .A(\FIFO[24][2] ), .B(\FIFO[25][2] ), .C(\FIFO[26][2] ), .D(
        \FIFO[27][2] ), .S0(n827), .S1(n818), .Q(n490) );
  IMUX40 U1040 ( .A(\FIFO[20][2] ), .B(\FIFO[21][2] ), .C(\FIFO[22][2] ), .D(
        \FIFO[23][2] ), .S0(n827), .S1(n818), .Q(n491) );
  IMUX40 U933 ( .A(n489), .B(n490), .C(n491), .D(n492), .S0(n814), .S1(n581), 
        .Q(n488) );
  IMUX40 U1007 ( .A(\FIFO[16][1] ), .B(\FIFO[17][1] ), .C(\FIFO[18][1] ), .D(
        \FIFO[19][1] ), .S0(n828), .S1(n817), .Q(n447) );
  IMUX40 U1005 ( .A(\FIFO[24][1] ), .B(\FIFO[25][1] ), .C(\FIFO[26][1] ), .D(
        \FIFO[27][1] ), .S0(n828), .S1(n817), .Q(n448) );
  IMUX40 U1006 ( .A(\FIFO[20][1] ), .B(\FIFO[21][1] ), .C(\FIFO[22][1] ), .D(
        \FIFO[23][1] ), .S0(n828), .S1(n817), .Q(n449) );
  IMUX40 U924 ( .A(n447), .B(n448), .C(n449), .D(n450), .S0(n813), .S1(n581), 
        .Q(n446) );
  IMUX40 U973 ( .A(\FIFO[16][0] ), .B(\FIFO[17][0] ), .C(\FIFO[18][0] ), .D(
        \FIFO[19][0] ), .S0(n824), .S1(n815), .Q(n405) );
  IMUX40 U971 ( .A(\FIFO[24][0] ), .B(\FIFO[25][0] ), .C(\FIFO[26][0] ), .D(
        \FIFO[27][0] ), .S0(n824), .S1(n815), .Q(n406) );
  IMUX40 U972 ( .A(\FIFO[20][0] ), .B(\FIFO[21][0] ), .C(\FIFO[22][0] ), .D(
        \FIFO[23][0] ), .S0(n824), .S1(n819), .Q(n407) );
  IMUX40 U915 ( .A(n405), .B(n406), .C(n407), .D(n408), .S0(n814), .S1(n581), 
        .Q(n404) );
  IMUX40 U949 ( .A(\FIFO[108][0] ), .B(\FIFO[109][0] ), .C(\FIFO[110][0] ), 
        .D(\FIFO[111][0] ), .S0(n827), .S1(n816), .Q(n383) );
  IMUX40 U950 ( .A(\FIFO[104][0] ), .B(\FIFO[105][0] ), .C(\FIFO[106][0] ), 
        .D(\FIFO[107][0] ), .S0(n826), .S1(n816), .Q(n381) );
  IMUX40 U952 ( .A(\FIFO[96][0] ), .B(\FIFO[97][0] ), .C(\FIFO[98][0] ), .D(
        \FIFO[99][0] ), .S0(n830), .S1(N40), .Q(n380) );
  IMUX40 U945 ( .A(\FIFO[124][0] ), .B(\FIFO[125][0] ), .C(\FIFO[126][0] ), 
        .D(\FIFO[127][0] ), .S0(n825), .S1(n818), .Q(n378) );
  IMUX40 U946 ( .A(\FIFO[120][0] ), .B(\FIFO[121][0] ), .C(\FIFO[122][0] ), 
        .D(\FIFO[123][0] ), .S0(n820), .S1(n817), .Q(n376) );
  IMUX40 U948 ( .A(\FIFO[112][0] ), .B(\FIFO[113][0] ), .C(\FIFO[114][0] ), 
        .D(\FIFO[115][0] ), .S0(n824), .S1(N40), .Q(n375) );
  IMUX40 U1072 ( .A(\FIFO[28][3] ), .B(\FIFO[29][3] ), .C(\FIFO[30][3] ), .D(
        \FIFO[31][3] ), .S0(n825), .S1(n818), .Q(n534) );
  IMUX40 U1067 ( .A(\FIFO[48][3] ), .B(\FIFO[49][3] ), .C(\FIFO[50][3] ), .D(
        \FIFO[51][3] ), .S0(n825), .S1(n819), .Q(n521) );
  IMUX40 U1068 ( .A(\FIFO[44][3] ), .B(\FIFO[45][3] ), .C(\FIFO[46][3] ), .D(
        \FIFO[47][3] ), .S0(n825), .S1(n816), .Q(n529) );
  IMUX40 U1076 ( .A(\FIFO[12][3] ), .B(\FIFO[13][3] ), .C(\FIFO[14][3] ), .D(
        \FIFO[15][3] ), .S0(n825), .S1(n819), .Q(n539) );
  IMUX40 U1055 ( .A(\FIFO[92][3] ), .B(\FIFO[93][3] ), .C(\FIFO[94][3] ), .D(
        \FIFO[95][3] ), .S0(n826), .S1(n819), .Q(n514) );
  IMUX40 U1056 ( .A(\FIFO[88][3] ), .B(\FIFO[89][3] ), .C(\FIFO[90][3] ), .D(
        \FIFO[91][3] ), .S0(n826), .S1(n818), .Q(n512) );
  IMUX40 U1058 ( .A(\FIFO[80][3] ), .B(\FIFO[81][3] ), .C(\FIFO[82][3] ), .D(
        \FIFO[83][3] ), .S0(n826), .S1(n816), .Q(n511) );
  IMUX40 U1051 ( .A(\FIFO[108][3] ), .B(\FIFO[109][3] ), .C(\FIFO[110][3] ), 
        .D(\FIFO[111][3] ), .S0(n820), .S1(n819), .Q(n509) );
  IMUX40 U1052 ( .A(\FIFO[104][3] ), .B(\FIFO[105][3] ), .C(\FIFO[106][3] ), 
        .D(\FIFO[107][3] ), .S0(n823), .S1(n819), .Q(n507) );
  IMUX40 U1054 ( .A(\FIFO[96][3] ), .B(\FIFO[97][3] ), .C(\FIFO[98][3] ), .D(
        \FIFO[99][3] ), .S0(n826), .S1(n818), .Q(n506) );
  IMUX40 U1059 ( .A(\FIFO[76][3] ), .B(\FIFO[77][3] ), .C(\FIFO[78][3] ), .D(
        \FIFO[79][3] ), .S0(n826), .S1(n819), .Q(n519) );
  IMUX40 U1060 ( .A(\FIFO[72][3] ), .B(\FIFO[73][3] ), .C(\FIFO[74][3] ), .D(
        \FIFO[75][3] ), .S0(n826), .S1(n819), .Q(n517) );
  IMUX40 U1062 ( .A(\FIFO[64][3] ), .B(\FIFO[65][3] ), .C(\FIFO[66][3] ), .D(
        \FIFO[67][3] ), .S0(n826), .S1(n816), .Q(n516) );
  IMUX40 U1050 ( .A(\FIFO[112][3] ), .B(\FIFO[113][3] ), .C(\FIFO[114][3] ), 
        .D(\FIFO[115][3] ), .S0(n822), .S1(n815), .Q(n501) );
  IMUX40 U1038 ( .A(\FIFO[28][2] ), .B(\FIFO[29][2] ), .C(\FIFO[30][2] ), .D(
        \FIFO[31][2] ), .S0(n827), .S1(n818), .Q(n492) );
  IMUX40 U1033 ( .A(\FIFO[48][2] ), .B(\FIFO[49][2] ), .C(\FIFO[50][2] ), .D(
        \FIFO[51][2] ), .S0(n827), .S1(n818), .Q(n479) );
  IMUX40 U1034 ( .A(\FIFO[44][2] ), .B(\FIFO[45][2] ), .C(\FIFO[46][2] ), .D(
        \FIFO[47][2] ), .S0(n827), .S1(n818), .Q(n487) );
  IMUX40 U1042 ( .A(\FIFO[12][2] ), .B(\FIFO[13][2] ), .C(\FIFO[14][2] ), .D(
        \FIFO[15][2] ), .S0(n821), .S1(n818), .Q(n497) );
  IMUX40 U1021 ( .A(\FIFO[92][2] ), .B(\FIFO[93][2] ), .C(\FIFO[94][2] ), .D(
        \FIFO[95][2] ), .S0(n821), .S1(n819), .Q(n472) );
  IMUX40 U1022 ( .A(\FIFO[88][2] ), .B(\FIFO[89][2] ), .C(\FIFO[90][2] ), .D(
        \FIFO[91][2] ), .S0(n821), .S1(n817), .Q(n470) );
  IMUX40 U1024 ( .A(\FIFO[80][2] ), .B(\FIFO[81][2] ), .C(\FIFO[82][2] ), .D(
        \FIFO[83][2] ), .S0(N39), .S1(n815), .Q(n469) );
  IMUX40 U1017 ( .A(\FIFO[108][2] ), .B(\FIFO[109][2] ), .C(\FIFO[110][2] ), 
        .D(\FIFO[111][2] ), .S0(n822), .S1(n819), .Q(n467) );
  IMUX40 U1018 ( .A(\FIFO[104][2] ), .B(\FIFO[105][2] ), .C(\FIFO[106][2] ), 
        .D(\FIFO[107][2] ), .S0(n820), .S1(n819), .Q(n465) );
  IMUX40 U1020 ( .A(\FIFO[96][2] ), .B(\FIFO[97][2] ), .C(\FIFO[98][2] ), .D(
        \FIFO[99][2] ), .S0(n820), .S1(n818), .Q(n464) );
  IMUX40 U1025 ( .A(\FIFO[76][2] ), .B(\FIFO[77][2] ), .C(\FIFO[78][2] ), .D(
        \FIFO[79][2] ), .S0(n824), .S1(n819), .Q(n477) );
  IMUX40 U1026 ( .A(\FIFO[72][2] ), .B(\FIFO[73][2] ), .C(\FIFO[74][2] ), .D(
        \FIFO[75][2] ), .S0(n823), .S1(n818), .Q(n475) );
  IMUX40 U1028 ( .A(\FIFO[64][2] ), .B(\FIFO[65][2] ), .C(\FIFO[66][2] ), .D(
        \FIFO[67][2] ), .S0(n827), .S1(n819), .Q(n474) );
  IMUX40 U1016 ( .A(\FIFO[112][2] ), .B(\FIFO[113][2] ), .C(\FIFO[114][2] ), 
        .D(\FIFO[115][2] ), .S0(n823), .S1(n817), .Q(n459) );
  IMUX40 U1004 ( .A(\FIFO[28][1] ), .B(\FIFO[29][1] ), .C(\FIFO[30][1] ), .D(
        \FIFO[31][1] ), .S0(n828), .S1(n817), .Q(n450) );
  IMUX40 U999 ( .A(\FIFO[48][1] ), .B(\FIFO[49][1] ), .C(\FIFO[50][1] ), .D(
        \FIFO[51][1] ), .S0(n829), .S1(n816), .Q(n437) );
  IMUX40 U1000 ( .A(\FIFO[44][1] ), .B(\FIFO[45][1] ), .C(\FIFO[46][1] ), .D(
        \FIFO[47][1] ), .S0(n829), .S1(n816), .Q(n445) );
  IMUX40 U1008 ( .A(\FIFO[12][1] ), .B(\FIFO[13][1] ), .C(\FIFO[14][1] ), .D(
        \FIFO[15][1] ), .S0(n828), .S1(n817), .Q(n455) );
  IMUX40 U987 ( .A(\FIFO[92][1] ), .B(\FIFO[93][1] ), .C(\FIFO[94][1] ), .D(
        \FIFO[95][1] ), .S0(n830), .S1(n816), .Q(n430) );
  IMUX40 U988 ( .A(\FIFO[88][1] ), .B(\FIFO[89][1] ), .C(\FIFO[90][1] ), .D(
        \FIFO[91][1] ), .S0(n830), .S1(n816), .Q(n428) );
  IMUX40 U990 ( .A(\FIFO[80][1] ), .B(\FIFO[81][1] ), .C(\FIFO[82][1] ), .D(
        \FIFO[83][1] ), .S0(n830), .S1(n816), .Q(n427) );
  IMUX40 U983 ( .A(\FIFO[108][1] ), .B(\FIFO[109][1] ), .C(\FIFO[110][1] ), 
        .D(\FIFO[111][1] ), .S0(n830), .S1(n817), .Q(n425) );
  IMUX40 U984 ( .A(\FIFO[104][1] ), .B(\FIFO[105][1] ), .C(\FIFO[106][1] ), 
        .D(\FIFO[107][1] ), .S0(n830), .S1(n817), .Q(n423) );
  IMUX40 U986 ( .A(\FIFO[96][1] ), .B(\FIFO[97][1] ), .C(\FIFO[98][1] ), .D(
        \FIFO[99][1] ), .S0(n830), .S1(n815), .Q(n422) );
  IMUX40 U991 ( .A(\FIFO[76][1] ), .B(\FIFO[77][1] ), .C(\FIFO[78][1] ), .D(
        \FIFO[79][1] ), .S0(n829), .S1(n816), .Q(n435) );
  IMUX40 U992 ( .A(\FIFO[72][1] ), .B(\FIFO[73][1] ), .C(\FIFO[74][1] ), .D(
        \FIFO[75][1] ), .S0(n829), .S1(n816), .Q(n433) );
  IMUX40 U994 ( .A(\FIFO[64][1] ), .B(\FIFO[65][1] ), .C(\FIFO[66][1] ), .D(
        \FIFO[67][1] ), .S0(n829), .S1(n816), .Q(n432) );
  IMUX40 U982 ( .A(\FIFO[112][1] ), .B(\FIFO[113][1] ), .C(\FIFO[114][1] ), 
        .D(\FIFO[115][1] ), .S0(n830), .S1(n817), .Q(n417) );
  IMUX40 U970 ( .A(\FIFO[28][0] ), .B(\FIFO[29][0] ), .C(\FIFO[30][0] ), .D(
        \FIFO[31][0] ), .S0(n824), .S1(n815), .Q(n408) );
  IMUX40 U965 ( .A(\FIFO[48][0] ), .B(\FIFO[49][0] ), .C(\FIFO[50][0] ), .D(
        \FIFO[51][0] ), .S0(n821), .S1(n815), .Q(n395) );
  IMUX40 U966 ( .A(\FIFO[44][0] ), .B(\FIFO[45][0] ), .C(\FIFO[46][0] ), .D(
        \FIFO[47][0] ), .S0(n824), .S1(n815), .Q(n403) );
  IMUX40 U974 ( .A(\FIFO[12][0] ), .B(\FIFO[13][0] ), .C(\FIFO[14][0] ), .D(
        \FIFO[15][0] ), .S0(n824), .S1(n816), .Q(n413) );
  IMUX40 U953 ( .A(\FIFO[92][0] ), .B(\FIFO[93][0] ), .C(\FIFO[94][0] ), .D(
        \FIFO[95][0] ), .S0(n829), .S1(n819), .Q(n388) );
  IMUX40 U954 ( .A(\FIFO[88][0] ), .B(\FIFO[89][0] ), .C(\FIFO[90][0] ), .D(
        \FIFO[91][0] ), .S0(n823), .S1(N40), .Q(n386) );
  IMUX40 U956 ( .A(\FIFO[80][0] ), .B(\FIFO[81][0] ), .C(\FIFO[82][0] ), .D(
        \FIFO[83][0] ), .S0(n822), .S1(N40), .Q(n385) );
  IMUX40 U960 ( .A(\FIFO[64][0] ), .B(\FIFO[65][0] ), .C(\FIFO[66][0] ), .D(
        \FIFO[67][0] ), .S0(n824), .S1(n815), .Q(n390) );
  IMUX40 U1079 ( .A(\FIFO[0][3] ), .B(\FIFO[1][3] ), .C(\FIFO[2][3] ), .D(
        \FIFO[3][3] ), .S0(n828), .S1(n819), .Q(n536) );
  IMUX40 U1077 ( .A(\FIFO[8][3] ), .B(\FIFO[9][3] ), .C(\FIFO[10][3] ), .D(
        \FIFO[11][3] ), .S0(n825), .S1(n819), .Q(n537) );
  IMUX40 U1078 ( .A(\FIFO[4][3] ), .B(\FIFO[5][3] ), .C(\FIFO[6][3] ), .D(
        \FIFO[7][3] ), .S0(n825), .S1(n819), .Q(n538) );
  IMUX40 U943 ( .A(n536), .B(n537), .C(n538), .D(n539), .S0(N42), .S1(n581), 
        .Q(n535) );
  IMUX40 U1065 ( .A(\FIFO[56][3] ), .B(\FIFO[57][3] ), .C(\FIFO[58][3] ), .D(
        \FIFO[59][3] ), .S0(n826), .S1(n819), .Q(n522) );
  IMUX40 U1064 ( .A(\FIFO[60][3] ), .B(\FIFO[61][3] ), .C(\FIFO[62][3] ), .D(
        \FIFO[63][3] ), .S0(n826), .S1(n818), .Q(n524) );
  IMUX40 U1066 ( .A(\FIFO[52][3] ), .B(\FIFO[53][3] ), .C(\FIFO[54][3] ), .D(
        \FIFO[55][3] ), .S0(n826), .S1(n817), .Q(n523) );
  IMUX40 U940 ( .A(n521), .B(n522), .C(n523), .D(n524), .S0(n814), .S1(N41), 
        .Q(n520) );
  IMUX40 U1071 ( .A(\FIFO[32][3] ), .B(\FIFO[33][3] ), .C(\FIFO[34][3] ), .D(
        \FIFO[35][3] ), .S0(n825), .S1(n816), .Q(n526) );
  IMUX40 U1069 ( .A(\FIFO[40][3] ), .B(\FIFO[41][3] ), .C(\FIFO[42][3] ), .D(
        \FIFO[43][3] ), .S0(n825), .S1(n815), .Q(n527) );
  IMUX40 U1070 ( .A(\FIFO[36][3] ), .B(\FIFO[37][3] ), .C(\FIFO[38][3] ), .D(
        \FIFO[39][3] ), .S0(n825), .S1(n816), .Q(n528) );
  IMUX40 U941 ( .A(n526), .B(n527), .C(n528), .D(n529), .S0(n813), .S1(N41), 
        .Q(n525) );
  IMUX40 U1048 ( .A(\FIFO[120][3] ), .B(\FIFO[121][3] ), .C(\FIFO[122][3] ), 
        .D(\FIFO[123][3] ), .S0(n820), .S1(n819), .Q(n502) );
  IMUX40 U1047 ( .A(\FIFO[124][3] ), .B(\FIFO[125][3] ), .C(\FIFO[126][3] ), 
        .D(\FIFO[127][3] ), .S0(n821), .S1(n819), .Q(n504) );
  IMUX40 U1049 ( .A(\FIFO[116][3] ), .B(\FIFO[117][3] ), .C(\FIFO[118][3] ), 
        .D(\FIFO[119][3] ), .S0(n829), .S1(n819), .Q(n503) );
  IMUX40 U936 ( .A(n501), .B(n502), .C(n503), .D(n504), .S0(n814), .S1(N41), 
        .Q(n500) );
  IMUX40 U1031 ( .A(\FIFO[56][2] ), .B(\FIFO[57][2] ), .C(\FIFO[58][2] ), .D(
        \FIFO[59][2] ), .S0(n827), .S1(n815), .Q(n480) );
  IMUX40 U1030 ( .A(\FIFO[60][2] ), .B(\FIFO[61][2] ), .C(\FIFO[62][2] ), .D(
        \FIFO[63][2] ), .S0(n827), .S1(n817), .Q(n482) );
  IMUX40 U1032 ( .A(\FIFO[52][2] ), .B(\FIFO[53][2] ), .C(\FIFO[54][2] ), .D(
        \FIFO[55][2] ), .S0(n827), .S1(n818), .Q(n481) );
  IMUX40 U931 ( .A(n479), .B(n480), .C(n481), .D(n482), .S0(n814), .S1(N41), 
        .Q(n478) );
  IMUX40 U1037 ( .A(\FIFO[32][2] ), .B(\FIFO[33][2] ), .C(\FIFO[34][2] ), .D(
        \FIFO[35][2] ), .S0(n827), .S1(n818), .Q(n484) );
  IMUX40 U1035 ( .A(\FIFO[40][2] ), .B(\FIFO[41][2] ), .C(\FIFO[42][2] ), .D(
        \FIFO[43][2] ), .S0(n827), .S1(n818), .Q(n485) );
  IMUX40 U1036 ( .A(\FIFO[36][2] ), .B(\FIFO[37][2] ), .C(\FIFO[38][2] ), .D(
        \FIFO[39][2] ), .S0(n827), .S1(n818), .Q(n486) );
  IMUX40 U932 ( .A(n484), .B(n485), .C(n486), .D(n487), .S0(n814), .S1(N41), 
        .Q(n483) );
  IMUX40 U1045 ( .A(\FIFO[0][2] ), .B(\FIFO[1][2] ), .C(\FIFO[2][2] ), .D(
        \FIFO[3][2] ), .S0(n821), .S1(n818), .Q(n494) );
  IMUX40 U1043 ( .A(\FIFO[8][2] ), .B(\FIFO[9][2] ), .C(\FIFO[10][2] ), .D(
        \FIFO[11][2] ), .S0(n823), .S1(n818), .Q(n495) );
  IMUX40 U1044 ( .A(\FIFO[4][2] ), .B(\FIFO[5][2] ), .C(\FIFO[6][2] ), .D(
        \FIFO[7][2] ), .S0(n824), .S1(n818), .Q(n496) );
  IMUX40 U934 ( .A(n494), .B(n495), .C(n496), .D(n497), .S0(N42), .S1(n581), 
        .Q(n493) );
  IMUX40 U1014 ( .A(\FIFO[120][2] ), .B(\FIFO[121][2] ), .C(\FIFO[122][2] ), 
        .D(\FIFO[123][2] ), .S0(n828), .S1(n817), .Q(n460) );
  IMUX40 U1013 ( .A(\FIFO[124][2] ), .B(\FIFO[125][2] ), .C(\FIFO[126][2] ), 
        .D(\FIFO[127][2] ), .S0(n828), .S1(n817), .Q(n462) );
  IMUX40 U1015 ( .A(\FIFO[116][2] ), .B(\FIFO[117][2] ), .C(\FIFO[118][2] ), 
        .D(\FIFO[119][2] ), .S0(n828), .S1(n817), .Q(n461) );
  IMUX40 U927 ( .A(n459), .B(n460), .C(n461), .D(n462), .S0(n813), .S1(n581), 
        .Q(n458) );
  IMUX40 U997 ( .A(\FIFO[56][1] ), .B(\FIFO[57][1] ), .C(\FIFO[58][1] ), .D(
        \FIFO[59][1] ), .S0(n829), .S1(n816), .Q(n438) );
  IMUX40 U996 ( .A(\FIFO[60][1] ), .B(\FIFO[61][1] ), .C(\FIFO[62][1] ), .D(
        \FIFO[63][1] ), .S0(n829), .S1(n816), .Q(n440) );
  IMUX40 U998 ( .A(\FIFO[52][1] ), .B(\FIFO[53][1] ), .C(\FIFO[54][1] ), .D(
        \FIFO[55][1] ), .S0(n829), .S1(n816), .Q(n439) );
  IMUX40 U922 ( .A(n437), .B(n438), .C(n439), .D(n440), .S0(n813), .S1(N41), 
        .Q(n436) );
  IMUX40 U1003 ( .A(\FIFO[32][1] ), .B(\FIFO[33][1] ), .C(\FIFO[34][1] ), .D(
        \FIFO[35][1] ), .S0(n829), .S1(n817), .Q(n442) );
  IMUX40 U1001 ( .A(\FIFO[40][1] ), .B(\FIFO[41][1] ), .C(\FIFO[42][1] ), .D(
        \FIFO[43][1] ), .S0(n829), .S1(n816), .Q(n443) );
  IMUX40 U1002 ( .A(\FIFO[36][1] ), .B(\FIFO[37][1] ), .C(\FIFO[38][1] ), .D(
        \FIFO[39][1] ), .S0(n829), .S1(n817), .Q(n444) );
  IMUX40 U923 ( .A(n442), .B(n443), .C(n444), .D(n445), .S0(n813), .S1(N41), 
        .Q(n441) );
  IMUX40 U1011 ( .A(\FIFO[0][1] ), .B(\FIFO[1][1] ), .C(\FIFO[2][1] ), .D(
        \FIFO[3][1] ), .S0(n828), .S1(n817), .Q(n452) );
  IMUX40 U1009 ( .A(\FIFO[8][1] ), .B(\FIFO[9][1] ), .C(\FIFO[10][1] ), .D(
        \FIFO[11][1] ), .S0(n828), .S1(n817), .Q(n453) );
  IMUX40 U1010 ( .A(\FIFO[4][1] ), .B(\FIFO[5][1] ), .C(\FIFO[6][1] ), .D(
        \FIFO[7][1] ), .S0(n828), .S1(n817), .Q(n454) );
  IMUX40 U925 ( .A(n452), .B(n453), .C(n454), .D(n455), .S0(n813), .S1(n581), 
        .Q(n451) );
  IMUX40 U980 ( .A(\FIFO[120][1] ), .B(\FIFO[121][1] ), .C(\FIFO[122][1] ), 
        .D(\FIFO[123][1] ), .S0(n830), .S1(n815), .Q(n418) );
  IMUX40 U979 ( .A(\FIFO[124][1] ), .B(\FIFO[125][1] ), .C(\FIFO[126][1] ), 
        .D(\FIFO[127][1] ), .S0(n830), .S1(n815), .Q(n420) );
  IMUX40 U981 ( .A(\FIFO[116][1] ), .B(\FIFO[117][1] ), .C(\FIFO[118][1] ), 
        .D(\FIFO[119][1] ), .S0(n830), .S1(n818), .Q(n419) );
  IMUX40 U918 ( .A(n417), .B(n418), .C(n419), .D(n420), .S0(n813), .S1(n581), 
        .Q(n416) );
  IMUX40 U963 ( .A(\FIFO[56][0] ), .B(\FIFO[57][0] ), .C(\FIFO[58][0] ), .D(
        \FIFO[59][0] ), .S0(n830), .S1(n815), .Q(n396) );
  IMUX40 U962 ( .A(\FIFO[60][0] ), .B(\FIFO[61][0] ), .C(\FIFO[62][0] ), .D(
        \FIFO[63][0] ), .S0(n824), .S1(n815), .Q(n398) );
  IMUX40 U964 ( .A(\FIFO[52][0] ), .B(\FIFO[53][0] ), .C(\FIFO[54][0] ), .D(
        \FIFO[55][0] ), .S0(n828), .S1(n815), .Q(n397) );
  IMUX40 U913 ( .A(n395), .B(n396), .C(n397), .D(n398), .S0(n814), .S1(N41), 
        .Q(n394) );
  IMUX40 U969 ( .A(\FIFO[32][0] ), .B(\FIFO[33][0] ), .C(\FIFO[34][0] ), .D(
        \FIFO[35][0] ), .S0(n824), .S1(n815), .Q(n400) );
  IMUX40 U967 ( .A(\FIFO[40][0] ), .B(\FIFO[41][0] ), .C(\FIFO[42][0] ), .D(
        \FIFO[43][0] ), .S0(n824), .S1(n815), .Q(n401) );
  IMUX40 U968 ( .A(\FIFO[36][0] ), .B(\FIFO[37][0] ), .C(\FIFO[38][0] ), .D(
        \FIFO[39][0] ), .S0(n824), .S1(n815), .Q(n402) );
  IMUX40 U914 ( .A(n400), .B(n401), .C(n402), .D(n403), .S0(n814), .S1(N41), 
        .Q(n399) );
  IMUX40 U977 ( .A(\FIFO[0][0] ), .B(\FIFO[1][0] ), .C(\FIFO[2][0] ), .D(
        \FIFO[3][0] ), .S0(n824), .S1(n818), .Q(n410) );
  IMUX40 U975 ( .A(\FIFO[8][0] ), .B(\FIFO[9][0] ), .C(\FIFO[10][0] ), .D(
        \FIFO[11][0] ), .S0(n824), .S1(n816), .Q(n411) );
  IMUX40 U976 ( .A(\FIFO[4][0] ), .B(\FIFO[5][0] ), .C(\FIFO[6][0] ), .D(
        \FIFO[7][0] ), .S0(n824), .S1(n817), .Q(n412) );
  IMUX40 U916 ( .A(n410), .B(n411), .C(n412), .D(n413), .S0(n814), .S1(n581), 
        .Q(n409) );
  IMUX40 U958 ( .A(\FIFO[72][0] ), .B(\FIFO[73][0] ), .C(\FIFO[74][0] ), .D(
        \FIFO[75][0] ), .S0(n827), .S1(n815), .Q(n391) );
  IMUX40 U957 ( .A(\FIFO[76][0] ), .B(\FIFO[77][0] ), .C(\FIFO[78][0] ), .D(
        \FIFO[79][0] ), .S0(n830), .S1(n815), .Q(n393) );
  IMUX40 U959 ( .A(\FIFO[68][0] ), .B(\FIFO[69][0] ), .C(\FIFO[70][0] ), .D(
        \FIFO[71][0] ), .S0(n824), .S1(n815), .Q(n392) );
  IMUX40 U912 ( .A(n390), .B(n391), .C(n392), .D(n393), .S0(n814), .S1(n581), 
        .Q(n389) );
  DFE1 \sigOutData_reg[3]  ( .D(N209), .E(N201), .C(inClock), .Q(outData[3])
         );
  DFE1 \sigOutData_reg[2]  ( .D(N208), .E(N201), .C(inClock), .Q(outData[2])
         );
  DFE1 \sigOutData_reg[1]  ( .D(N207), .E(N201), .C(inClock), .Q(outData[1])
         );
  DFE1 \sigOutData_reg[0]  ( .D(N206), .E(N201), .C(inClock), .Q(outData[0])
         );
  IMUX40 U939 ( .A(n516), .B(n517), .C(n518), .D(n519), .S0(N42), .S1(n581), 
        .Q(n515) );
  IMUX40 U937 ( .A(n506), .B(n507), .C(n508), .D(n509), .S0(N42), .S1(N41), 
        .Q(n505) );
  IMUX40 U938 ( .A(n511), .B(n512), .C(n513), .D(n514), .S0(N42), .S1(n581), 
        .Q(n510) );
  IMUX40 U1063 ( .A(n515), .B(n505), .C(n510), .D(n500), .S0(n579), .S1(n580), 
        .Q(n541) );
  IMUX40 U930 ( .A(n474), .B(n475), .C(n476), .D(n477), .S0(n813), .S1(n581), 
        .Q(n473) );
  IMUX40 U928 ( .A(n464), .B(n465), .C(n466), .D(n467), .S0(n813), .S1(N41), 
        .Q(n463) );
  IMUX40 U929 ( .A(n469), .B(n470), .C(n471), .D(n472), .S0(n813), .S1(n581), 
        .Q(n468) );
  IMUX40 U1029 ( .A(n473), .B(n463), .C(n468), .D(n458), .S0(n579), .S1(n580), 
        .Q(n499) );
  IMUX40 U921 ( .A(n432), .B(n433), .C(n434), .D(n435), .S0(n813), .S1(n581), 
        .Q(n431) );
  IMUX40 U919 ( .A(n422), .B(n423), .C(n424), .D(n425), .S0(n813), .S1(N41), 
        .Q(n421) );
  IMUX40 U920 ( .A(n427), .B(n428), .C(n429), .D(n430), .S0(n813), .S1(n581), 
        .Q(n426) );
  IMUX40 U995 ( .A(n431), .B(n421), .C(n426), .D(n416), .S0(n579), .S1(n580), 
        .Q(n457) );
  IMUX40 U911 ( .A(n385), .B(n386), .C(n387), .D(n388), .S0(n814), .S1(n581), 
        .Q(n384) );
  IMUX40 U909 ( .A(n375), .B(n376), .C(n377), .D(n378), .S0(n814), .S1(n581), 
        .Q(n374) );
  IMUX40 U910 ( .A(n380), .B(n381), .C(n382), .D(n383), .S0(n814), .S1(N41), 
        .Q(n379) );
  IMUX40 U961 ( .A(n389), .B(n379), .C(n384), .D(n374), .S0(n579), .S1(n580), 
        .Q(n415) );
  DFE1 sigWError_reg ( .D(N1277), .E(N1804), .C(inClock), .Q(outWriteError) );
  DFE1 sigRError_reg ( .D(N1276), .E(N1806), .C(inClock), .Q(outReadError) );
  NOR21 U1081 ( .A(n576), .B(n809), .Q(N165) );
  NOR21 U1082 ( .A(n577), .B(n807), .Q(N228) );
  MUX22 U1083 ( .A(n414), .B(n415), .S(N45), .Q(n559) );
  MUX22 U1084 ( .A(n456), .B(n457), .S(N45), .Q(n560) );
  MUX22 U1085 ( .A(n498), .B(n499), .S(N45), .Q(n561) );
  MUX22 U1086 ( .A(n540), .B(n541), .S(N45), .Q(n562) );
  BUF2 U1087 ( .A(n177), .Q(n603) );
  BUF2 U1088 ( .A(n177), .Q(n602) );
  NAND22 U1089 ( .A(n856), .B(n150), .Q(n180) );
  BUF2 U1090 ( .A(n171), .Q(n605) );
  BUF2 U1091 ( .A(n171), .Q(n604) );
  BUF2 U1092 ( .A(n169), .Q(n609) );
  BUF2 U1093 ( .A(n170), .Q(n606) );
  BUF2 U1094 ( .A(n851), .Q(n640) );
  BUF2 U1095 ( .A(n169), .Q(n610) );
  BUF2 U1096 ( .A(n169), .Q(n611) );
  BUF2 U1097 ( .A(n170), .Q(n607) );
  BUF2 U1098 ( .A(n170), .Q(n608) );
  BUF2 U1099 ( .A(n851), .Q(n639) );
  BUF2 U1100 ( .A(n851), .Q(n638) );
  BUF2 U1101 ( .A(n851), .Q(n637) );
  BUF2 U1102 ( .A(n851), .Q(n636) );
  BUF2 U1103 ( .A(n851), .Q(n635) );
  BUF2 U1104 ( .A(n851), .Q(n634) );
  BUF2 U1105 ( .A(n851), .Q(n633) );
  INV3 U1106 ( .A(n648), .Q(n647) );
  INV3 U1107 ( .A(n650), .Q(n649) );
  INV3 U1108 ( .A(n642), .Q(n641) );
  INV3 U1109 ( .A(n654), .Q(n653) );
  INV3 U1110 ( .A(n646), .Q(n645) );
  INV3 U1111 ( .A(n652), .Q(n651) );
  INV3 U1112 ( .A(n644), .Q(n643) );
  INV3 U1113 ( .A(n660), .Q(n659) );
  INV3 U1114 ( .A(n658), .Q(n657) );
  INV3 U1115 ( .A(n656), .Q(n655) );
  INV3 U1116 ( .A(n662), .Q(n661) );
  INV3 U1117 ( .A(n143), .Q(n863) );
  BUF2 U1118 ( .A(n168), .Q(n613) );
  BUF2 U1119 ( .A(n168), .Q(n612) );
  NAND22 U1120 ( .A(n856), .B(N198), .Q(n177) );
  BUF2 U1121 ( .A(n738), .Q(n737) );
  BUF2 U1122 ( .A(n738), .Q(n736) );
  BUF2 U1123 ( .A(n739), .Q(n735) );
  BUF2 U1124 ( .A(n739), .Q(n734) );
  BUF2 U1125 ( .A(n740), .Q(n733) );
  BUF2 U1126 ( .A(n740), .Q(n732) );
  BUF2 U1127 ( .A(n741), .Q(n731) );
  BUF2 U1128 ( .A(n741), .Q(n730) );
  BUF2 U1129 ( .A(n742), .Q(n729) );
  BUF2 U1130 ( .A(n742), .Q(n728) );
  BUF2 U1131 ( .A(n743), .Q(n727) );
  BUF2 U1132 ( .A(n743), .Q(n726) );
  BUF2 U1133 ( .A(n744), .Q(n725) );
  BUF2 U1134 ( .A(n744), .Q(n724) );
  BUF2 U1135 ( .A(n745), .Q(n723) );
  BUF2 U1136 ( .A(n745), .Q(n722) );
  BUF2 U1137 ( .A(n746), .Q(n721) );
  BUF2 U1138 ( .A(n746), .Q(n720) );
  BUF2 U1139 ( .A(n747), .Q(n719) );
  BUF2 U1140 ( .A(n747), .Q(n718) );
  BUF2 U1141 ( .A(n748), .Q(n717) );
  BUF2 U1142 ( .A(n748), .Q(n716) );
  BUF2 U1143 ( .A(n749), .Q(n715) );
  BUF2 U1144 ( .A(n749), .Q(n714) );
  BUF2 U1145 ( .A(n750), .Q(n713) );
  BUF2 U1146 ( .A(n750), .Q(n712) );
  BUF2 U1147 ( .A(n751), .Q(n711) );
  BUF2 U1148 ( .A(n751), .Q(n710) );
  BUF2 U1149 ( .A(n752), .Q(n709) );
  BUF2 U1150 ( .A(n752), .Q(n708) );
  BUF2 U1151 ( .A(n753), .Q(n707) );
  BUF2 U1152 ( .A(n753), .Q(n706) );
  BUF2 U1153 ( .A(n754), .Q(n705) );
  BUF2 U1154 ( .A(n754), .Q(n704) );
  BUF2 U1155 ( .A(n755), .Q(n703) );
  BUF2 U1156 ( .A(n755), .Q(n702) );
  BUF2 U1157 ( .A(n756), .Q(n701) );
  BUF2 U1158 ( .A(n756), .Q(n700) );
  BUF2 U1159 ( .A(n757), .Q(n699) );
  BUF2 U1160 ( .A(n757), .Q(n698) );
  BUF2 U1161 ( .A(n758), .Q(n697) );
  BUF2 U1162 ( .A(n758), .Q(n696) );
  BUF2 U1163 ( .A(n759), .Q(n695) );
  BUF2 U1164 ( .A(n759), .Q(n694) );
  BUF2 U1165 ( .A(n760), .Q(n693) );
  BUF2 U1166 ( .A(n760), .Q(n692) );
  BUF2 U1167 ( .A(n761), .Q(n691) );
  BUF2 U1168 ( .A(n761), .Q(n690) );
  BUF2 U1169 ( .A(n762), .Q(n689) );
  BUF2 U1170 ( .A(n762), .Q(n688) );
  BUF2 U1171 ( .A(n763), .Q(n687) );
  BUF2 U1172 ( .A(n763), .Q(n686) );
  BUF2 U1173 ( .A(n764), .Q(n685) );
  BUF2 U1174 ( .A(n764), .Q(n684) );
  BUF2 U1175 ( .A(n765), .Q(n683) );
  BUF2 U1176 ( .A(n765), .Q(n682) );
  BUF2 U1177 ( .A(n766), .Q(n681) );
  BUF2 U1178 ( .A(n766), .Q(n680) );
  BUF2 U1179 ( .A(n767), .Q(n679) );
  BUF2 U1180 ( .A(n767), .Q(n678) );
  BUF2 U1181 ( .A(n768), .Q(n677) );
  BUF2 U1182 ( .A(n768), .Q(n676) );
  BUF2 U1183 ( .A(n769), .Q(n675) );
  BUF2 U1184 ( .A(n769), .Q(n674) );
  NOR21 U1185 ( .A(n184), .B(n640), .Q(n150) );
  NAND22 U1186 ( .A(n856), .B(n145), .Q(n178) );
  NAND22 U1187 ( .A(n856), .B(n146), .Q(n179) );
  INV3 U1188 ( .A(N183), .Q(n851) );
  NAND22 U1189 ( .A(n175), .B(n145), .Q(n169) );
  NAND22 U1190 ( .A(n175), .B(n146), .Q(n170) );
  NAND22 U1191 ( .A(n175), .B(n150), .Q(n171) );
  BUF2 U1192 ( .A(n152), .Q(n628) );
  BUF2 U1193 ( .A(n152), .Q(n627) );
  BUF2 U1194 ( .A(n153), .Q(n626) );
  BUF2 U1195 ( .A(n153), .Q(n625) );
  BUF2 U1196 ( .A(n164), .Q(n617) );
  BUF2 U1197 ( .A(n164), .Q(n616) );
  BUF2 U1198 ( .A(n154), .Q(n624) );
  BUF2 U1199 ( .A(n154), .Q(n623) );
  BUF2 U1200 ( .A(n165), .Q(n615) );
  BUF2 U1201 ( .A(n165), .Q(n614) );
  BUF2 U1202 ( .A(n163), .Q(n618) );
  NOR21 U1203 ( .A(n880), .B(n807), .Q(N227) );
  INV3 U1204 ( .A(N220), .Q(n880) );
  NOR21 U1205 ( .A(n881), .B(n807), .Q(N226) );
  INV3 U1206 ( .A(N219), .Q(n881) );
  BUF2 U1207 ( .A(n163), .Q(n619) );
  BUF2 U1208 ( .A(n163), .Q(n620) );
  NOR21 U1209 ( .A(n118), .B(n807), .Q(n116) );
  NAND22 U1210 ( .A(n358), .B(n328), .Q(n143) );
  NAND22 U1211 ( .A(n358), .B(n328), .Q(n586) );
  NAND22 U1212 ( .A(n358), .B(n328), .Q(n585) );
  INV3 U1213 ( .A(n198), .Q(n856) );
  NOR21 U1214 ( .A(n198), .B(n184), .Q(n186) );
  INV3 U1215 ( .A(n142), .Q(n865) );
  INV3 U1216 ( .A(n140), .Q(n866) );
  INV3 U1217 ( .A(n141), .Q(n862) );
  INV3 U1218 ( .A(n131), .Q(n656) );
  INV3 U1219 ( .A(n135), .Q(n648) );
  INV3 U1220 ( .A(n139), .Q(n864) );
  INV3 U1221 ( .A(n130), .Q(n658) );
  INV3 U1222 ( .A(n124), .Q(n662) );
  INV3 U1223 ( .A(n129), .Q(n660) );
  INV3 U1224 ( .A(n134), .Q(n650) );
  INV3 U1225 ( .A(n138), .Q(n642) );
  INV3 U1226 ( .A(n132), .Q(n654) );
  INV3 U1227 ( .A(n136), .Q(n646) );
  INV3 U1228 ( .A(n133), .Q(n652) );
  INV3 U1229 ( .A(n137), .Q(n644) );
  BUF2 U1230 ( .A(n151), .Q(n630) );
  BUF2 U1231 ( .A(n151), .Q(n629) );
  BUF2 U1232 ( .A(n162), .Q(n622) );
  BUF2 U1233 ( .A(n162), .Q(n621) );
  BUF2 U1234 ( .A(n202), .Q(n601) );
  BUF2 U1235 ( .A(n202), .Q(n600) );
  BUF2 U1236 ( .A(n255), .Q(n597) );
  BUF2 U1237 ( .A(n255), .Q(n596) );
  BUF2 U1238 ( .A(n308), .Q(n590) );
  BUF2 U1239 ( .A(n308), .Q(n589) );
  BUF2 U1240 ( .A(n125), .Q(n631) );
  BUF2 U1241 ( .A(n125), .Q(n632) );
  NAND22 U1242 ( .A(n175), .B(N198), .Q(n168) );
  INV3 U1243 ( .A(n598), .Q(n599) );
  INV3 U1244 ( .A(n587), .Q(n588) );
  INV3 U1245 ( .A(n118), .Q(n875) );
  INV3 U1246 ( .A(n117), .Q(n831) );
  NOR21 U1247 ( .A(n882), .B(n807), .Q(N225) );
  INV3 U1248 ( .A(N218), .Q(n882) );
  NOR21 U1249 ( .A(n883), .B(n807), .Q(N224) );
  INV3 U1250 ( .A(N217), .Q(n883) );
  NOR21 U1251 ( .A(n884), .B(n807), .Q(N223) );
  INV3 U1252 ( .A(N216), .Q(n884) );
  NOR21 U1253 ( .A(n639), .B(n187), .Q(N1497) );
  AOI211 U1254 ( .A(n188), .B(n866), .C(n808), .Q(n187) );
  NOR21 U1255 ( .A(n639), .B(n189), .Q(N1496) );
  AOI211 U1256 ( .A(n190), .B(n866), .C(n808), .Q(n189) );
  NOR21 U1257 ( .A(n639), .B(n191), .Q(N1495) );
  AOI211 U1258 ( .A(n186), .B(n866), .C(n808), .Q(n191) );
  NOR21 U1259 ( .A(n639), .B(n192), .Q(N1493) );
  AOI211 U1260 ( .A(n188), .B(n862), .C(n808), .Q(n192) );
  NOR21 U1261 ( .A(n639), .B(n193), .Q(N1492) );
  AOI211 U1262 ( .A(n190), .B(n862), .C(n808), .Q(n193) );
  NOR21 U1263 ( .A(n639), .B(n194), .Q(N1491) );
  AOI211 U1264 ( .A(n186), .B(n862), .C(n808), .Q(n194) );
  NOR21 U1265 ( .A(n639), .B(n195), .Q(N1489) );
  AOI211 U1266 ( .A(n188), .B(n865), .C(n808), .Q(n195) );
  NOR21 U1267 ( .A(n639), .B(n196), .Q(N1488) );
  AOI211 U1268 ( .A(n190), .B(n865), .C(n808), .Q(n196) );
  NOR21 U1269 ( .A(n639), .B(n197), .Q(N1487) );
  AOI211 U1270 ( .A(n186), .B(n865), .C(n808), .Q(n197) );
  NOR21 U1271 ( .A(n639), .B(n199), .Q(N1485) );
  AOI211 U1272 ( .A(n188), .B(n863), .C(n808), .Q(n199) );
  NOR21 U1273 ( .A(n639), .B(n200), .Q(N1484) );
  AOI211 U1274 ( .A(n190), .B(n863), .C(n808), .Q(n200) );
  NOR21 U1275 ( .A(n639), .B(n201), .Q(N1483) );
  AOI211 U1276 ( .A(n186), .B(n863), .C(n808), .Q(n201) );
  NOR21 U1277 ( .A(n639), .B(n203), .Q(N1481) );
  AOI211 U1278 ( .A(n599), .B(n662), .C(n808), .Q(n203) );
  NOR21 U1279 ( .A(n638), .B(n205), .Q(N1480) );
  AOI211 U1280 ( .A(n206), .B(n662), .C(n808), .Q(n205) );
  NOR21 U1281 ( .A(n638), .B(n207), .Q(N1479) );
  AOI211 U1282 ( .A(n208), .B(n662), .C(n807), .Q(n207) );
  NOR21 U1283 ( .A(n638), .B(n209), .Q(N1477) );
  AOI211 U1284 ( .A(n204), .B(n660), .C(n808), .Q(n209) );
  NOR21 U1285 ( .A(n638), .B(n210), .Q(N1476) );
  AOI211 U1286 ( .A(n206), .B(n660), .C(n810), .Q(n210) );
  NOR21 U1287 ( .A(n638), .B(n211), .Q(N1475) );
  AOI211 U1288 ( .A(n208), .B(n660), .C(n809), .Q(n211) );
  NOR21 U1289 ( .A(n638), .B(n212), .Q(N1473) );
  AOI211 U1290 ( .A(n599), .B(n658), .C(n810), .Q(n212) );
  NOR21 U1291 ( .A(n638), .B(n213), .Q(N1472) );
  AOI211 U1292 ( .A(n206), .B(n658), .C(n812), .Q(n213) );
  NOR21 U1293 ( .A(n638), .B(n214), .Q(N1471) );
  AOI211 U1294 ( .A(n208), .B(n658), .C(n811), .Q(n214) );
  NOR21 U1295 ( .A(n638), .B(n215), .Q(N1469) );
  AOI211 U1296 ( .A(n204), .B(n656), .C(n810), .Q(n215) );
  NOR21 U1297 ( .A(n638), .B(n216), .Q(N1468) );
  AOI211 U1298 ( .A(n206), .B(n656), .C(n807), .Q(n216) );
  NOR21 U1299 ( .A(n638), .B(n217), .Q(N1467) );
  AOI211 U1300 ( .A(n208), .B(n656), .C(n808), .Q(n217) );
  NOR21 U1301 ( .A(n638), .B(n218), .Q(N1465) );
  AOI211 U1302 ( .A(n599), .B(n654), .C(n812), .Q(n218) );
  NOR21 U1303 ( .A(n638), .B(n219), .Q(N1464) );
  AOI211 U1304 ( .A(n206), .B(n654), .C(n809), .Q(n219) );
  NOR21 U1305 ( .A(n637), .B(n220), .Q(N1463) );
  AOI211 U1306 ( .A(n208), .B(n654), .C(n810), .Q(n220) );
  NOR21 U1307 ( .A(n637), .B(n221), .Q(N1461) );
  AOI211 U1308 ( .A(n204), .B(n652), .C(n812), .Q(n221) );
  NOR21 U1309 ( .A(n637), .B(n222), .Q(N1460) );
  AOI211 U1310 ( .A(n206), .B(n652), .C(n811), .Q(n222) );
  NOR21 U1311 ( .A(n637), .B(n223), .Q(N1459) );
  AOI211 U1312 ( .A(n208), .B(n652), .C(n812), .Q(n223) );
  NOR21 U1313 ( .A(n637), .B(n224), .Q(N1457) );
  AOI211 U1314 ( .A(n599), .B(n650), .C(n807), .Q(n224) );
  NOR21 U1315 ( .A(n637), .B(n225), .Q(N1456) );
  AOI211 U1316 ( .A(n206), .B(n650), .C(n808), .Q(n225) );
  NOR21 U1317 ( .A(n637), .B(n226), .Q(N1455) );
  AOI211 U1318 ( .A(n208), .B(n650), .C(n809), .Q(n226) );
  NOR21 U1319 ( .A(n637), .B(n227), .Q(N1453) );
  AOI211 U1320 ( .A(n204), .B(n648), .C(n810), .Q(n227) );
  NOR21 U1321 ( .A(n637), .B(n228), .Q(N1452) );
  AOI211 U1322 ( .A(n206), .B(n648), .C(n812), .Q(n228) );
  NOR21 U1323 ( .A(n637), .B(n229), .Q(N1451) );
  AOI211 U1324 ( .A(n208), .B(n648), .C(n811), .Q(n229) );
  NOR21 U1325 ( .A(n637), .B(n230), .Q(N1449) );
  AOI211 U1326 ( .A(n599), .B(n646), .C(n811), .Q(n230) );
  NOR21 U1327 ( .A(n637), .B(n231), .Q(N1448) );
  AOI211 U1328 ( .A(n206), .B(n646), .C(n812), .Q(n231) );
  NOR21 U1329 ( .A(n637), .B(n232), .Q(N1447) );
  AOI211 U1330 ( .A(n208), .B(n646), .C(n807), .Q(n232) );
  NOR21 U1331 ( .A(n636), .B(n233), .Q(N1445) );
  AOI211 U1332 ( .A(n204), .B(n644), .C(n811), .Q(n233) );
  NOR21 U1333 ( .A(n636), .B(n234), .Q(N1444) );
  AOI211 U1334 ( .A(n206), .B(n644), .C(n809), .Q(n234) );
  NOR21 U1335 ( .A(n636), .B(n235), .Q(N1443) );
  AOI211 U1336 ( .A(n208), .B(n644), .C(n810), .Q(n235) );
  NOR21 U1337 ( .A(n636), .B(n236), .Q(N1441) );
  AOI211 U1338 ( .A(n599), .B(n642), .C(n812), .Q(n236) );
  NOR21 U1339 ( .A(n636), .B(n237), .Q(N1440) );
  AOI211 U1340 ( .A(n206), .B(n642), .C(n811), .Q(n237) );
  NOR21 U1341 ( .A(n636), .B(n238), .Q(N1439) );
  AOI211 U1342 ( .A(n208), .B(n642), .C(n809), .Q(n238) );
  NOR21 U1343 ( .A(n636), .B(n239), .Q(N1437) );
  AOI211 U1344 ( .A(n599), .B(n864), .C(n811), .Q(n239) );
  NOR21 U1345 ( .A(n636), .B(n240), .Q(N1436) );
  AOI211 U1346 ( .A(n206), .B(n864), .C(n807), .Q(n240) );
  NOR21 U1347 ( .A(n636), .B(n241), .Q(N1435) );
  AOI211 U1348 ( .A(n208), .B(n864), .C(n808), .Q(n241) );
  NOR21 U1349 ( .A(n636), .B(n242), .Q(N1433) );
  AOI211 U1350 ( .A(n599), .B(n866), .C(n807), .Q(n242) );
  NOR21 U1351 ( .A(n636), .B(n243), .Q(N1432) );
  AOI211 U1352 ( .A(n206), .B(n866), .C(n809), .Q(n243) );
  NOR21 U1353 ( .A(n636), .B(n244), .Q(N1431) );
  AOI211 U1354 ( .A(n208), .B(n866), .C(n810), .Q(n244) );
  NOR21 U1355 ( .A(n636), .B(n245), .Q(N1429) );
  AOI211 U1356 ( .A(n599), .B(n862), .C(n809), .Q(n245) );
  NOR21 U1357 ( .A(n635), .B(n246), .Q(N1428) );
  AOI211 U1358 ( .A(n206), .B(n862), .C(n809), .Q(n246) );
  NOR21 U1359 ( .A(n635), .B(n247), .Q(N1427) );
  AOI211 U1360 ( .A(n208), .B(n862), .C(n809), .Q(n247) );
  NOR21 U1361 ( .A(n635), .B(n248), .Q(N1425) );
  AOI211 U1362 ( .A(n599), .B(n865), .C(n809), .Q(n248) );
  NOR21 U1363 ( .A(n635), .B(n249), .Q(N1424) );
  AOI211 U1364 ( .A(n206), .B(n865), .C(n809), .Q(n249) );
  NOR21 U1365 ( .A(n635), .B(n250), .Q(N1423) );
  AOI211 U1366 ( .A(n208), .B(n865), .C(n809), .Q(n250) );
  NOR21 U1367 ( .A(n635), .B(n252), .Q(N1421) );
  AOI211 U1368 ( .A(n599), .B(n863), .C(n809), .Q(n252) );
  NOR21 U1369 ( .A(n635), .B(n253), .Q(N1420) );
  AOI211 U1370 ( .A(n206), .B(n863), .C(n809), .Q(n253) );
  NOR21 U1371 ( .A(n635), .B(n254), .Q(N1419) );
  AOI211 U1372 ( .A(n208), .B(n863), .C(n809), .Q(n254) );
  NOR21 U1373 ( .A(n635), .B(n256), .Q(N1417) );
  AOI211 U1374 ( .A(n257), .B(n662), .C(n809), .Q(n256) );
  NOR21 U1375 ( .A(n635), .B(n258), .Q(N1416) );
  AOI211 U1376 ( .A(n259), .B(n662), .C(n809), .Q(n258) );
  NOR21 U1377 ( .A(n635), .B(n260), .Q(N1415) );
  AOI211 U1378 ( .A(n261), .B(n662), .C(n809), .Q(n260) );
  NOR21 U1379 ( .A(n635), .B(n262), .Q(N1413) );
  AOI211 U1380 ( .A(n257), .B(n660), .C(n809), .Q(n262) );
  NOR21 U1381 ( .A(n635), .B(n263), .Q(N1412) );
  AOI211 U1382 ( .A(n259), .B(n660), .C(n809), .Q(n263) );
  NOR21 U1383 ( .A(n634), .B(n264), .Q(N1411) );
  AOI211 U1384 ( .A(n261), .B(n660), .C(n809), .Q(n264) );
  NOR21 U1385 ( .A(n634), .B(n265), .Q(N1409) );
  AOI211 U1386 ( .A(n257), .B(n658), .C(n809), .Q(n265) );
  NOR21 U1387 ( .A(n634), .B(n266), .Q(N1408) );
  AOI211 U1388 ( .A(n259), .B(n658), .C(n809), .Q(n266) );
  NOR21 U1389 ( .A(n634), .B(n267), .Q(N1407) );
  AOI211 U1390 ( .A(n261), .B(n658), .C(n809), .Q(n267) );
  NOR21 U1391 ( .A(n634), .B(n268), .Q(N1405) );
  AOI211 U1392 ( .A(n257), .B(n656), .C(n810), .Q(n268) );
  NOR21 U1393 ( .A(n634), .B(n269), .Q(N1404) );
  AOI211 U1394 ( .A(n259), .B(n656), .C(n810), .Q(n269) );
  NOR21 U1395 ( .A(n634), .B(n270), .Q(N1403) );
  AOI211 U1396 ( .A(n261), .B(n656), .C(n810), .Q(n270) );
  NOR21 U1397 ( .A(n634), .B(n271), .Q(N1401) );
  AOI211 U1398 ( .A(n257), .B(n654), .C(n810), .Q(n271) );
  NOR21 U1399 ( .A(n634), .B(n272), .Q(N1400) );
  AOI211 U1400 ( .A(n259), .B(n654), .C(n810), .Q(n272) );
  NOR21 U1401 ( .A(n634), .B(n273), .Q(N1399) );
  AOI211 U1402 ( .A(n261), .B(n654), .C(n810), .Q(n273) );
  NOR21 U1403 ( .A(n634), .B(n274), .Q(N1397) );
  AOI211 U1404 ( .A(n257), .B(n652), .C(n810), .Q(n274) );
  NOR21 U1405 ( .A(n634), .B(n275), .Q(N1396) );
  AOI211 U1406 ( .A(n259), .B(n652), .C(n810), .Q(n275) );
  NOR21 U1407 ( .A(n634), .B(n276), .Q(N1395) );
  AOI211 U1408 ( .A(n261), .B(n652), .C(n810), .Q(n276) );
  NOR21 U1409 ( .A(n633), .B(n277), .Q(N1393) );
  AOI211 U1410 ( .A(n257), .B(n650), .C(n810), .Q(n277) );
  NOR21 U1411 ( .A(n633), .B(n278), .Q(N1392) );
  AOI211 U1412 ( .A(n259), .B(n650), .C(n810), .Q(n278) );
  NOR21 U1413 ( .A(n633), .B(n279), .Q(N1391) );
  AOI211 U1414 ( .A(n261), .B(n650), .C(n810), .Q(n279) );
  NOR21 U1415 ( .A(n633), .B(n280), .Q(N1389) );
  AOI211 U1416 ( .A(n257), .B(n648), .C(n810), .Q(n280) );
  NOR21 U1417 ( .A(n633), .B(n281), .Q(N1388) );
  AOI211 U1418 ( .A(n259), .B(n648), .C(n810), .Q(n281) );
  NOR21 U1419 ( .A(n633), .B(n282), .Q(N1387) );
  AOI211 U1420 ( .A(n261), .B(n648), .C(n810), .Q(n282) );
  NOR21 U1421 ( .A(n633), .B(n283), .Q(N1385) );
  AOI211 U1422 ( .A(n257), .B(n646), .C(n810), .Q(n283) );
  NOR21 U1423 ( .A(n633), .B(n284), .Q(N1384) );
  AOI211 U1424 ( .A(n259), .B(n646), .C(n810), .Q(n284) );
  NOR21 U1425 ( .A(n633), .B(n285), .Q(N1383) );
  AOI211 U1426 ( .A(n261), .B(n646), .C(n810), .Q(n285) );
  NOR21 U1427 ( .A(n633), .B(n286), .Q(N1381) );
  AOI211 U1428 ( .A(n257), .B(n644), .C(n810), .Q(n286) );
  NOR21 U1429 ( .A(n633), .B(n287), .Q(N1380) );
  AOI211 U1430 ( .A(n259), .B(n644), .C(n811), .Q(n287) );
  NOR21 U1431 ( .A(n633), .B(n288), .Q(N1379) );
  AOI211 U1432 ( .A(n261), .B(n644), .C(n811), .Q(n288) );
  NOR21 U1433 ( .A(n633), .B(n289), .Q(N1377) );
  AOI211 U1434 ( .A(n257), .B(n642), .C(n811), .Q(n289) );
  NOR21 U1435 ( .A(n633), .B(n290), .Q(N1376) );
  AOI211 U1436 ( .A(n259), .B(n642), .C(n811), .Q(n290) );
  NOR21 U1437 ( .A(n637), .B(n291), .Q(N1375) );
  AOI211 U1438 ( .A(n261), .B(n642), .C(n811), .Q(n291) );
  NOR21 U1439 ( .A(n636), .B(n292), .Q(N1373) );
  AOI211 U1440 ( .A(n257), .B(n864), .C(n811), .Q(n292) );
  NOR21 U1441 ( .A(n635), .B(n293), .Q(N1372) );
  AOI211 U1442 ( .A(n259), .B(n864), .C(n811), .Q(n293) );
  NOR21 U1443 ( .A(n634), .B(n294), .Q(N1371) );
  AOI211 U1444 ( .A(n261), .B(n864), .C(n811), .Q(n294) );
  NOR21 U1445 ( .A(n633), .B(n295), .Q(N1369) );
  AOI211 U1446 ( .A(n257), .B(n866), .C(n811), .Q(n295) );
  NOR21 U1447 ( .A(n639), .B(n296), .Q(N1368) );
  AOI211 U1448 ( .A(n259), .B(n866), .C(n811), .Q(n296) );
  NOR21 U1449 ( .A(n638), .B(n297), .Q(N1367) );
  AOI211 U1450 ( .A(n261), .B(n866), .C(n811), .Q(n297) );
  NOR21 U1451 ( .A(n639), .B(n298), .Q(N1365) );
  AOI211 U1452 ( .A(n257), .B(n862), .C(n811), .Q(n298) );
  NOR21 U1453 ( .A(n637), .B(n299), .Q(N1364) );
  AOI211 U1454 ( .A(n259), .B(n862), .C(n811), .Q(n299) );
  NOR21 U1455 ( .A(n636), .B(n300), .Q(N1363) );
  AOI211 U1456 ( .A(n261), .B(n862), .C(n811), .Q(n300) );
  NOR21 U1457 ( .A(n635), .B(n301), .Q(N1361) );
  AOI211 U1458 ( .A(n257), .B(n865), .C(n811), .Q(n301) );
  NOR21 U1459 ( .A(n634), .B(n302), .Q(N1360) );
  AOI211 U1460 ( .A(n259), .B(n865), .C(n811), .Q(n302) );
  NOR21 U1461 ( .A(n637), .B(n303), .Q(N1359) );
  AOI211 U1462 ( .A(n261), .B(n865), .C(n811), .Q(n303) );
  NOR21 U1463 ( .A(n636), .B(n305), .Q(N1357) );
  AOI211 U1464 ( .A(n257), .B(n863), .C(n811), .Q(n305) );
  NOR21 U1465 ( .A(n635), .B(n306), .Q(N1356) );
  AOI211 U1466 ( .A(n259), .B(n863), .C(n811), .Q(n306) );
  NOR21 U1467 ( .A(n634), .B(n307), .Q(N1355) );
  AOI211 U1468 ( .A(n261), .B(n863), .C(n812), .Q(n307) );
  NOR21 U1469 ( .A(n639), .B(n309), .Q(N1353) );
  AOI211 U1470 ( .A(n588), .B(n662), .C(n812), .Q(n309) );
  NOR21 U1471 ( .A(n638), .B(n311), .Q(N1352) );
  AOI211 U1472 ( .A(n312), .B(n662), .C(n812), .Q(n311) );
  NOR21 U1473 ( .A(n633), .B(n313), .Q(N1351) );
  AOI211 U1474 ( .A(n314), .B(n662), .C(n812), .Q(n313) );
  NOR21 U1475 ( .A(n637), .B(n317), .Q(N1349) );
  AOI211 U1476 ( .A(n588), .B(n660), .C(n812), .Q(n317) );
  NOR21 U1477 ( .A(n636), .B(n318), .Q(N1348) );
  AOI211 U1478 ( .A(n312), .B(n660), .C(n812), .Q(n318) );
  NOR21 U1479 ( .A(n635), .B(n319), .Q(N1347) );
  AOI211 U1480 ( .A(n314), .B(n660), .C(n812), .Q(n319) );
  NOR21 U1481 ( .A(n634), .B(n321), .Q(N1345) );
  AOI211 U1482 ( .A(n588), .B(n658), .C(n812), .Q(n321) );
  NOR21 U1483 ( .A(n639), .B(n322), .Q(N1344) );
  AOI211 U1484 ( .A(n312), .B(n658), .C(n812), .Q(n322) );
  NOR21 U1485 ( .A(n638), .B(n323), .Q(N1343) );
  AOI211 U1486 ( .A(n314), .B(n658), .C(n812), .Q(n323) );
  NOR21 U1487 ( .A(n638), .B(n325), .Q(N1341) );
  AOI211 U1488 ( .A(n310), .B(n656), .C(n812), .Q(n325) );
  NOR21 U1489 ( .A(n639), .B(n326), .Q(N1340) );
  AOI211 U1490 ( .A(n312), .B(n656), .C(n812), .Q(n326) );
  NOR21 U1491 ( .A(n638), .B(n327), .Q(N1339) );
  AOI211 U1492 ( .A(n314), .B(n656), .C(n812), .Q(n327) );
  NOR21 U1493 ( .A(n633), .B(n329), .Q(N1337) );
  AOI211 U1494 ( .A(n588), .B(n654), .C(n812), .Q(n329) );
  NOR21 U1495 ( .A(n637), .B(n330), .Q(N1336) );
  AOI211 U1496 ( .A(n312), .B(n654), .C(n812), .Q(n330) );
  NOR21 U1497 ( .A(n636), .B(n331), .Q(N1335) );
  AOI211 U1498 ( .A(n314), .B(n654), .C(n812), .Q(n331) );
  NOR21 U1499 ( .A(n635), .B(n333), .Q(N1333) );
  AOI211 U1500 ( .A(n310), .B(n652), .C(n812), .Q(n333) );
  NOR21 U1501 ( .A(n634), .B(n334), .Q(N1332) );
  AOI211 U1502 ( .A(n312), .B(n652), .C(n812), .Q(n334) );
  NOR21 U1503 ( .A(n633), .B(n335), .Q(N1331) );
  AOI211 U1504 ( .A(n314), .B(n652), .C(n812), .Q(n335) );
  NOR21 U1505 ( .A(n637), .B(n336), .Q(N1329) );
  AOI211 U1506 ( .A(n588), .B(n650), .C(n807), .Q(n336) );
  NOR21 U1507 ( .A(n639), .B(n337), .Q(N1328) );
  AOI211 U1508 ( .A(n312), .B(n650), .C(n808), .Q(n337) );
  NOR21 U1509 ( .A(n638), .B(n338), .Q(N1327) );
  AOI211 U1510 ( .A(n314), .B(n650), .C(n810), .Q(n338) );
  NOR21 U1511 ( .A(n639), .B(n339), .Q(N1325) );
  AOI211 U1512 ( .A(n310), .B(n648), .C(n812), .Q(n339) );
  NOR21 U1513 ( .A(n636), .B(n340), .Q(N1324) );
  AOI211 U1514 ( .A(n312), .B(n648), .C(n811), .Q(n340) );
  NOR21 U1515 ( .A(n635), .B(n341), .Q(N1323) );
  AOI211 U1516 ( .A(n314), .B(n648), .C(n809), .Q(n341) );
  NOR21 U1517 ( .A(n634), .B(n342), .Q(N1321) );
  AOI211 U1518 ( .A(n588), .B(n646), .C(n807), .Q(n342) );
  NOR21 U1519 ( .A(n633), .B(n343), .Q(N1320) );
  AOI211 U1520 ( .A(n312), .B(n646), .C(n808), .Q(n343) );
  NOR21 U1521 ( .A(n636), .B(n344), .Q(N1319) );
  AOI211 U1522 ( .A(n314), .B(n646), .C(n810), .Q(n344) );
  NOR21 U1523 ( .A(n638), .B(n346), .Q(N1317) );
  AOI211 U1524 ( .A(n310), .B(n644), .C(n812), .Q(n346) );
  NOR21 U1525 ( .A(n639), .B(n347), .Q(N1316) );
  AOI211 U1526 ( .A(n312), .B(n644), .C(n811), .Q(n347) );
  NOR21 U1527 ( .A(n637), .B(n348), .Q(N1315) );
  AOI211 U1528 ( .A(n314), .B(n644), .C(n809), .Q(n348) );
  NOR21 U1529 ( .A(n636), .B(n349), .Q(N1313) );
  AOI211 U1530 ( .A(n588), .B(n642), .C(n807), .Q(n349) );
  NOR21 U1531 ( .A(n635), .B(n350), .Q(N1312) );
  AOI211 U1532 ( .A(n312), .B(n642), .C(n808), .Q(n350) );
  NOR21 U1533 ( .A(n634), .B(n351), .Q(N1311) );
  AOI211 U1534 ( .A(n314), .B(n642), .C(n810), .Q(n351) );
  NOR21 U1535 ( .A(n633), .B(n352), .Q(N1309) );
  AOI211 U1536 ( .A(n310), .B(n864), .C(n812), .Q(n352) );
  NOR21 U1537 ( .A(n635), .B(n353), .Q(N1308) );
  AOI211 U1538 ( .A(n312), .B(n864), .C(n811), .Q(n353) );
  NOR21 U1539 ( .A(n639), .B(n354), .Q(N1307) );
  AOI211 U1540 ( .A(n314), .B(n864), .C(n809), .Q(n354) );
  NOR21 U1541 ( .A(n638), .B(n355), .Q(N1305) );
  AOI211 U1542 ( .A(n588), .B(n866), .C(n807), .Q(n355) );
  NOR21 U1543 ( .A(n637), .B(n356), .Q(N1304) );
  AOI211 U1544 ( .A(n312), .B(n866), .C(n807), .Q(n356) );
  NOR21 U1545 ( .A(n636), .B(n357), .Q(N1303) );
  AOI211 U1546 ( .A(n314), .B(n866), .C(n809), .Q(n357) );
  NOR21 U1547 ( .A(n635), .B(n359), .Q(N1301) );
  AOI211 U1548 ( .A(n588), .B(n862), .C(n807), .Q(n359) );
  NOR21 U1549 ( .A(n634), .B(n360), .Q(N1300) );
  AOI211 U1550 ( .A(n312), .B(n862), .C(n807), .Q(n360) );
  NOR21 U1551 ( .A(n633), .B(n361), .Q(N1299) );
  AOI211 U1552 ( .A(n314), .B(n862), .C(n807), .Q(n361) );
  NOR21 U1553 ( .A(n634), .B(n362), .Q(N1297) );
  AOI211 U1554 ( .A(n588), .B(n865), .C(n808), .Q(n362) );
  NOR21 U1555 ( .A(n633), .B(n363), .Q(N1296) );
  AOI211 U1556 ( .A(n312), .B(n865), .C(n807), .Q(n363) );
  NOR21 U1557 ( .A(n638), .B(n364), .Q(N1295) );
  AOI211 U1558 ( .A(n314), .B(n865), .C(n810), .Q(n364) );
  NOR21 U1559 ( .A(n637), .B(n367), .Q(N1293) );
  AOI211 U1560 ( .A(n588), .B(n863), .C(n807), .Q(n367) );
  NOR21 U1561 ( .A(n639), .B(n368), .Q(N1292) );
  AOI211 U1562 ( .A(n312), .B(n863), .C(n812), .Q(n368) );
  NOR21 U1563 ( .A(n638), .B(n369), .Q(N1291) );
  AOI211 U1564 ( .A(n314), .B(n863), .C(n808), .Q(n369) );
  NOR21 U1565 ( .A(n640), .B(n185), .Q(N1499) );
  AOI211 U1566 ( .A(n186), .B(n864), .C(n808), .Q(n185) );
  INV3 U1567 ( .A(n107), .Q(n877) );
  BUF2 U1568 ( .A(n663), .Q(n738) );
  BUF2 U1569 ( .A(n663), .Q(n739) );
  BUF2 U1570 ( .A(n663), .Q(n740) );
  BUF2 U1571 ( .A(n664), .Q(n741) );
  BUF2 U1572 ( .A(n664), .Q(n742) );
  BUF2 U1573 ( .A(n664), .Q(n743) );
  BUF2 U1574 ( .A(n665), .Q(n744) );
  BUF2 U1575 ( .A(n665), .Q(n745) );
  BUF2 U1576 ( .A(n665), .Q(n746) );
  BUF2 U1577 ( .A(n666), .Q(n747) );
  BUF2 U1578 ( .A(n666), .Q(n748) );
  BUF2 U1579 ( .A(n666), .Q(n749) );
  BUF2 U1580 ( .A(n667), .Q(n750) );
  BUF2 U1581 ( .A(n667), .Q(n751) );
  BUF2 U1582 ( .A(n667), .Q(n752) );
  BUF2 U1583 ( .A(n668), .Q(n753) );
  BUF2 U1584 ( .A(n668), .Q(n754) );
  BUF2 U1585 ( .A(n668), .Q(n755) );
  BUF2 U1586 ( .A(n669), .Q(n756) );
  BUF2 U1587 ( .A(n669), .Q(n757) );
  BUF2 U1588 ( .A(n669), .Q(n758) );
  BUF2 U1589 ( .A(n670), .Q(n759) );
  BUF2 U1590 ( .A(n670), .Q(n760) );
  BUF2 U1591 ( .A(n670), .Q(n761) );
  BUF2 U1592 ( .A(n671), .Q(n762) );
  BUF2 U1593 ( .A(n671), .Q(n763) );
  BUF2 U1594 ( .A(n671), .Q(n764) );
  BUF2 U1595 ( .A(n672), .Q(n765) );
  BUF2 U1596 ( .A(n672), .Q(n766) );
  BUF2 U1597 ( .A(n672), .Q(n767) );
  BUF2 U1598 ( .A(n673), .Q(n768) );
  BUF2 U1599 ( .A(n673), .Q(n769) );
  NOR40 U1600 ( .A(n872), .B(n905), .C(N145), .D(N144), .Q(N1269) );
  NAND22 U1601 ( .A(N150), .B(n873), .Q(n905) );
  INV3 U1602 ( .A(n904), .Q(n872) );
  INV3 U1603 ( .A(N143), .Q(n873) );
  NOR40 U1604 ( .A(N149), .B(N148), .C(N147), .D(N146), .Q(n904) );
  AOI211 U1605 ( .A(n103), .B(n867), .C(n106), .Q(n104) );
  INV3 U1606 ( .A(N1270), .Q(n867) );
  INV3 U1607 ( .A(n155), .Q(n838) );
  AOI221 U1608 ( .A(N125), .B(n148), .C(N149), .D(n149), .Q(n155) );
  NOR21 U1609 ( .A(n119), .B(n640), .Q(n146) );
  NOR21 U1610 ( .A(n120), .B(n640), .Q(n145) );
  NAND22 U1611 ( .A(n774), .B(n365), .Q(N183) );
  INV3 U1612 ( .A(n545), .Q(n581) );
  NAND22 U1613 ( .A(n167), .B(n145), .Q(n163) );
  NAND22 U1614 ( .A(n161), .B(n145), .Q(n152) );
  NAND22 U1615 ( .A(n161), .B(n146), .Q(n153) );
  NAND22 U1616 ( .A(n167), .B(n146), .Q(n164) );
  NAND22 U1617 ( .A(n161), .B(n150), .Q(n154) );
  NAND22 U1618 ( .A(n167), .B(n150), .Q(n165) );
  NAND22 U1619 ( .A(n146), .B(n144), .Q(n127) );
  NAND22 U1620 ( .A(n145), .B(n144), .Q(n126) );
  NAND22 U1621 ( .A(n150), .B(n144), .Q(n128) );
  INV3 U1622 ( .A(n903), .Q(n868) );
  XNR21 U1623 ( .A(\add_256/carry [6]), .B(n583), .Q(n576) );
  NOR21 U1624 ( .A(n857), .B(n810), .Q(N164) );
  INV3 U1625 ( .A(N132), .Q(n857) );
  INV3 U1626 ( .A(n157), .Q(n836) );
  AOI221 U1627 ( .A(N123), .B(n148), .C(N147), .D(n149), .Q(n157) );
  INV3 U1628 ( .A(n156), .Q(n837) );
  AOI221 U1629 ( .A(N124), .B(n148), .C(N148), .D(n149), .Q(n156) );
  NOR21 U1630 ( .A(n557), .B(n543), .Q(n358) );
  NOR21 U1631 ( .A(n556), .B(n542), .Q(n328) );
  AOI211 U1632 ( .A(n116), .B(n572), .C(n370), .Q(N1286) );
  NAND31 U1633 ( .A(n544), .B(n563), .C(n583), .Q(n198) );
  NOR31 U1634 ( .A(n544), .B(n583), .C(n563), .Q(n175) );
  NAND22 U1635 ( .A(n569), .B(n547), .Q(n184) );
  NAND22 U1636 ( .A(n345), .B(n328), .Q(n139) );
  NAND22 U1637 ( .A(n358), .B(n324), .Q(n142) );
  NAND22 U1638 ( .A(n345), .B(n328), .Q(n595) );
  AOI211 U1639 ( .A(n546), .B(n102), .C(n875), .Q(n122) );
  NAND22 U1640 ( .A(n358), .B(n315), .Q(n140) );
  NAND22 U1641 ( .A(n358), .B(n320), .Q(n141) );
  NAND22 U1642 ( .A(n332), .B(n328), .Q(n135) );
  NAND22 U1643 ( .A(n332), .B(n324), .Q(n134) );
  NAND22 U1644 ( .A(n345), .B(n324), .Q(n138) );
  NAND22 U1645 ( .A(n332), .B(n315), .Q(n132) );
  NAND22 U1646 ( .A(n345), .B(n315), .Q(n136) );
  NAND22 U1647 ( .A(n332), .B(n320), .Q(n133) );
  NAND22 U1648 ( .A(n345), .B(n320), .Q(n137) );
  NAND22 U1649 ( .A(n358), .B(n315), .Q(n594) );
  NAND22 U1650 ( .A(n315), .B(n316), .Q(n124) );
  NAND22 U1651 ( .A(n320), .B(n316), .Q(n129) );
  NAND22 U1652 ( .A(n324), .B(n316), .Q(n130) );
  NAND22 U1653 ( .A(n328), .B(n316), .Q(n131) );
  NAND22 U1654 ( .A(n358), .B(n320), .Q(n593) );
  NAND22 U1655 ( .A(n102), .B(n548), .Q(n118) );
  NAND22 U1656 ( .A(n358), .B(n324), .Q(n592) );
  NAND22 U1657 ( .A(n358), .B(n324), .Q(n591) );
  BUF2 U1658 ( .A(n823), .Q(n830) );
  BUF2 U1659 ( .A(n823), .Q(n829) );
  BUF2 U1660 ( .A(n821), .Q(n827) );
  BUF2 U1661 ( .A(n822), .Q(n828) );
  BUF2 U1662 ( .A(n820), .Q(n826) );
  BUF2 U1663 ( .A(n820), .Q(n825) );
  NOR21 U1664 ( .A(n148), .B(n370), .Q(N1287) );
  AOI211 U1665 ( .A(n546), .B(n116), .C(n117), .Q(n105) );
  NOR21 U1666 ( .A(n198), .B(n119), .Q(n190) );
  NOR21 U1667 ( .A(n198), .B(n120), .Q(n188) );
  NAND31 U1668 ( .A(n771), .B(n121), .C(n122), .Q(N1806) );
  NAND31 U1669 ( .A(n770), .B(n123), .C(n122), .Q(N1804) );
  AOI211 U1670 ( .A(n112), .B(sig_fsm_start_R), .C(n877), .Q(n115) );
  BUF2 U1671 ( .A(n582), .Q(n815) );
  BUF2 U1672 ( .A(n582), .Q(n816) );
  BUF2 U1673 ( .A(n582), .Q(n817) );
  BUF2 U1674 ( .A(n582), .Q(n818) );
  NOR21 U1675 ( .A(n365), .B(n807), .Q(n117) );
  NAND22 U1676 ( .A(N198), .B(n144), .Q(n125) );
  NAND22 U1677 ( .A(n161), .B(N198), .Q(n151) );
  NAND22 U1678 ( .A(n167), .B(N198), .Q(n162) );
  NOR31 U1679 ( .A(n547), .B(n831), .C(n569), .Q(N198) );
  INV3 U1680 ( .A(n204), .Q(n598) );
  NOR21 U1681 ( .A(n251), .B(n120), .Q(n204) );
  NOR21 U1682 ( .A(n251), .B(n119), .Q(n206) );
  NOR21 U1683 ( .A(n251), .B(n184), .Q(n208) );
  NOR21 U1684 ( .A(n304), .B(n120), .Q(n257) );
  NOR21 U1685 ( .A(n304), .B(n119), .Q(n259) );
  NOR21 U1686 ( .A(n304), .B(n184), .Q(n261) );
  INV3 U1687 ( .A(n310), .Q(n587) );
  NOR21 U1688 ( .A(n366), .B(n120), .Q(n310) );
  NOR21 U1689 ( .A(n366), .B(n119), .Q(n312) );
  NOR21 U1690 ( .A(n366), .B(n184), .Q(n314) );
  NAND22 U1691 ( .A(n855), .B(N198), .Q(n202) );
  INV3 U1692 ( .A(n251), .Q(n855) );
  NAND22 U1693 ( .A(n854), .B(N198), .Q(n255) );
  INV3 U1694 ( .A(n304), .Q(n854) );
  NAND22 U1695 ( .A(n853), .B(N198), .Q(n308) );
  INV3 U1696 ( .A(n366), .Q(n853) );
  NOR21 U1697 ( .A(n858), .B(n812), .Q(N163) );
  INV3 U1698 ( .A(N131), .Q(n858) );
  NOR21 U1699 ( .A(n859), .B(n811), .Q(N162) );
  INV3 U1700 ( .A(N130), .Q(n859) );
  NOR21 U1701 ( .A(n860), .B(n811), .Q(N161) );
  INV3 U1702 ( .A(N129), .Q(n860) );
  BUF2 U1703 ( .A(n582), .Q(n819) );
  INV3 U1704 ( .A(n160), .Q(n833) );
  AOI221 U1705 ( .A(N120), .B(n148), .C(N144), .D(n149), .Q(n160) );
  INV3 U1706 ( .A(n158), .Q(n835) );
  AOI221 U1707 ( .A(N122), .B(n148), .C(N146), .D(n149), .Q(n158) );
  INV3 U1708 ( .A(n159), .Q(n834) );
  AOI221 U1709 ( .A(N121), .B(n148), .C(N145), .D(n149), .Q(n159) );
  INV3 U1710 ( .A(n899), .Q(n870) );
  NAND22 U1711 ( .A(n549), .B(n900), .Q(n899) );
  INV3 U1712 ( .A(n173), .Q(n845) );
  NAND22 U1713 ( .A(n116), .B(N140), .Q(n173) );
  INV3 U1714 ( .A(n174), .Q(n844) );
  NAND22 U1715 ( .A(n116), .B(N139), .Q(n174) );
  INV3 U1716 ( .A(n176), .Q(n843) );
  NAND22 U1717 ( .A(n116), .B(N138), .Q(n176) );
  INV3 U1718 ( .A(n181), .Q(n842) );
  NAND22 U1719 ( .A(n116), .B(N137), .Q(n181) );
  INV3 U1720 ( .A(n182), .Q(n841) );
  NAND22 U1721 ( .A(n116), .B(N136), .Q(n182) );
  INV3 U1722 ( .A(n183), .Q(n840) );
  NAND22 U1723 ( .A(n116), .B(n550), .Q(n183) );
  NAND31 U1724 ( .A(n548), .B(n575), .C(n113), .Q(n107) );
  NAND22 U1725 ( .A(n773), .B(n118), .Q(N213) );
  AOI211 U1726 ( .A(n119), .B(n120), .C(n808), .Q(N192) );
  NOR21 U1727 ( .A(n572), .B(n807), .Q(n148) );
  INV3 U1728 ( .A(n108), .Q(n878) );
  NOR21 U1729 ( .A(n807), .B(n121), .Q(N1276) );
  NOR21 U1730 ( .A(n807), .B(n123), .Q(N1277) );
  NOR21 U1731 ( .A(n824), .B(n807), .Q(N222) );
  NOR21 U1732 ( .A(n861), .B(n808), .Q(N160) );
  INV3 U1733 ( .A(N128), .Q(n861) );
  INV3 U1734 ( .A(n112), .Q(n879) );
  INV3 U1735 ( .A(n166), .Q(n832) );
  AOI221 U1736 ( .A(n552), .B(n148), .C(N143), .D(n149), .Q(n166) );
  INV3 U1737 ( .A(n773), .Q(n808) );
  INV3 U1738 ( .A(n773), .Q(n807) );
  INV3 U1739 ( .A(n771), .Q(n809) );
  INV3 U1740 ( .A(n771), .Q(n810) );
  INV3 U1741 ( .A(n770), .Q(n811) );
  INV3 U1742 ( .A(n771), .Q(n812) );
  AOI2111 U1743 ( .A(N148), .B(n909), .C(N150), .D(N149), .Q(N1285) );
  NAND22 U1744 ( .A(n908), .B(n907), .Q(n909) );
  NOR21 U1745 ( .A(N144), .B(N143), .Q(n908) );
  NOR31 U1746 ( .A(N145), .B(N147), .C(N146), .Q(n907) );
  BUF2 U1747 ( .A(N918), .Q(n663) );
  BUF2 U1748 ( .A(N918), .Q(n664) );
  BUF2 U1749 ( .A(N918), .Q(n665) );
  BUF2 U1750 ( .A(N918), .Q(n666) );
  BUF2 U1751 ( .A(N918), .Q(n667) );
  BUF2 U1752 ( .A(N918), .Q(n668) );
  BUF2 U1753 ( .A(N918), .Q(n669) );
  BUF2 U1754 ( .A(N918), .Q(n670) );
  BUF2 U1755 ( .A(N918), .Q(n671) );
  BUF2 U1756 ( .A(N918), .Q(n672) );
  BUF2 U1757 ( .A(N918), .Q(n673) );
  INV3 U1758 ( .A(n906), .Q(outAlmostFull) );
  AOI211 U1759 ( .A(N149), .B(N148), .C(N150), .Q(n906) );
  INV3 U1760 ( .A(n578), .Q(\r98/carry [1]) );
  NOR21 U1761 ( .A(n550), .B(outWriteCount[0]), .Q(n578) );
  XNR21 U1762 ( .A(\r98/carry [7]), .B(outWriteCount[7]), .Q(N150) );
  AOI211 U1763 ( .A(n100), .B(n101), .C(n809), .Q(N50) );
  AOI221 U1764 ( .A(currentState[1]), .B(n102), .C(n868), .D(n878), .Q(n101)
         );
  AOI221 U1765 ( .A(N1269), .B(n877), .C(N1270), .D(n103), .Q(n100) );
  INV3 U1766 ( .A(n147), .Q(n839) );
  AOI221 U1767 ( .A(N126), .B(n148), .C(N150), .D(n149), .Q(n147) );
  XOR21 U1768 ( .A(\add_255/carry [7]), .B(outWriteCount[7]), .Q(N126) );
  NOR40 U1769 ( .A(n902), .B(n903), .C(n874), .D(n901), .Q(N1270) );
  INV3 U1770 ( .A(n898), .Q(n874) );
  NAND41 U1771 ( .A(n896), .B(n890), .C(n889), .D(n886), .Q(n902) );
  AOI211 U1772 ( .A(outWriteCount[1]), .B(n900), .C(n870), .Q(n901) );
  NAND31 U1773 ( .A(n102), .B(n546), .C(currentState[0]), .Q(n365) );
  OAI2111 U1774 ( .A(n892), .B(n891), .C(n890), .D(n889), .Q(n894) );
  NOR21 U1775 ( .A(outReadCount[3]), .B(n565), .Q(n892) );
  OAI2111 U1776 ( .A(n887), .B(n549), .C(n869), .D(n886), .Q(n888) );
  NOR21 U1777 ( .A(n558), .B(currentState[3]), .Q(n102) );
  AOI2111 U1778 ( .A(N1270), .B(n103), .C(n878), .D(n110), .Q(n109) );
  NOR31 U1779 ( .A(n879), .B(currentState[2]), .C(n111), .Q(n110) );
  XNR21 U1780 ( .A(sig_fsm_start_W), .B(sig_fsm_start_R), .Q(n111) );
  AOI311 U1781 ( .A(n898), .B(n896), .C(n895), .D(outWriteCount[7]), .Q(n897)
         );
  OAI2111 U1782 ( .A(outReadCount[5]), .B(n566), .C(n894), .D(n893), .Q(n895)
         );
  NAND22 U1783 ( .A(outWriteCount[4]), .B(n554), .Q(n893) );
  NOR21 U1784 ( .A(n552), .B(outReadCount[0]), .Q(n887) );
  BUF2 U1785 ( .A(N40), .Q(n582) );
  XNR21 U1786 ( .A(\add_360/carry [6]), .B(N45), .Q(n577) );
  INV3 U1787 ( .A(n885), .Q(n869) );
  AOI211 U1788 ( .A(n549), .B(n887), .C(outWriteCount[1]), .Q(n885) );
  INV3 U1789 ( .A(n172), .Q(n846) );
  NAND22 U1790 ( .A(n116), .B(N141), .Q(n172) );
  XOR21 U1791 ( .A(\add_260/carry [6]), .B(outReadCount[6]), .Q(N141) );
  NOR31 U1792 ( .A(i_FIFO[5]), .B(n583), .C(n544), .Q(n161) );
  NOR31 U1793 ( .A(i_FIFO[4]), .B(n583), .C(n563), .Q(n167) );
  NAND31 U1794 ( .A(i_FIFO[4]), .B(n563), .C(n583), .Q(n251) );
  NAND31 U1795 ( .A(i_FIFO[5]), .B(n544), .C(n583), .Q(n304) );
  NAND31 U1796 ( .A(i_FIFO[5]), .B(i_FIFO[4]), .C(n583), .Q(n366) );
  NOR31 U1797 ( .A(i_FIFO[5]), .B(n583), .C(i_FIFO[4]), .Q(n144) );
  NOR21 U1798 ( .A(n556), .B(i_FIFO[0]), .Q(n324) );
  NOR21 U1799 ( .A(i_FIFO[1]), .B(i_FIFO[0]), .Q(n315) );
  NOR21 U1800 ( .A(n542), .B(i_FIFO[1]), .Q(n320) );
  NAND22 U1801 ( .A(k_FIFO[1]), .B(n547), .Q(n120) );
  NAND22 U1802 ( .A(k_FIFO[0]), .B(n569), .Q(n119) );
  XNR21 U1803 ( .A(outWriteCount[0]), .B(n550), .Q(N143) );
  NOR21 U1804 ( .A(n557), .B(i_FIFO[2]), .Q(n345) );
  AOI2111 U1805 ( .A(n371), .B(n372), .C(n584), .D(n875), .Q(n370) );
  NOR40 U1806 ( .A(outWriteCount[2]), .B(outWriteCount[1]), .C(
        outWriteCount[0]), .D(n571), .Q(n371) );
  NOR40 U1807 ( .A(outWriteCount[6]), .B(outWriteCount[5]), .C(
        outWriteCount[4]), .D(outWriteCount[3]), .Q(n372) );
  NOR21 U1808 ( .A(i_FIFO[3]), .B(i_FIFO[2]), .Q(n316) );
  BUF2 U1809 ( .A(N42), .Q(n813) );
  NOR21 U1810 ( .A(n543), .B(i_FIFO[3]), .Q(n332) );
  BUF2 U1811 ( .A(N42), .Q(n814) );
  BUF2 U1812 ( .A(i_FIFO[6]), .Q(n583) );
  NAND22 U1813 ( .A(outReadCount[0]), .B(n552), .Q(n900) );
  NAND22 U1814 ( .A(outReadCount[6]), .B(n564), .Q(n898) );
  NAND22 U1815 ( .A(outReadCount[5]), .B(n566), .Q(n896) );
  NOR21 U1816 ( .A(n559), .B(n810), .Q(N206) );
  NOR21 U1817 ( .A(n560), .B(n812), .Q(N207) );
  NOR21 U1818 ( .A(n561), .B(n811), .Q(N208) );
  NOR21 U1819 ( .A(n562), .B(n809), .Q(N209) );
  NAND22 U1820 ( .A(outReadCount[3]), .B(n565), .Q(n889) );
  NAND22 U1821 ( .A(outReadCount[2]), .B(n553), .Q(n886) );
  NAND22 U1822 ( .A(outReadCount[4]), .B(n568), .Q(n890) );
  BUF2 U1823 ( .A(N43), .Q(n580) );
  INV3 U1824 ( .A(n149), .Q(n584) );
  NOR21 U1825 ( .A(n807), .B(sigEnableCounter), .Q(n149) );
  BUF2 U1826 ( .A(N39), .Q(n824) );
  BUF2 U1827 ( .A(N39), .Q(n823) );
  BUF2 U1828 ( .A(N39), .Q(n821) );
  BUF2 U1829 ( .A(N39), .Q(n822) );
  BUF2 U1830 ( .A(N39), .Q(n820) );
  NAND31 U1831 ( .A(n546), .B(n558), .C(currentState[0]), .Q(n114) );
  NAND31 U1832 ( .A(n113), .B(n575), .C(currentState[0]), .Q(n108) );
  NAND31 U1833 ( .A(currentState[3]), .B(n548), .C(n113), .Q(n121) );
  NOR21 U1834 ( .A(n546), .B(currentState[2]), .Q(n113) );
  NOR31 U1835 ( .A(currentState[1]), .B(currentState[3]), .C(currentState[0]), 
        .Q(n112) );
  NOR21 U1836 ( .A(n114), .B(currentState[3]), .Q(n103) );
  BUF2 U1837 ( .A(N44), .Q(n579) );
  NOR21 U1838 ( .A(\os1/sigQout2 ), .B(n573), .Q(sig_fsm_start_R) );
  NOR21 U1839 ( .A(i_FIFO[0]), .B(n807), .Q(N159) );
  NOR21 U1840 ( .A(k_FIFO[0]), .B(n808), .Q(N191) );
  NOR21 U1841 ( .A(\os2/sigQout2 ), .B(n574), .Q(sig_fsm_start_W) );
  NAND22 U1842 ( .A(n876), .B(currentState[3]), .Q(n123) );
  INV3 U1843 ( .A(n114), .Q(n876) );
  INV3 U1844 ( .A(n910), .Q(n847) );
  NAND22 U1845 ( .A(n773), .B(\os1/sigQout1 ), .Q(n910) );
  INV3 U1846 ( .A(n912), .Q(n849) );
  NAND22 U1847 ( .A(n774), .B(\os2/sigQout1 ), .Q(n912) );
  NOR21 U1848 ( .A(n807), .B(n852), .Q(N918) );
  INV3 U1849 ( .A(inData), .Q(n852) );
  NOR40 U1850 ( .A(currentState[2]), .B(currentState[1]), .C(currentState[0]), 
        .D(n575), .Q(outDone) );
  BUF2 U1851 ( .A(inReset), .Q(n771) );
  BUF2 U1852 ( .A(inReset), .Q(n770) );
  BUF2 U1853 ( .A(inReset), .Q(n772) );
  BUF2 U1854 ( .A(inReset), .Q(n773) );
  BUF2 U1855 ( .A(inReset), .Q(n790) );
  BUF2 U1856 ( .A(inReset), .Q(n791) );
  BUF2 U1857 ( .A(inReset), .Q(n792) );
  BUF2 U1858 ( .A(inReset), .Q(n793) );
  BUF2 U1859 ( .A(inReset), .Q(n794) );
  BUF2 U1860 ( .A(inReset), .Q(n795) );
  BUF2 U1861 ( .A(inReset), .Q(n796) );
  BUF2 U1862 ( .A(inReset), .Q(n797) );
  BUF2 U1863 ( .A(inReset), .Q(n798) );
  BUF2 U1864 ( .A(inReset), .Q(n799) );
  BUF2 U1865 ( .A(inReset), .Q(n800) );
  BUF2 U1866 ( .A(inReset), .Q(n801) );
  BUF2 U1867 ( .A(inReset), .Q(n802) );
  BUF2 U1868 ( .A(inReset), .Q(n803) );
  BUF2 U1869 ( .A(inReset), .Q(n804) );
  BUF2 U1870 ( .A(inReset), .Q(n805) );
  BUF2 U1871 ( .A(inReset), .Q(n781) );
  BUF2 U1872 ( .A(inReset), .Q(n780) );
  BUF2 U1873 ( .A(inReset), .Q(n779) );
  BUF2 U1874 ( .A(inReset), .Q(n777) );
  BUF2 U1875 ( .A(inReset), .Q(n776) );
  BUF2 U1876 ( .A(inReset), .Q(n775) );
  BUF2 U1877 ( .A(inReset), .Q(n778) );
  BUF2 U1878 ( .A(inReset), .Q(n782) );
  BUF2 U1879 ( .A(inReset), .Q(n783) );
  BUF2 U1880 ( .A(inReset), .Q(n784) );
  BUF2 U1881 ( .A(inReset), .Q(n785) );
  BUF2 U1882 ( .A(inReset), .Q(n786) );
  BUF2 U1883 ( .A(inReset), .Q(n787) );
  BUF2 U1884 ( .A(inReset), .Q(n788) );
  BUF2 U1885 ( .A(inReset), .Q(n789) );
  BUF2 U1886 ( .A(inReset), .Q(n774) );
  BUF2 U1887 ( .A(inReset), .Q(n806) );
  INV3 U1888 ( .A(n911), .Q(n848) );
  NAND22 U1889 ( .A(n773), .B(inWriteEnable), .Q(n911) );
  INV3 U1890 ( .A(\os1/dff1/n2 ), .Q(n850) );
  NAND22 U1891 ( .A(n774), .B(inReadEnable), .Q(\os1/dff1/n2 ) );
  OAI212 U1892 ( .A(outReadCount[2]), .B(n553), .C(n888), .Q(n891) );
  OAI212 U1893 ( .A(outReadCount[6]), .B(n564), .C(n897), .Q(n903) );
endmodule

