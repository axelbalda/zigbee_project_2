
module inFIFO ( inClock, inReset, inReadEnable, inWriteEnable, inData, 
        outWriteCount, outReadCount, outReadError, outWriteError, outFull, 
        outEmpty, outAlmostEmpty, outAlmostFull, outDone, outData );
  input [3:0] inData;
  output [7:0] outWriteCount;
  output [6:0] outReadCount;
  input inClock, inReset, inReadEnable, inWriteEnable;
  output outReadError, outWriteError, outFull, outEmpty, outAlmostEmpty,
         outAlmostFull, outDone, outData;
  wire   N38, N40, N41, N42, N43, N44, N45, sig_fsm_start_W, N47, N48, N49,
         N50, N119, N120, N121, N122, N123, N124, N126, N127, N128, N129, N130,
         N131, N133, N134, N135, N136, N137, N138, N139, N140, N143, N144,
         N145, N146, N147, N148, N149, N190, N196, N199, \FIFO[127][3] ,
         \FIFO[127][2] , \FIFO[127][1] , \FIFO[127][0] , \FIFO[126][3] ,
         \FIFO[126][2] , \FIFO[126][1] , \FIFO[126][0] , \FIFO[125][3] ,
         \FIFO[125][2] , \FIFO[125][1] , \FIFO[125][0] , \FIFO[124][3] ,
         \FIFO[124][2] , \FIFO[124][1] , \FIFO[124][0] , \FIFO[123][3] ,
         \FIFO[123][2] , \FIFO[123][1] , \FIFO[123][0] , \FIFO[122][3] ,
         \FIFO[122][2] , \FIFO[122][1] , \FIFO[122][0] , \FIFO[121][3] ,
         \FIFO[121][2] , \FIFO[121][1] , \FIFO[121][0] , \FIFO[120][3] ,
         \FIFO[120][2] , \FIFO[120][1] , \FIFO[120][0] , \FIFO[119][3] ,
         \FIFO[119][2] , \FIFO[119][1] , \FIFO[119][0] , \FIFO[118][3] ,
         \FIFO[118][2] , \FIFO[118][1] , \FIFO[118][0] , \FIFO[117][3] ,
         \FIFO[117][2] , \FIFO[117][1] , \FIFO[117][0] , \FIFO[116][3] ,
         \FIFO[116][2] , \FIFO[116][1] , \FIFO[116][0] , \FIFO[115][3] ,
         \FIFO[115][2] , \FIFO[115][1] , \FIFO[115][0] , \FIFO[114][3] ,
         \FIFO[114][2] , \FIFO[114][1] , \FIFO[114][0] , \FIFO[113][3] ,
         \FIFO[113][2] , \FIFO[113][1] , \FIFO[113][0] , \FIFO[112][3] ,
         \FIFO[112][2] , \FIFO[112][1] , \FIFO[112][0] , \FIFO[111][3] ,
         \FIFO[111][2] , \FIFO[111][1] , \FIFO[111][0] , \FIFO[110][3] ,
         \FIFO[110][2] , \FIFO[110][1] , \FIFO[110][0] , \FIFO[109][3] ,
         \FIFO[109][2] , \FIFO[109][1] , \FIFO[109][0] , \FIFO[108][3] ,
         \FIFO[108][2] , \FIFO[108][1] , \FIFO[108][0] , \FIFO[107][3] ,
         \FIFO[107][2] , \FIFO[107][1] , \FIFO[107][0] , \FIFO[106][3] ,
         \FIFO[106][2] , \FIFO[106][1] , \FIFO[106][0] , \FIFO[105][3] ,
         \FIFO[105][2] , \FIFO[105][1] , \FIFO[105][0] , \FIFO[104][3] ,
         \FIFO[104][2] , \FIFO[104][1] , \FIFO[104][0] , \FIFO[103][3] ,
         \FIFO[103][2] , \FIFO[103][1] , \FIFO[103][0] , \FIFO[102][3] ,
         \FIFO[102][2] , \FIFO[102][1] , \FIFO[102][0] , \FIFO[101][3] ,
         \FIFO[101][2] , \FIFO[101][1] , \FIFO[101][0] , \FIFO[100][3] ,
         \FIFO[100][2] , \FIFO[100][1] , \FIFO[100][0] , \FIFO[99][3] ,
         \FIFO[99][2] , \FIFO[99][1] , \FIFO[99][0] , \FIFO[98][3] ,
         \FIFO[98][2] , \FIFO[98][1] , \FIFO[98][0] , \FIFO[97][3] ,
         \FIFO[97][2] , \FIFO[97][1] , \FIFO[97][0] , \FIFO[96][3] ,
         \FIFO[96][2] , \FIFO[96][1] , \FIFO[96][0] , \FIFO[95][3] ,
         \FIFO[95][2] , \FIFO[95][1] , \FIFO[95][0] , \FIFO[94][3] ,
         \FIFO[94][2] , \FIFO[94][1] , \FIFO[94][0] , \FIFO[93][3] ,
         \FIFO[93][2] , \FIFO[93][1] , \FIFO[93][0] , \FIFO[92][3] ,
         \FIFO[92][2] , \FIFO[92][1] , \FIFO[92][0] , \FIFO[91][3] ,
         \FIFO[91][2] , \FIFO[91][1] , \FIFO[91][0] , \FIFO[90][3] ,
         \FIFO[90][2] , \FIFO[90][1] , \FIFO[90][0] , \FIFO[89][3] ,
         \FIFO[89][2] , \FIFO[89][1] , \FIFO[89][0] , \FIFO[88][3] ,
         \FIFO[88][2] , \FIFO[88][1] , \FIFO[88][0] , \FIFO[87][3] ,
         \FIFO[87][2] , \FIFO[87][1] , \FIFO[87][0] , \FIFO[86][3] ,
         \FIFO[86][2] , \FIFO[86][1] , \FIFO[86][0] , \FIFO[85][3] ,
         \FIFO[85][2] , \FIFO[85][1] , \FIFO[85][0] , \FIFO[84][3] ,
         \FIFO[84][2] , \FIFO[84][1] , \FIFO[84][0] , \FIFO[83][3] ,
         \FIFO[83][2] , \FIFO[83][1] , \FIFO[83][0] , \FIFO[82][3] ,
         \FIFO[82][2] , \FIFO[82][1] , \FIFO[82][0] , \FIFO[81][3] ,
         \FIFO[81][2] , \FIFO[81][1] , \FIFO[81][0] , \FIFO[80][3] ,
         \FIFO[80][2] , \FIFO[80][1] , \FIFO[80][0] , \FIFO[79][3] ,
         \FIFO[79][2] , \FIFO[79][1] , \FIFO[79][0] , \FIFO[78][3] ,
         \FIFO[78][2] , \FIFO[78][1] , \FIFO[78][0] , \FIFO[77][3] ,
         \FIFO[77][2] , \FIFO[77][1] , \FIFO[77][0] , \FIFO[76][3] ,
         \FIFO[76][2] , \FIFO[76][1] , \FIFO[76][0] , \FIFO[75][3] ,
         \FIFO[75][2] , \FIFO[75][1] , \FIFO[75][0] , \FIFO[74][3] ,
         \FIFO[74][2] , \FIFO[74][1] , \FIFO[74][0] , \FIFO[73][3] ,
         \FIFO[73][2] , \FIFO[73][1] , \FIFO[73][0] , \FIFO[72][3] ,
         \FIFO[72][2] , \FIFO[72][1] , \FIFO[72][0] , \FIFO[71][3] ,
         \FIFO[71][2] , \FIFO[71][1] , \FIFO[71][0] , \FIFO[70][3] ,
         \FIFO[70][2] , \FIFO[70][1] , \FIFO[70][0] , \FIFO[69][3] ,
         \FIFO[69][2] , \FIFO[69][1] , \FIFO[69][0] , \FIFO[68][3] ,
         \FIFO[68][2] , \FIFO[68][1] , \FIFO[68][0] , \FIFO[67][3] ,
         \FIFO[67][2] , \FIFO[67][1] , \FIFO[67][0] , \FIFO[66][3] ,
         \FIFO[66][2] , \FIFO[66][1] , \FIFO[66][0] , \FIFO[65][3] ,
         \FIFO[65][2] , \FIFO[65][1] , \FIFO[65][0] , \FIFO[64][3] ,
         \FIFO[64][2] , \FIFO[64][1] , \FIFO[64][0] , \FIFO[63][3] ,
         \FIFO[63][2] , \FIFO[63][1] , \FIFO[63][0] , \FIFO[62][3] ,
         \FIFO[62][2] , \FIFO[62][1] , \FIFO[62][0] , \FIFO[61][3] ,
         \FIFO[61][2] , \FIFO[61][1] , \FIFO[61][0] , \FIFO[60][3] ,
         \FIFO[60][2] , \FIFO[60][1] , \FIFO[60][0] , \FIFO[59][3] ,
         \FIFO[59][2] , \FIFO[59][1] , \FIFO[59][0] , \FIFO[58][3] ,
         \FIFO[58][2] , \FIFO[58][1] , \FIFO[58][0] , \FIFO[57][3] ,
         \FIFO[57][2] , \FIFO[57][1] , \FIFO[57][0] , \FIFO[56][3] ,
         \FIFO[56][2] , \FIFO[56][1] , \FIFO[56][0] , \FIFO[55][3] ,
         \FIFO[55][2] , \FIFO[55][1] , \FIFO[55][0] , \FIFO[54][3] ,
         \FIFO[54][2] , \FIFO[54][1] , \FIFO[54][0] , \FIFO[53][3] ,
         \FIFO[53][2] , \FIFO[53][1] , \FIFO[53][0] , \FIFO[52][3] ,
         \FIFO[52][2] , \FIFO[52][1] , \FIFO[52][0] , \FIFO[51][3] ,
         \FIFO[51][2] , \FIFO[51][1] , \FIFO[51][0] , \FIFO[50][3] ,
         \FIFO[50][2] , \FIFO[50][1] , \FIFO[50][0] , \FIFO[49][3] ,
         \FIFO[49][2] , \FIFO[49][1] , \FIFO[49][0] , \FIFO[48][3] ,
         \FIFO[48][2] , \FIFO[48][1] , \FIFO[48][0] , \FIFO[47][3] ,
         \FIFO[47][2] , \FIFO[47][1] , \FIFO[47][0] , \FIFO[46][3] ,
         \FIFO[46][2] , \FIFO[46][1] , \FIFO[46][0] , \FIFO[45][3] ,
         \FIFO[45][2] , \FIFO[45][1] , \FIFO[45][0] , \FIFO[44][3] ,
         \FIFO[44][2] , \FIFO[44][1] , \FIFO[44][0] , \FIFO[43][3] ,
         \FIFO[43][2] , \FIFO[43][1] , \FIFO[43][0] , \FIFO[42][3] ,
         \FIFO[42][2] , \FIFO[42][1] , \FIFO[42][0] , \FIFO[41][3] ,
         \FIFO[41][2] , \FIFO[41][1] , \FIFO[41][0] , \FIFO[40][3] ,
         \FIFO[40][2] , \FIFO[40][1] , \FIFO[40][0] , \FIFO[39][3] ,
         \FIFO[39][2] , \FIFO[39][1] , \FIFO[39][0] , \FIFO[38][3] ,
         \FIFO[38][2] , \FIFO[38][1] , \FIFO[38][0] , \FIFO[37][3] ,
         \FIFO[37][2] , \FIFO[37][1] , \FIFO[37][0] , \FIFO[36][3] ,
         \FIFO[36][2] , \FIFO[36][1] , \FIFO[36][0] , \FIFO[35][3] ,
         \FIFO[35][2] , \FIFO[35][1] , \FIFO[35][0] , \FIFO[34][3] ,
         \FIFO[34][2] , \FIFO[34][1] , \FIFO[34][0] , \FIFO[33][3] ,
         \FIFO[33][2] , \FIFO[33][1] , \FIFO[33][0] , \FIFO[32][3] ,
         \FIFO[32][2] , \FIFO[32][1] , \FIFO[32][0] , \FIFO[31][3] ,
         \FIFO[31][2] , \FIFO[31][1] , \FIFO[31][0] , \FIFO[30][3] ,
         \FIFO[30][2] , \FIFO[30][1] , \FIFO[30][0] , \FIFO[29][3] ,
         \FIFO[29][2] , \FIFO[29][1] , \FIFO[29][0] , \FIFO[28][3] ,
         \FIFO[28][2] , \FIFO[28][1] , \FIFO[28][0] , \FIFO[27][3] ,
         \FIFO[27][2] , \FIFO[27][1] , \FIFO[27][0] , \FIFO[26][3] ,
         \FIFO[26][2] , \FIFO[26][1] , \FIFO[26][0] , \FIFO[25][3] ,
         \FIFO[25][2] , \FIFO[25][1] , \FIFO[25][0] , \FIFO[24][3] ,
         \FIFO[24][2] , \FIFO[24][1] , \FIFO[24][0] , \FIFO[23][3] ,
         \FIFO[23][2] , \FIFO[23][1] , \FIFO[23][0] , \FIFO[22][3] ,
         \FIFO[22][2] , \FIFO[22][1] , \FIFO[22][0] , \FIFO[21][3] ,
         \FIFO[21][2] , \FIFO[21][1] , \FIFO[21][0] , \FIFO[20][3] ,
         \FIFO[20][2] , \FIFO[20][1] , \FIFO[20][0] , \FIFO[19][3] ,
         \FIFO[19][2] , \FIFO[19][1] , \FIFO[19][0] , \FIFO[18][3] ,
         \FIFO[18][2] , \FIFO[18][1] , \FIFO[18][0] , \FIFO[17][3] ,
         \FIFO[17][2] , \FIFO[17][1] , \FIFO[17][0] , \FIFO[16][3] ,
         \FIFO[16][2] , \FIFO[16][1] , \FIFO[16][0] , \FIFO[15][3] ,
         \FIFO[15][2] , \FIFO[15][1] , \FIFO[15][0] , \FIFO[14][3] ,
         \FIFO[14][2] , \FIFO[14][1] , \FIFO[14][0] , \FIFO[13][3] ,
         \FIFO[13][2] , \FIFO[13][1] , \FIFO[13][0] , \FIFO[12][3] ,
         \FIFO[12][2] , \FIFO[12][1] , \FIFO[12][0] , \FIFO[11][3] ,
         \FIFO[11][2] , \FIFO[11][1] , \FIFO[11][0] , \FIFO[10][3] ,
         \FIFO[10][2] , \FIFO[10][1] , \FIFO[10][0] , \FIFO[9][3] ,
         \FIFO[9][2] , \FIFO[9][1] , \FIFO[9][0] , \FIFO[8][3] , \FIFO[8][2] ,
         \FIFO[8][1] , \FIFO[8][0] , \FIFO[7][3] , \FIFO[7][2] , \FIFO[7][1] ,
         \FIFO[7][0] , \FIFO[6][3] , \FIFO[6][2] , \FIFO[6][1] , \FIFO[6][0] ,
         \FIFO[5][3] , \FIFO[5][2] , \FIFO[5][1] , \FIFO[5][0] , \FIFO[4][3] ,
         \FIFO[4][2] , \FIFO[4][1] , \FIFO[4][0] , \FIFO[3][3] , \FIFO[3][2] ,
         \FIFO[3][1] , \FIFO[3][0] , \FIFO[2][3] , \FIFO[2][2] , \FIFO[2][1] ,
         \FIFO[2][0] , \FIFO[1][3] , \FIFO[1][2] , \FIFO[1][1] , \FIFO[1][0] ,
         \FIFO[0][3] , \FIFO[0][2] , \FIFO[0][1] , \FIFO[0][0] , N200, N201,
         N202, N203, N204, N212, N213, N214, N215, N216, N225, N226, N227,
         N228, N229, N230, N231, N375, N381, N382, N390, N391, N392, N393,
         N396, N397, N398, N399, N400, N401, N402, N403, N404, N405, N406,
         N407, N408, N409, N410, N411, N412, N413, N414, N415, N416, N417,
         N418, N419, N420, N422, N423, N424, N425, N426, N427, N428, N429,
         N430, N431, N432, N433, N434, N435, N436, N437, N438, N439, N440,
         N441, N442, N443, N444, N445, N446, N448, N449, N450, N451, N452,
         N453, N454, N455, N456, N457, N458, N459, N460, N461, N462, N463,
         N464, N465, N466, N467, N468, N469, N470, N471, N472, N474, N475,
         N476, N477, N478, N479, N480, N481, N482, N483, N484, N485, N486,
         N487, N488, N489, N490, N491, N492, N493, N494, N495, N496, N497,
         N498, N499, N500, N501, N502, N503, N504, N505, N506, N507, N508,
         N509, N510, N511, N512, N513, N514, N515, N516, N517, N518, N519,
         N520, N521, N522, N524, N525, N526, N527, N528, N530, N532, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120,
         n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
         n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
         n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175,
         n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186,
         n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197,
         n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208,
         n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         \os1/sigQout1 , \os1/dff1/n2 , \os2/sigQout2 , \os2/sigQout1 , n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715;
  wire   [3:0] currentState;
  wire   [6:0] j_FIFO;
  wire   [6:2] \add_357/carry ;
  wire   [7:2] \add_263/carry ;
  wire   [6:2] \add_253/carry ;
  wire   [6:2] \add_252/carry ;
  wire   [8:0] \r96/carry ;
  assign outFull = N375;
  assign outAlmostEmpty = N390;
  assign outEmpty = N391;

  OAI222 U73 ( .A(n665), .B(n657), .C(n133), .D(n505), .Q(n132) );
  OAI212 U95 ( .A(n146), .B(n601), .C(n621), .Q(N49) );
  OAI212 U119 ( .A(n159), .B(n601), .C(n621), .Q(N48) );
  OAI222 U120 ( .A(currentState[0]), .B(n161), .C(n601), .D(n162), .Q(n160) );
  ADD22 \add_357/U1_1_1  ( .A(j_FIFO[1]), .B(j_FIFO[0]), .CO(
        \add_357/carry [2]), .S(N212) );
  ADD22 \add_357/U1_1_2  ( .A(j_FIFO[2]), .B(\add_357/carry [2]), .CO(
        \add_357/carry [3]), .S(N213) );
  ADD22 \add_357/U1_1_3  ( .A(j_FIFO[3]), .B(\add_357/carry [3]), .CO(
        \add_357/carry [4]), .S(N214) );
  ADD22 \add_357/U1_1_4  ( .A(j_FIFO[4]), .B(\add_357/carry [4]), .CO(
        \add_357/carry [5]), .S(N215) );
  ADD22 \add_357/U1_1_5  ( .A(j_FIFO[5]), .B(\add_357/carry [5]), .CO(
        \add_357/carry [6]), .S(N216) );
  ADD22 \add_263/U1_1_1  ( .A(outWriteCount[1]), .B(outWriteCount[0]), .CO(
        \add_263/carry [2]), .S(N143) );
  ADD22 \add_263/U1_1_2  ( .A(outWriteCount[2]), .B(\add_263/carry [2]), .CO(
        \add_263/carry [3]), .S(N144) );
  ADD22 \add_263/U1_1_3  ( .A(outWriteCount[3]), .B(\add_263/carry [3]), .CO(
        \add_263/carry [4]), .S(N145) );
  ADD22 \add_263/U1_1_4  ( .A(outWriteCount[4]), .B(\add_263/carry [4]), .CO(
        \add_263/carry [5]), .S(N146) );
  ADD22 \add_263/U1_1_5  ( .A(outWriteCount[5]), .B(\add_263/carry [5]), .CO(
        \add_263/carry [6]), .S(N147) );
  ADD22 \add_263/U1_1_6  ( .A(outWriteCount[6]), .B(\add_263/carry [6]), .CO(
        \add_263/carry [7]), .S(N148) );
  ADD22 \add_253/U1_1_1  ( .A(n523), .B(n620), .CO(\add_253/carry [2]), .S(
        N126) );
  ADD22 \add_253/U1_1_2  ( .A(n522), .B(\add_253/carry [2]), .CO(
        \add_253/carry [3]), .S(N127) );
  ADD22 \add_253/U1_1_3  ( .A(n605), .B(\add_253/carry [3]), .CO(
        \add_253/carry [4]), .S(N128) );
  ADD22 \add_253/U1_1_4  ( .A(n521), .B(\add_253/carry [4]), .CO(
        \add_253/carry [5]), .S(N129) );
  ADD22 \add_253/U1_1_5  ( .A(n520), .B(\add_253/carry [5]), .CO(
        \add_253/carry [6]), .S(N130) );
  ADD22 \add_252/U1_1_1  ( .A(outReadCount[1]), .B(outReadCount[0]), .CO(
        \add_252/carry [2]), .S(N119) );
  ADD22 \add_252/U1_1_2  ( .A(outReadCount[2]), .B(\add_252/carry [2]), .CO(
        \add_252/carry [3]), .S(N120) );
  ADD22 \add_252/U1_1_3  ( .A(outReadCount[3]), .B(\add_252/carry [3]), .CO(
        \add_252/carry [4]), .S(N121) );
  ADD22 \add_252/U1_1_4  ( .A(outReadCount[4]), .B(\add_252/carry [4]), .CO(
        \add_252/carry [5]), .S(N122) );
  ADD22 \add_252/U1_1_5  ( .A(outReadCount[5]), .B(\add_252/carry [5]), .CO(
        \add_252/carry [6]), .S(N123) );
  ADD32 \r96/U2_1  ( .A(outWriteCount[1]), .B(n493), .CI(\r96/carry [1]), .CO(
        \r96/carry [2]), .S(N134) );
  ADD32 \r96/U2_2  ( .A(outWriteCount[2]), .B(n495), .CI(\r96/carry [2]), .CO(
        \r96/carry [3]), .S(N135) );
  ADD32 \r96/U2_3  ( .A(outWriteCount[3]), .B(n498), .CI(\r96/carry [3]), .CO(
        \r96/carry [4]), .S(N136) );
  ADD32 \r96/U2_4  ( .A(outWriteCount[4]), .B(n496), .CI(\r96/carry [4]), .CO(
        \r96/carry [5]), .S(N137) );
  ADD32 \r96/U2_5  ( .A(outWriteCount[5]), .B(n497), .CI(\r96/carry [5]), .CO(
        \r96/carry [6]), .S(N138) );
  ADD32 \r96/U2_6  ( .A(outWriteCount[6]), .B(n501), .CI(\r96/carry [6]), .CO(
        \r96/carry [7]), .S(N139) );
  DF3 sigEnableCounter_reg ( .D(N196), .C(inClock), .QN(n510) );
  DF3 \currentState_reg[3]  ( .D(N50), .C(inClock), .Q(currentState[3]), .QN(
        n489) );
  DF3 \currentState_reg[0]  ( .D(N47), .C(inClock), .Q(currentState[0]), .QN(
        n505) );
  DF3 \currentState_reg[1]  ( .D(N48), .C(inClock), .Q(currentState[1]), .QN(
        n513) );
  DF3 \currentState_reg[2]  ( .D(N49), .C(inClock), .Q(currentState[2]) );
  DF3 \os1/dff1/s_qout_reg  ( .D(n640), .C(inClock), .Q(\os1/sigQout1 ) );
  DF3 \os2/dff2/s_qout_reg  ( .D(n639), .C(inClock), .Q(\os2/sigQout2 ) );
  DF3 \os2/dff1/s_qout_reg  ( .D(n638), .C(inClock), .Q(\os2/sigQout1 ), .QN(
        n515) );
  DF3 \os1/dff2/s_qout_reg  ( .D(n637), .C(inClock), .QN(n518) );
  DFE1 \k_FIFO_reg[0]  ( .D(n648), .E(N199), .C(inClock), .Q(N44), .QN(n514)
         );
  DFE1 \k_FIFO_reg[1]  ( .D(N190), .E(N199), .C(inClock), .Q(N45), .QN(n492)
         );
  DFE1 \FIFO_reg[126][3]  ( .D(n576), .E(N398), .C(inClock), .Q(\FIFO[126][3] ) );
  DFE1 \FIFO_reg[126][2]  ( .D(n560), .E(N398), .C(inClock), .Q(\FIFO[126][2] ) );
  DFE1 \FIFO_reg[126][1]  ( .D(n544), .E(N398), .C(inClock), .Q(\FIFO[126][1] ) );
  DFE1 \FIFO_reg[126][0]  ( .D(n528), .E(N398), .C(inClock), .Q(\FIFO[126][0] ) );
  DFE1 \FIFO_reg[122][3]  ( .D(n576), .E(N402), .C(inClock), .Q(\FIFO[122][3] ) );
  DFE1 \FIFO_reg[122][2]  ( .D(n560), .E(N402), .C(inClock), .Q(\FIFO[122][2] ) );
  DFE1 \FIFO_reg[122][1]  ( .D(n544), .E(N402), .C(inClock), .Q(\FIFO[122][1] ) );
  DFE1 \FIFO_reg[122][0]  ( .D(n528), .E(N402), .C(inClock), .Q(\FIFO[122][0] ) );
  DFE1 \FIFO_reg[118][3]  ( .D(n577), .E(N406), .C(inClock), .Q(\FIFO[118][3] ) );
  DFE1 \FIFO_reg[118][2]  ( .D(n561), .E(N406), .C(inClock), .Q(\FIFO[118][2] ) );
  DFE1 \FIFO_reg[118][1]  ( .D(n545), .E(N406), .C(inClock), .Q(\FIFO[118][1] ) );
  DFE1 \FIFO_reg[118][0]  ( .D(n529), .E(N406), .C(inClock), .Q(\FIFO[118][0] ) );
  DFE1 \FIFO_reg[114][3]  ( .D(n577), .E(N410), .C(inClock), .Q(\FIFO[114][3] ) );
  DFE1 \FIFO_reg[114][2]  ( .D(n561), .E(N410), .C(inClock), .Q(\FIFO[114][2] ) );
  DFE1 \FIFO_reg[114][1]  ( .D(n545), .E(N410), .C(inClock), .Q(\FIFO[114][1] ) );
  DFE1 \FIFO_reg[114][0]  ( .D(n529), .E(N410), .C(inClock), .Q(\FIFO[114][0] ) );
  DFE1 \FIFO_reg[110][3]  ( .D(n578), .E(N414), .C(inClock), .Q(\FIFO[110][3] ) );
  DFE1 \FIFO_reg[110][2]  ( .D(n562), .E(N414), .C(inClock), .Q(\FIFO[110][2] ) );
  DFE1 \FIFO_reg[110][1]  ( .D(n546), .E(N414), .C(inClock), .Q(\FIFO[110][1] ) );
  DFE1 \FIFO_reg[110][0]  ( .D(n530), .E(N414), .C(inClock), .Q(\FIFO[110][0] ) );
  DFE1 \FIFO_reg[106][3]  ( .D(n578), .E(N418), .C(inClock), .Q(\FIFO[106][3] ) );
  DFE1 \FIFO_reg[106][2]  ( .D(n562), .E(N418), .C(inClock), .Q(\FIFO[106][2] ) );
  DFE1 \FIFO_reg[106][1]  ( .D(n546), .E(N418), .C(inClock), .Q(\FIFO[106][1] ) );
  DFE1 \FIFO_reg[106][0]  ( .D(n530), .E(N418), .C(inClock), .Q(\FIFO[106][0] ) );
  DFE1 \FIFO_reg[102][3]  ( .D(n579), .E(N423), .C(inClock), .Q(\FIFO[102][3] ) );
  DFE1 \FIFO_reg[102][2]  ( .D(n563), .E(N423), .C(inClock), .Q(\FIFO[102][2] ) );
  DFE1 \FIFO_reg[102][1]  ( .D(n547), .E(N423), .C(inClock), .Q(\FIFO[102][1] ) );
  DFE1 \FIFO_reg[102][0]  ( .D(n531), .E(N423), .C(inClock), .Q(\FIFO[102][0] ) );
  DFE1 \FIFO_reg[98][3]  ( .D(n579), .E(N427), .C(inClock), .Q(\FIFO[98][3] )
         );
  DFE1 \FIFO_reg[98][2]  ( .D(n563), .E(N427), .C(inClock), .Q(\FIFO[98][2] )
         );
  DFE1 \FIFO_reg[98][1]  ( .D(n547), .E(N427), .C(inClock), .Q(\FIFO[98][1] )
         );
  DFE1 \FIFO_reg[98][0]  ( .D(n531), .E(N427), .C(inClock), .Q(\FIFO[98][0] )
         );
  DFE1 \FIFO_reg[94][3]  ( .D(n580), .E(N431), .C(inClock), .Q(\FIFO[94][3] )
         );
  DFE1 \FIFO_reg[94][2]  ( .D(n564), .E(N431), .C(inClock), .Q(\FIFO[94][2] )
         );
  DFE1 \FIFO_reg[94][1]  ( .D(n548), .E(N431), .C(inClock), .Q(\FIFO[94][1] )
         );
  DFE1 \FIFO_reg[94][0]  ( .D(n532), .E(N431), .C(inClock), .Q(\FIFO[94][0] )
         );
  DFE1 \FIFO_reg[90][3]  ( .D(n580), .E(N435), .C(inClock), .Q(\FIFO[90][3] )
         );
  DFE1 \FIFO_reg[90][2]  ( .D(n564), .E(N435), .C(inClock), .Q(\FIFO[90][2] )
         );
  DFE1 \FIFO_reg[90][1]  ( .D(n548), .E(N435), .C(inClock), .Q(\FIFO[90][1] )
         );
  DFE1 \FIFO_reg[90][0]  ( .D(n532), .E(N435), .C(inClock), .Q(\FIFO[90][0] )
         );
  DFE1 \FIFO_reg[86][3]  ( .D(n581), .E(N439), .C(inClock), .Q(\FIFO[86][3] )
         );
  DFE1 \FIFO_reg[86][2]  ( .D(n565), .E(N439), .C(inClock), .Q(\FIFO[86][2] )
         );
  DFE1 \FIFO_reg[86][1]  ( .D(n549), .E(N439), .C(inClock), .Q(\FIFO[86][1] )
         );
  DFE1 \FIFO_reg[86][0]  ( .D(n533), .E(N439), .C(inClock), .Q(\FIFO[86][0] )
         );
  DFE1 \FIFO_reg[82][3]  ( .D(n581), .E(N443), .C(inClock), .Q(\FIFO[82][3] )
         );
  DFE1 \FIFO_reg[82][2]  ( .D(n565), .E(N443), .C(inClock), .Q(\FIFO[82][2] )
         );
  DFE1 \FIFO_reg[82][1]  ( .D(n549), .E(N443), .C(inClock), .Q(\FIFO[82][1] )
         );
  DFE1 \FIFO_reg[82][0]  ( .D(n533), .E(N443), .C(inClock), .Q(\FIFO[82][0] )
         );
  DFE1 \FIFO_reg[78][3]  ( .D(n582), .E(N448), .C(inClock), .Q(\FIFO[78][3] )
         );
  DFE1 \FIFO_reg[78][2]  ( .D(n566), .E(N448), .C(inClock), .Q(\FIFO[78][2] )
         );
  DFE1 \FIFO_reg[78][1]  ( .D(n550), .E(N448), .C(inClock), .Q(\FIFO[78][1] )
         );
  DFE1 \FIFO_reg[78][0]  ( .D(n534), .E(N448), .C(inClock), .Q(\FIFO[78][0] )
         );
  DFE1 \FIFO_reg[74][3]  ( .D(n582), .E(N452), .C(inClock), .Q(\FIFO[74][3] )
         );
  DFE1 \FIFO_reg[74][2]  ( .D(n566), .E(N452), .C(inClock), .Q(\FIFO[74][2] )
         );
  DFE1 \FIFO_reg[74][1]  ( .D(n550), .E(N452), .C(inClock), .Q(\FIFO[74][1] )
         );
  DFE1 \FIFO_reg[74][0]  ( .D(n534), .E(N452), .C(inClock), .Q(\FIFO[74][0] )
         );
  DFE1 \FIFO_reg[70][3]  ( .D(n583), .E(N456), .C(inClock), .Q(\FIFO[70][3] )
         );
  DFE1 \FIFO_reg[70][2]  ( .D(n567), .E(N456), .C(inClock), .Q(\FIFO[70][2] )
         );
  DFE1 \FIFO_reg[70][1]  ( .D(n551), .E(N456), .C(inClock), .Q(\FIFO[70][1] )
         );
  DFE1 \FIFO_reg[70][0]  ( .D(n535), .E(N456), .C(inClock), .Q(\FIFO[70][0] )
         );
  DFE1 \FIFO_reg[66][3]  ( .D(n583), .E(N460), .C(inClock), .Q(\FIFO[66][3] )
         );
  DFE1 \FIFO_reg[66][2]  ( .D(n567), .E(N460), .C(inClock), .Q(\FIFO[66][2] )
         );
  DFE1 \FIFO_reg[66][1]  ( .D(n551), .E(N460), .C(inClock), .Q(\FIFO[66][1] )
         );
  DFE1 \FIFO_reg[66][0]  ( .D(n535), .E(N460), .C(inClock), .Q(\FIFO[66][0] )
         );
  DFE1 \FIFO_reg[62][3]  ( .D(n584), .E(N464), .C(inClock), .Q(\FIFO[62][3] )
         );
  DFE1 \FIFO_reg[62][2]  ( .D(n568), .E(N464), .C(inClock), .Q(\FIFO[62][2] )
         );
  DFE1 \FIFO_reg[62][1]  ( .D(n552), .E(N464), .C(inClock), .Q(\FIFO[62][1] )
         );
  DFE1 \FIFO_reg[62][0]  ( .D(n536), .E(N464), .C(inClock), .Q(\FIFO[62][0] )
         );
  DFE1 \FIFO_reg[58][3]  ( .D(n584), .E(N468), .C(inClock), .Q(\FIFO[58][3] )
         );
  DFE1 \FIFO_reg[58][2]  ( .D(n568), .E(N468), .C(inClock), .Q(\FIFO[58][2] )
         );
  DFE1 \FIFO_reg[58][1]  ( .D(n552), .E(N468), .C(inClock), .Q(\FIFO[58][1] )
         );
  DFE1 \FIFO_reg[58][0]  ( .D(n536), .E(N468), .C(inClock), .Q(\FIFO[58][0] )
         );
  DFE1 \FIFO_reg[54][3]  ( .D(n585), .E(N472), .C(inClock), .Q(\FIFO[54][3] )
         );
  DFE1 \FIFO_reg[54][2]  ( .D(n569), .E(N472), .C(inClock), .Q(\FIFO[54][2] )
         );
  DFE1 \FIFO_reg[54][1]  ( .D(n553), .E(N472), .C(inClock), .Q(\FIFO[54][1] )
         );
  DFE1 \FIFO_reg[54][0]  ( .D(n537), .E(N472), .C(inClock), .Q(\FIFO[54][0] )
         );
  DFE1 \FIFO_reg[50][3]  ( .D(n585), .E(N477), .C(inClock), .Q(\FIFO[50][3] )
         );
  DFE1 \FIFO_reg[50][2]  ( .D(n569), .E(N477), .C(inClock), .Q(\FIFO[50][2] )
         );
  DFE1 \FIFO_reg[50][1]  ( .D(n553), .E(N477), .C(inClock), .Q(\FIFO[50][1] )
         );
  DFE1 \FIFO_reg[50][0]  ( .D(n537), .E(N477), .C(inClock), .Q(\FIFO[50][0] )
         );
  DFE1 \FIFO_reg[46][3]  ( .D(n586), .E(N481), .C(inClock), .Q(\FIFO[46][3] )
         );
  DFE1 \FIFO_reg[46][2]  ( .D(n570), .E(N481), .C(inClock), .Q(\FIFO[46][2] )
         );
  DFE1 \FIFO_reg[46][1]  ( .D(n554), .E(N481), .C(inClock), .Q(\FIFO[46][1] )
         );
  DFE1 \FIFO_reg[46][0]  ( .D(n538), .E(N481), .C(inClock), .Q(\FIFO[46][0] )
         );
  DFE1 \FIFO_reg[42][3]  ( .D(n586), .E(N485), .C(inClock), .Q(\FIFO[42][3] )
         );
  DFE1 \FIFO_reg[42][2]  ( .D(n570), .E(N485), .C(inClock), .Q(\FIFO[42][2] )
         );
  DFE1 \FIFO_reg[42][1]  ( .D(n554), .E(N485), .C(inClock), .Q(\FIFO[42][1] )
         );
  DFE1 \FIFO_reg[42][0]  ( .D(n538), .E(N485), .C(inClock), .Q(\FIFO[42][0] )
         );
  DFE1 \FIFO_reg[38][3]  ( .D(n587), .E(N489), .C(inClock), .Q(\FIFO[38][3] )
         );
  DFE1 \FIFO_reg[38][2]  ( .D(n571), .E(N489), .C(inClock), .Q(\FIFO[38][2] )
         );
  DFE1 \FIFO_reg[38][1]  ( .D(n555), .E(N489), .C(inClock), .Q(\FIFO[38][1] )
         );
  DFE1 \FIFO_reg[38][0]  ( .D(n539), .E(N489), .C(inClock), .Q(\FIFO[38][0] )
         );
  DFE1 \FIFO_reg[34][3]  ( .D(n587), .E(N493), .C(inClock), .Q(\FIFO[34][3] )
         );
  DFE1 \FIFO_reg[34][2]  ( .D(n571), .E(N493), .C(inClock), .Q(\FIFO[34][2] )
         );
  DFE1 \FIFO_reg[34][1]  ( .D(n555), .E(N493), .C(inClock), .Q(\FIFO[34][1] )
         );
  DFE1 \FIFO_reg[34][0]  ( .D(n539), .E(N493), .C(inClock), .Q(\FIFO[34][0] )
         );
  DFE1 \FIFO_reg[30][3]  ( .D(n588), .E(N497), .C(inClock), .Q(\FIFO[30][3] )
         );
  DFE1 \FIFO_reg[30][2]  ( .D(n572), .E(N497), .C(inClock), .Q(\FIFO[30][2] )
         );
  DFE1 \FIFO_reg[30][1]  ( .D(n556), .E(N497), .C(inClock), .Q(\FIFO[30][1] )
         );
  DFE1 \FIFO_reg[30][0]  ( .D(n540), .E(N497), .C(inClock), .Q(\FIFO[30][0] )
         );
  DFE1 \FIFO_reg[26][3]  ( .D(n588), .E(N501), .C(inClock), .Q(\FIFO[26][3] )
         );
  DFE1 \FIFO_reg[26][2]  ( .D(n572), .E(N501), .C(inClock), .Q(\FIFO[26][2] )
         );
  DFE1 \FIFO_reg[26][1]  ( .D(n556), .E(N501), .C(inClock), .Q(\FIFO[26][1] )
         );
  DFE1 \FIFO_reg[26][0]  ( .D(n540), .E(N501), .C(inClock), .Q(\FIFO[26][0] )
         );
  DFE1 \FIFO_reg[22][3]  ( .D(n589), .E(N505), .C(inClock), .Q(\FIFO[22][3] )
         );
  DFE1 \FIFO_reg[22][2]  ( .D(n573), .E(N505), .C(inClock), .Q(\FIFO[22][2] )
         );
  DFE1 \FIFO_reg[22][1]  ( .D(n557), .E(N505), .C(inClock), .Q(\FIFO[22][1] )
         );
  DFE1 \FIFO_reg[22][0]  ( .D(n541), .E(N505), .C(inClock), .Q(\FIFO[22][0] )
         );
  DFE1 \FIFO_reg[18][3]  ( .D(n589), .E(N509), .C(inClock), .Q(\FIFO[18][3] )
         );
  DFE1 \FIFO_reg[18][2]  ( .D(n573), .E(N509), .C(inClock), .Q(\FIFO[18][2] )
         );
  DFE1 \FIFO_reg[18][1]  ( .D(n557), .E(N509), .C(inClock), .Q(\FIFO[18][1] )
         );
  DFE1 \FIFO_reg[18][0]  ( .D(n541), .E(N509), .C(inClock), .Q(\FIFO[18][0] )
         );
  DFE1 \FIFO_reg[14][3]  ( .D(n590), .E(N513), .C(inClock), .Q(\FIFO[14][3] )
         );
  DFE1 \FIFO_reg[14][2]  ( .D(n574), .E(N513), .C(inClock), .Q(\FIFO[14][2] )
         );
  DFE1 \FIFO_reg[14][1]  ( .D(n558), .E(N513), .C(inClock), .Q(\FIFO[14][1] )
         );
  DFE1 \FIFO_reg[14][0]  ( .D(n542), .E(N513), .C(inClock), .Q(\FIFO[14][0] )
         );
  DFE1 \FIFO_reg[10][3]  ( .D(n590), .E(N517), .C(inClock), .Q(\FIFO[10][3] )
         );
  DFE1 \FIFO_reg[10][2]  ( .D(n574), .E(N517), .C(inClock), .Q(\FIFO[10][2] )
         );
  DFE1 \FIFO_reg[10][1]  ( .D(n558), .E(N517), .C(inClock), .Q(\FIFO[10][1] )
         );
  DFE1 \FIFO_reg[10][0]  ( .D(n542), .E(N517), .C(inClock), .Q(\FIFO[10][0] )
         );
  DFE1 \FIFO_reg[6][3]  ( .D(n591), .E(N521), .C(inClock), .Q(\FIFO[6][3] ) );
  DFE1 \FIFO_reg[6][2]  ( .D(n575), .E(N521), .C(inClock), .Q(\FIFO[6][2] ) );
  DFE1 \FIFO_reg[6][1]  ( .D(n559), .E(N521), .C(inClock), .Q(\FIFO[6][1] ) );
  DFE1 \FIFO_reg[6][0]  ( .D(n543), .E(N521), .C(inClock), .Q(\FIFO[6][0] ) );
  DFE1 \FIFO_reg[2][3]  ( .D(n591), .E(N526), .C(inClock), .Q(\FIFO[2][3] ) );
  DFE1 \FIFO_reg[2][2]  ( .D(n575), .E(N526), .C(inClock), .Q(\FIFO[2][2] ) );
  DFE1 \FIFO_reg[2][1]  ( .D(n559), .E(N526), .C(inClock), .Q(\FIFO[2][1] ) );
  DFE1 \FIFO_reg[2][0]  ( .D(n543), .E(N526), .C(inClock), .Q(\FIFO[2][0] ) );
  DFE1 \FIFO_reg[127][3]  ( .D(n576), .E(N397), .C(inClock), .Q(\FIFO[127][3] ) );
  DFE1 \FIFO_reg[127][2]  ( .D(n560), .E(N397), .C(inClock), .Q(\FIFO[127][2] ) );
  DFE1 \FIFO_reg[127][1]  ( .D(n544), .E(N397), .C(inClock), .Q(\FIFO[127][1] ) );
  DFE1 \FIFO_reg[127][0]  ( .D(n528), .E(N397), .C(inClock), .Q(\FIFO[127][0] ) );
  DFE1 \FIFO_reg[125][3]  ( .D(n576), .E(N399), .C(inClock), .Q(\FIFO[125][3] ) );
  DFE1 \FIFO_reg[125][2]  ( .D(n560), .E(N399), .C(inClock), .Q(\FIFO[125][2] ) );
  DFE1 \FIFO_reg[125][1]  ( .D(n544), .E(N399), .C(inClock), .Q(\FIFO[125][1] ) );
  DFE1 \FIFO_reg[125][0]  ( .D(n528), .E(N399), .C(inClock), .Q(\FIFO[125][0] ) );
  DFE1 \FIFO_reg[124][3]  ( .D(n576), .E(N400), .C(inClock), .Q(\FIFO[124][3] ) );
  DFE1 \FIFO_reg[124][2]  ( .D(n560), .E(N400), .C(inClock), .Q(\FIFO[124][2] ) );
  DFE1 \FIFO_reg[124][1]  ( .D(n544), .E(N400), .C(inClock), .Q(\FIFO[124][1] ) );
  DFE1 \FIFO_reg[124][0]  ( .D(n528), .E(N400), .C(inClock), .Q(\FIFO[124][0] ) );
  DFE1 \FIFO_reg[123][3]  ( .D(n576), .E(N401), .C(inClock), .Q(\FIFO[123][3] ) );
  DFE1 \FIFO_reg[123][2]  ( .D(n560), .E(N401), .C(inClock), .Q(\FIFO[123][2] ) );
  DFE1 \FIFO_reg[123][1]  ( .D(n544), .E(N401), .C(inClock), .Q(\FIFO[123][1] ) );
  DFE1 \FIFO_reg[123][0]  ( .D(n528), .E(N401), .C(inClock), .Q(\FIFO[123][0] ) );
  DFE1 \FIFO_reg[121][3]  ( .D(n576), .E(N403), .C(inClock), .Q(\FIFO[121][3] ) );
  DFE1 \FIFO_reg[121][2]  ( .D(n560), .E(N403), .C(inClock), .Q(\FIFO[121][2] ) );
  DFE1 \FIFO_reg[121][1]  ( .D(n544), .E(N403), .C(inClock), .Q(\FIFO[121][1] ) );
  DFE1 \FIFO_reg[121][0]  ( .D(n528), .E(N403), .C(inClock), .Q(\FIFO[121][0] ) );
  DFE1 \FIFO_reg[120][3]  ( .D(n576), .E(N404), .C(inClock), .Q(\FIFO[120][3] ) );
  DFE1 \FIFO_reg[120][2]  ( .D(n560), .E(N404), .C(inClock), .Q(\FIFO[120][2] ) );
  DFE1 \FIFO_reg[120][1]  ( .D(n544), .E(N404), .C(inClock), .Q(\FIFO[120][1] ) );
  DFE1 \FIFO_reg[120][0]  ( .D(n528), .E(N404), .C(inClock), .Q(\FIFO[120][0] ) );
  DFE1 \FIFO_reg[119][3]  ( .D(n577), .E(N405), .C(inClock), .Q(\FIFO[119][3] ) );
  DFE1 \FIFO_reg[119][2]  ( .D(n561), .E(N405), .C(inClock), .Q(\FIFO[119][2] ) );
  DFE1 \FIFO_reg[119][1]  ( .D(n545), .E(N405), .C(inClock), .Q(\FIFO[119][1] ) );
  DFE1 \FIFO_reg[119][0]  ( .D(n529), .E(N405), .C(inClock), .Q(\FIFO[119][0] ) );
  DFE1 \FIFO_reg[117][3]  ( .D(n577), .E(N407), .C(inClock), .Q(\FIFO[117][3] ) );
  DFE1 \FIFO_reg[117][2]  ( .D(n561), .E(N407), .C(inClock), .Q(\FIFO[117][2] ) );
  DFE1 \FIFO_reg[117][1]  ( .D(n545), .E(N407), .C(inClock), .Q(\FIFO[117][1] ) );
  DFE1 \FIFO_reg[117][0]  ( .D(n529), .E(N407), .C(inClock), .Q(\FIFO[117][0] ) );
  DFE1 \FIFO_reg[116][3]  ( .D(n577), .E(N408), .C(inClock), .Q(\FIFO[116][3] ) );
  DFE1 \FIFO_reg[116][2]  ( .D(n561), .E(N408), .C(inClock), .Q(\FIFO[116][2] ) );
  DFE1 \FIFO_reg[116][1]  ( .D(n545), .E(N408), .C(inClock), .Q(\FIFO[116][1] ) );
  DFE1 \FIFO_reg[116][0]  ( .D(n529), .E(N408), .C(inClock), .Q(\FIFO[116][0] ) );
  DFE1 \FIFO_reg[115][3]  ( .D(n577), .E(N409), .C(inClock), .Q(\FIFO[115][3] ) );
  DFE1 \FIFO_reg[115][2]  ( .D(n561), .E(N409), .C(inClock), .Q(\FIFO[115][2] ) );
  DFE1 \FIFO_reg[115][1]  ( .D(n545), .E(N409), .C(inClock), .Q(\FIFO[115][1] ) );
  DFE1 \FIFO_reg[115][0]  ( .D(n529), .E(N409), .C(inClock), .Q(\FIFO[115][0] ) );
  DFE1 \FIFO_reg[113][3]  ( .D(n577), .E(N411), .C(inClock), .Q(\FIFO[113][3] ) );
  DFE1 \FIFO_reg[113][2]  ( .D(n561), .E(N411), .C(inClock), .Q(\FIFO[113][2] ) );
  DFE1 \FIFO_reg[113][1]  ( .D(n545), .E(N411), .C(inClock), .Q(\FIFO[113][1] ) );
  DFE1 \FIFO_reg[113][0]  ( .D(n529), .E(N411), .C(inClock), .Q(\FIFO[113][0] ) );
  DFE1 \FIFO_reg[112][3]  ( .D(n577), .E(N412), .C(inClock), .Q(\FIFO[112][3] ) );
  DFE1 \FIFO_reg[112][2]  ( .D(n561), .E(N412), .C(inClock), .Q(\FIFO[112][2] ) );
  DFE1 \FIFO_reg[112][1]  ( .D(n545), .E(N412), .C(inClock), .Q(\FIFO[112][1] ) );
  DFE1 \FIFO_reg[112][0]  ( .D(n529), .E(N412), .C(inClock), .Q(\FIFO[112][0] ) );
  DFE1 \FIFO_reg[111][3]  ( .D(n578), .E(N413), .C(inClock), .Q(\FIFO[111][3] ) );
  DFE1 \FIFO_reg[111][2]  ( .D(n562), .E(N413), .C(inClock), .Q(\FIFO[111][2] ) );
  DFE1 \FIFO_reg[111][1]  ( .D(n546), .E(N413), .C(inClock), .Q(\FIFO[111][1] ) );
  DFE1 \FIFO_reg[111][0]  ( .D(n530), .E(N413), .C(inClock), .Q(\FIFO[111][0] ) );
  DFE1 \FIFO_reg[109][3]  ( .D(n578), .E(N415), .C(inClock), .Q(\FIFO[109][3] ) );
  DFE1 \FIFO_reg[109][2]  ( .D(n562), .E(N415), .C(inClock), .Q(\FIFO[109][2] ) );
  DFE1 \FIFO_reg[109][1]  ( .D(n546), .E(N415), .C(inClock), .Q(\FIFO[109][1] ) );
  DFE1 \FIFO_reg[109][0]  ( .D(n530), .E(N415), .C(inClock), .Q(\FIFO[109][0] ) );
  DFE1 \FIFO_reg[108][3]  ( .D(n578), .E(N416), .C(inClock), .Q(\FIFO[108][3] ) );
  DFE1 \FIFO_reg[108][2]  ( .D(n562), .E(N416), .C(inClock), .Q(\FIFO[108][2] ) );
  DFE1 \FIFO_reg[108][1]  ( .D(n546), .E(N416), .C(inClock), .Q(\FIFO[108][1] ) );
  DFE1 \FIFO_reg[108][0]  ( .D(n530), .E(N416), .C(inClock), .Q(\FIFO[108][0] ) );
  DFE1 \FIFO_reg[107][3]  ( .D(n578), .E(N417), .C(inClock), .Q(\FIFO[107][3] ) );
  DFE1 \FIFO_reg[107][2]  ( .D(n562), .E(N417), .C(inClock), .Q(\FIFO[107][2] ) );
  DFE1 \FIFO_reg[107][1]  ( .D(n546), .E(N417), .C(inClock), .Q(\FIFO[107][1] ) );
  DFE1 \FIFO_reg[107][0]  ( .D(n530), .E(N417), .C(inClock), .Q(\FIFO[107][0] ) );
  DFE1 \FIFO_reg[105][3]  ( .D(n578), .E(N419), .C(inClock), .Q(\FIFO[105][3] ) );
  DFE1 \FIFO_reg[105][2]  ( .D(n562), .E(N419), .C(inClock), .Q(\FIFO[105][2] ) );
  DFE1 \FIFO_reg[105][1]  ( .D(n546), .E(N419), .C(inClock), .Q(\FIFO[105][1] ) );
  DFE1 \FIFO_reg[105][0]  ( .D(n530), .E(N419), .C(inClock), .Q(\FIFO[105][0] ) );
  DFE1 \FIFO_reg[104][3]  ( .D(n578), .E(N420), .C(inClock), .Q(\FIFO[104][3] ) );
  DFE1 \FIFO_reg[104][2]  ( .D(n562), .E(N420), .C(inClock), .Q(\FIFO[104][2] ) );
  DFE1 \FIFO_reg[104][1]  ( .D(n546), .E(N420), .C(inClock), .Q(\FIFO[104][1] ) );
  DFE1 \FIFO_reg[104][0]  ( .D(n530), .E(N420), .C(inClock), .Q(\FIFO[104][0] ) );
  DFE1 \FIFO_reg[103][3]  ( .D(n579), .E(N422), .C(inClock), .Q(\FIFO[103][3] ) );
  DFE1 \FIFO_reg[103][2]  ( .D(n563), .E(N422), .C(inClock), .Q(\FIFO[103][2] ) );
  DFE1 \FIFO_reg[103][1]  ( .D(n547), .E(N422), .C(inClock), .Q(\FIFO[103][1] ) );
  DFE1 \FIFO_reg[103][0]  ( .D(n531), .E(N422), .C(inClock), .Q(\FIFO[103][0] ) );
  DFE1 \FIFO_reg[101][3]  ( .D(n579), .E(N424), .C(inClock), .Q(\FIFO[101][3] ) );
  DFE1 \FIFO_reg[101][2]  ( .D(n563), .E(N424), .C(inClock), .Q(\FIFO[101][2] ) );
  DFE1 \FIFO_reg[101][1]  ( .D(n547), .E(N424), .C(inClock), .Q(\FIFO[101][1] ) );
  DFE1 \FIFO_reg[101][0]  ( .D(n531), .E(N424), .C(inClock), .Q(\FIFO[101][0] ) );
  DFE1 \FIFO_reg[100][3]  ( .D(n579), .E(N425), .C(inClock), .Q(\FIFO[100][3] ) );
  DFE1 \FIFO_reg[100][2]  ( .D(n563), .E(N425), .C(inClock), .Q(\FIFO[100][2] ) );
  DFE1 \FIFO_reg[100][1]  ( .D(n547), .E(N425), .C(inClock), .Q(\FIFO[100][1] ) );
  DFE1 \FIFO_reg[100][0]  ( .D(n531), .E(N425), .C(inClock), .Q(\FIFO[100][0] ) );
  DFE1 \FIFO_reg[99][3]  ( .D(n579), .E(N426), .C(inClock), .Q(\FIFO[99][3] )
         );
  DFE1 \FIFO_reg[99][2]  ( .D(n563), .E(N426), .C(inClock), .Q(\FIFO[99][2] )
         );
  DFE1 \FIFO_reg[99][1]  ( .D(n547), .E(N426), .C(inClock), .Q(\FIFO[99][1] )
         );
  DFE1 \FIFO_reg[99][0]  ( .D(n531), .E(N426), .C(inClock), .Q(\FIFO[99][0] )
         );
  DFE1 \FIFO_reg[97][3]  ( .D(n579), .E(N428), .C(inClock), .Q(\FIFO[97][3] )
         );
  DFE1 \FIFO_reg[97][2]  ( .D(n563), .E(N428), .C(inClock), .Q(\FIFO[97][2] )
         );
  DFE1 \FIFO_reg[97][1]  ( .D(n547), .E(N428), .C(inClock), .Q(\FIFO[97][1] )
         );
  DFE1 \FIFO_reg[97][0]  ( .D(n531), .E(N428), .C(inClock), .Q(\FIFO[97][0] )
         );
  DFE1 \FIFO_reg[96][3]  ( .D(n579), .E(N429), .C(inClock), .Q(\FIFO[96][3] )
         );
  DFE1 \FIFO_reg[96][2]  ( .D(n563), .E(N429), .C(inClock), .Q(\FIFO[96][2] )
         );
  DFE1 \FIFO_reg[96][1]  ( .D(n547), .E(N429), .C(inClock), .Q(\FIFO[96][1] )
         );
  DFE1 \FIFO_reg[96][0]  ( .D(n531), .E(N429), .C(inClock), .Q(\FIFO[96][0] )
         );
  DFE1 \FIFO_reg[95][3]  ( .D(n580), .E(N430), .C(inClock), .Q(\FIFO[95][3] )
         );
  DFE1 \FIFO_reg[95][2]  ( .D(n564), .E(N430), .C(inClock), .Q(\FIFO[95][2] )
         );
  DFE1 \FIFO_reg[95][1]  ( .D(n548), .E(N430), .C(inClock), .Q(\FIFO[95][1] )
         );
  DFE1 \FIFO_reg[95][0]  ( .D(n532), .E(N430), .C(inClock), .Q(\FIFO[95][0] )
         );
  DFE1 \FIFO_reg[93][3]  ( .D(n580), .E(N432), .C(inClock), .Q(\FIFO[93][3] )
         );
  DFE1 \FIFO_reg[93][2]  ( .D(n564), .E(N432), .C(inClock), .Q(\FIFO[93][2] )
         );
  DFE1 \FIFO_reg[93][1]  ( .D(n548), .E(N432), .C(inClock), .Q(\FIFO[93][1] )
         );
  DFE1 \FIFO_reg[93][0]  ( .D(n532), .E(N432), .C(inClock), .Q(\FIFO[93][0] )
         );
  DFE1 \FIFO_reg[92][3]  ( .D(n580), .E(N433), .C(inClock), .Q(\FIFO[92][3] )
         );
  DFE1 \FIFO_reg[92][2]  ( .D(n564), .E(N433), .C(inClock), .Q(\FIFO[92][2] )
         );
  DFE1 \FIFO_reg[92][1]  ( .D(n548), .E(N433), .C(inClock), .Q(\FIFO[92][1] )
         );
  DFE1 \FIFO_reg[92][0]  ( .D(n532), .E(N433), .C(inClock), .Q(\FIFO[92][0] )
         );
  DFE1 \FIFO_reg[91][3]  ( .D(n580), .E(N434), .C(inClock), .Q(\FIFO[91][3] )
         );
  DFE1 \FIFO_reg[91][2]  ( .D(n564), .E(N434), .C(inClock), .Q(\FIFO[91][2] )
         );
  DFE1 \FIFO_reg[91][1]  ( .D(n548), .E(N434), .C(inClock), .Q(\FIFO[91][1] )
         );
  DFE1 \FIFO_reg[91][0]  ( .D(n532), .E(N434), .C(inClock), .Q(\FIFO[91][0] )
         );
  DFE1 \FIFO_reg[89][3]  ( .D(n580), .E(N436), .C(inClock), .Q(\FIFO[89][3] )
         );
  DFE1 \FIFO_reg[89][2]  ( .D(n564), .E(N436), .C(inClock), .Q(\FIFO[89][2] )
         );
  DFE1 \FIFO_reg[89][1]  ( .D(n548), .E(N436), .C(inClock), .Q(\FIFO[89][1] )
         );
  DFE1 \FIFO_reg[89][0]  ( .D(n532), .E(N436), .C(inClock), .Q(\FIFO[89][0] )
         );
  DFE1 \FIFO_reg[88][3]  ( .D(n580), .E(N437), .C(inClock), .Q(\FIFO[88][3] )
         );
  DFE1 \FIFO_reg[88][2]  ( .D(n564), .E(N437), .C(inClock), .Q(\FIFO[88][2] )
         );
  DFE1 \FIFO_reg[88][1]  ( .D(n548), .E(N437), .C(inClock), .Q(\FIFO[88][1] )
         );
  DFE1 \FIFO_reg[88][0]  ( .D(n532), .E(N437), .C(inClock), .Q(\FIFO[88][0] )
         );
  DFE1 \FIFO_reg[87][3]  ( .D(n581), .E(N438), .C(inClock), .Q(\FIFO[87][3] )
         );
  DFE1 \FIFO_reg[87][2]  ( .D(n565), .E(N438), .C(inClock), .Q(\FIFO[87][2] )
         );
  DFE1 \FIFO_reg[87][1]  ( .D(n549), .E(N438), .C(inClock), .Q(\FIFO[87][1] )
         );
  DFE1 \FIFO_reg[87][0]  ( .D(n533), .E(N438), .C(inClock), .Q(\FIFO[87][0] )
         );
  DFE1 \FIFO_reg[85][3]  ( .D(n581), .E(N440), .C(inClock), .Q(\FIFO[85][3] )
         );
  DFE1 \FIFO_reg[85][2]  ( .D(n565), .E(N440), .C(inClock), .Q(\FIFO[85][2] )
         );
  DFE1 \FIFO_reg[85][1]  ( .D(n549), .E(N440), .C(inClock), .Q(\FIFO[85][1] )
         );
  DFE1 \FIFO_reg[85][0]  ( .D(n533), .E(N440), .C(inClock), .Q(\FIFO[85][0] )
         );
  DFE1 \FIFO_reg[84][3]  ( .D(n581), .E(N441), .C(inClock), .Q(\FIFO[84][3] )
         );
  DFE1 \FIFO_reg[84][2]  ( .D(n565), .E(N441), .C(inClock), .Q(\FIFO[84][2] )
         );
  DFE1 \FIFO_reg[84][1]  ( .D(n549), .E(N441), .C(inClock), .Q(\FIFO[84][1] )
         );
  DFE1 \FIFO_reg[84][0]  ( .D(n533), .E(N441), .C(inClock), .Q(\FIFO[84][0] )
         );
  DFE1 \FIFO_reg[83][3]  ( .D(n581), .E(N442), .C(inClock), .Q(\FIFO[83][3] )
         );
  DFE1 \FIFO_reg[83][2]  ( .D(n565), .E(N442), .C(inClock), .Q(\FIFO[83][2] )
         );
  DFE1 \FIFO_reg[83][1]  ( .D(n549), .E(N442), .C(inClock), .Q(\FIFO[83][1] )
         );
  DFE1 \FIFO_reg[83][0]  ( .D(n533), .E(N442), .C(inClock), .Q(\FIFO[83][0] )
         );
  DFE1 \FIFO_reg[81][3]  ( .D(n581), .E(N444), .C(inClock), .Q(\FIFO[81][3] )
         );
  DFE1 \FIFO_reg[81][2]  ( .D(n565), .E(N444), .C(inClock), .Q(\FIFO[81][2] )
         );
  DFE1 \FIFO_reg[81][1]  ( .D(n549), .E(N444), .C(inClock), .Q(\FIFO[81][1] )
         );
  DFE1 \FIFO_reg[81][0]  ( .D(n533), .E(N444), .C(inClock), .Q(\FIFO[81][0] )
         );
  DFE1 \FIFO_reg[80][3]  ( .D(n581), .E(N445), .C(inClock), .Q(\FIFO[80][3] )
         );
  DFE1 \FIFO_reg[80][2]  ( .D(n565), .E(N445), .C(inClock), .Q(\FIFO[80][2] )
         );
  DFE1 \FIFO_reg[80][1]  ( .D(n549), .E(N445), .C(inClock), .Q(\FIFO[80][1] )
         );
  DFE1 \FIFO_reg[80][0]  ( .D(n533), .E(N445), .C(inClock), .Q(\FIFO[80][0] )
         );
  DFE1 \FIFO_reg[79][3]  ( .D(n582), .E(N446), .C(inClock), .Q(\FIFO[79][3] )
         );
  DFE1 \FIFO_reg[79][2]  ( .D(n566), .E(N446), .C(inClock), .Q(\FIFO[79][2] )
         );
  DFE1 \FIFO_reg[79][1]  ( .D(n550), .E(N446), .C(inClock), .Q(\FIFO[79][1] )
         );
  DFE1 \FIFO_reg[79][0]  ( .D(n534), .E(N446), .C(inClock), .Q(\FIFO[79][0] )
         );
  DFE1 \FIFO_reg[77][3]  ( .D(n582), .E(N449), .C(inClock), .Q(\FIFO[77][3] )
         );
  DFE1 \FIFO_reg[77][2]  ( .D(n566), .E(N449), .C(inClock), .Q(\FIFO[77][2] )
         );
  DFE1 \FIFO_reg[77][1]  ( .D(n550), .E(N449), .C(inClock), .Q(\FIFO[77][1] )
         );
  DFE1 \FIFO_reg[77][0]  ( .D(n534), .E(N449), .C(inClock), .Q(\FIFO[77][0] )
         );
  DFE1 \FIFO_reg[76][3]  ( .D(n582), .E(N450), .C(inClock), .Q(\FIFO[76][3] )
         );
  DFE1 \FIFO_reg[76][2]  ( .D(n566), .E(N450), .C(inClock), .Q(\FIFO[76][2] )
         );
  DFE1 \FIFO_reg[76][1]  ( .D(n550), .E(N450), .C(inClock), .Q(\FIFO[76][1] )
         );
  DFE1 \FIFO_reg[76][0]  ( .D(n534), .E(N450), .C(inClock), .Q(\FIFO[76][0] )
         );
  DFE1 \FIFO_reg[75][3]  ( .D(n582), .E(N451), .C(inClock), .Q(\FIFO[75][3] )
         );
  DFE1 \FIFO_reg[75][2]  ( .D(n566), .E(N451), .C(inClock), .Q(\FIFO[75][2] )
         );
  DFE1 \FIFO_reg[75][1]  ( .D(n550), .E(N451), .C(inClock), .Q(\FIFO[75][1] )
         );
  DFE1 \FIFO_reg[75][0]  ( .D(n534), .E(N451), .C(inClock), .Q(\FIFO[75][0] )
         );
  DFE1 \FIFO_reg[73][3]  ( .D(n582), .E(N453), .C(inClock), .Q(\FIFO[73][3] )
         );
  DFE1 \FIFO_reg[73][2]  ( .D(n566), .E(N453), .C(inClock), .Q(\FIFO[73][2] )
         );
  DFE1 \FIFO_reg[73][1]  ( .D(n550), .E(N453), .C(inClock), .Q(\FIFO[73][1] )
         );
  DFE1 \FIFO_reg[73][0]  ( .D(n534), .E(N453), .C(inClock), .Q(\FIFO[73][0] )
         );
  DFE1 \FIFO_reg[72][3]  ( .D(n582), .E(N454), .C(inClock), .Q(\FIFO[72][3] )
         );
  DFE1 \FIFO_reg[72][2]  ( .D(n566), .E(N454), .C(inClock), .Q(\FIFO[72][2] )
         );
  DFE1 \FIFO_reg[72][1]  ( .D(n550), .E(N454), .C(inClock), .Q(\FIFO[72][1] )
         );
  DFE1 \FIFO_reg[72][0]  ( .D(n534), .E(N454), .C(inClock), .Q(\FIFO[72][0] )
         );
  DFE1 \FIFO_reg[71][3]  ( .D(n583), .E(N455), .C(inClock), .Q(\FIFO[71][3] )
         );
  DFE1 \FIFO_reg[71][2]  ( .D(n567), .E(N455), .C(inClock), .Q(\FIFO[71][2] )
         );
  DFE1 \FIFO_reg[71][1]  ( .D(n551), .E(N455), .C(inClock), .Q(\FIFO[71][1] )
         );
  DFE1 \FIFO_reg[71][0]  ( .D(n535), .E(N455), .C(inClock), .Q(\FIFO[71][0] )
         );
  DFE1 \FIFO_reg[69][3]  ( .D(n583), .E(N457), .C(inClock), .Q(\FIFO[69][3] )
         );
  DFE1 \FIFO_reg[69][2]  ( .D(n567), .E(N457), .C(inClock), .Q(\FIFO[69][2] )
         );
  DFE1 \FIFO_reg[69][1]  ( .D(n551), .E(N457), .C(inClock), .Q(\FIFO[69][1] )
         );
  DFE1 \FIFO_reg[69][0]  ( .D(n535), .E(N457), .C(inClock), .Q(\FIFO[69][0] )
         );
  DFE1 \FIFO_reg[68][3]  ( .D(n583), .E(N458), .C(inClock), .Q(\FIFO[68][3] )
         );
  DFE1 \FIFO_reg[68][2]  ( .D(n567), .E(N458), .C(inClock), .Q(\FIFO[68][2] )
         );
  DFE1 \FIFO_reg[68][1]  ( .D(n551), .E(N458), .C(inClock), .Q(\FIFO[68][1] )
         );
  DFE1 \FIFO_reg[68][0]  ( .D(n535), .E(N458), .C(inClock), .Q(\FIFO[68][0] )
         );
  DFE1 \FIFO_reg[67][3]  ( .D(n583), .E(N459), .C(inClock), .Q(\FIFO[67][3] )
         );
  DFE1 \FIFO_reg[67][2]  ( .D(n567), .E(N459), .C(inClock), .Q(\FIFO[67][2] )
         );
  DFE1 \FIFO_reg[67][1]  ( .D(n551), .E(N459), .C(inClock), .Q(\FIFO[67][1] )
         );
  DFE1 \FIFO_reg[67][0]  ( .D(n535), .E(N459), .C(inClock), .Q(\FIFO[67][0] )
         );
  DFE1 \FIFO_reg[65][3]  ( .D(n583), .E(N461), .C(inClock), .Q(\FIFO[65][3] )
         );
  DFE1 \FIFO_reg[65][2]  ( .D(n567), .E(N461), .C(inClock), .Q(\FIFO[65][2] )
         );
  DFE1 \FIFO_reg[65][1]  ( .D(n551), .E(N461), .C(inClock), .Q(\FIFO[65][1] )
         );
  DFE1 \FIFO_reg[65][0]  ( .D(n535), .E(N461), .C(inClock), .Q(\FIFO[65][0] )
         );
  DFE1 \FIFO_reg[64][3]  ( .D(n583), .E(N462), .C(inClock), .Q(\FIFO[64][3] )
         );
  DFE1 \FIFO_reg[64][2]  ( .D(n567), .E(N462), .C(inClock), .Q(\FIFO[64][2] )
         );
  DFE1 \FIFO_reg[64][1]  ( .D(n551), .E(N462), .C(inClock), .Q(\FIFO[64][1] )
         );
  DFE1 \FIFO_reg[64][0]  ( .D(n535), .E(N462), .C(inClock), .Q(\FIFO[64][0] )
         );
  DFE1 \FIFO_reg[63][3]  ( .D(n584), .E(N463), .C(inClock), .Q(\FIFO[63][3] )
         );
  DFE1 \FIFO_reg[63][2]  ( .D(n568), .E(N463), .C(inClock), .Q(\FIFO[63][2] )
         );
  DFE1 \FIFO_reg[63][1]  ( .D(n552), .E(N463), .C(inClock), .Q(\FIFO[63][1] )
         );
  DFE1 \FIFO_reg[63][0]  ( .D(n536), .E(N463), .C(inClock), .Q(\FIFO[63][0] )
         );
  DFE1 \FIFO_reg[61][3]  ( .D(n584), .E(N465), .C(inClock), .Q(\FIFO[61][3] )
         );
  DFE1 \FIFO_reg[61][2]  ( .D(n568), .E(N465), .C(inClock), .Q(\FIFO[61][2] )
         );
  DFE1 \FIFO_reg[61][1]  ( .D(n552), .E(N465), .C(inClock), .Q(\FIFO[61][1] )
         );
  DFE1 \FIFO_reg[61][0]  ( .D(n536), .E(N465), .C(inClock), .Q(\FIFO[61][0] )
         );
  DFE1 \FIFO_reg[60][3]  ( .D(n584), .E(N466), .C(inClock), .Q(\FIFO[60][3] )
         );
  DFE1 \FIFO_reg[60][2]  ( .D(n568), .E(N466), .C(inClock), .Q(\FIFO[60][2] )
         );
  DFE1 \FIFO_reg[60][1]  ( .D(n552), .E(N466), .C(inClock), .Q(\FIFO[60][1] )
         );
  DFE1 \FIFO_reg[60][0]  ( .D(n536), .E(N466), .C(inClock), .Q(\FIFO[60][0] )
         );
  DFE1 \FIFO_reg[59][3]  ( .D(n584), .E(N467), .C(inClock), .Q(\FIFO[59][3] )
         );
  DFE1 \FIFO_reg[59][2]  ( .D(n568), .E(N467), .C(inClock), .Q(\FIFO[59][2] )
         );
  DFE1 \FIFO_reg[59][1]  ( .D(n552), .E(N467), .C(inClock), .Q(\FIFO[59][1] )
         );
  DFE1 \FIFO_reg[59][0]  ( .D(n536), .E(N467), .C(inClock), .Q(\FIFO[59][0] )
         );
  DFE1 \FIFO_reg[57][3]  ( .D(n584), .E(N469), .C(inClock), .Q(\FIFO[57][3] )
         );
  DFE1 \FIFO_reg[57][2]  ( .D(n568), .E(N469), .C(inClock), .Q(\FIFO[57][2] )
         );
  DFE1 \FIFO_reg[57][1]  ( .D(n552), .E(N469), .C(inClock), .Q(\FIFO[57][1] )
         );
  DFE1 \FIFO_reg[57][0]  ( .D(n536), .E(N469), .C(inClock), .Q(\FIFO[57][0] )
         );
  DFE1 \FIFO_reg[56][3]  ( .D(n584), .E(N470), .C(inClock), .Q(\FIFO[56][3] )
         );
  DFE1 \FIFO_reg[56][2]  ( .D(n568), .E(N470), .C(inClock), .Q(\FIFO[56][2] )
         );
  DFE1 \FIFO_reg[56][1]  ( .D(n552), .E(N470), .C(inClock), .Q(\FIFO[56][1] )
         );
  DFE1 \FIFO_reg[56][0]  ( .D(n536), .E(N470), .C(inClock), .Q(\FIFO[56][0] )
         );
  DFE1 \FIFO_reg[55][3]  ( .D(n585), .E(N471), .C(inClock), .Q(\FIFO[55][3] )
         );
  DFE1 \FIFO_reg[55][2]  ( .D(n569), .E(N471), .C(inClock), .Q(\FIFO[55][2] )
         );
  DFE1 \FIFO_reg[55][1]  ( .D(n553), .E(N471), .C(inClock), .Q(\FIFO[55][1] )
         );
  DFE1 \FIFO_reg[55][0]  ( .D(n537), .E(N471), .C(inClock), .Q(\FIFO[55][0] )
         );
  DFE1 \FIFO_reg[53][3]  ( .D(n585), .E(N474), .C(inClock), .Q(\FIFO[53][3] )
         );
  DFE1 \FIFO_reg[53][2]  ( .D(n569), .E(N474), .C(inClock), .Q(\FIFO[53][2] )
         );
  DFE1 \FIFO_reg[53][1]  ( .D(n553), .E(N474), .C(inClock), .Q(\FIFO[53][1] )
         );
  DFE1 \FIFO_reg[53][0]  ( .D(n537), .E(N474), .C(inClock), .Q(\FIFO[53][0] )
         );
  DFE1 \FIFO_reg[52][3]  ( .D(n585), .E(N475), .C(inClock), .Q(\FIFO[52][3] )
         );
  DFE1 \FIFO_reg[52][2]  ( .D(n569), .E(N475), .C(inClock), .Q(\FIFO[52][2] )
         );
  DFE1 \FIFO_reg[52][1]  ( .D(n553), .E(N475), .C(inClock), .Q(\FIFO[52][1] )
         );
  DFE1 \FIFO_reg[52][0]  ( .D(n537), .E(N475), .C(inClock), .Q(\FIFO[52][0] )
         );
  DFE1 \FIFO_reg[51][3]  ( .D(n585), .E(N476), .C(inClock), .Q(\FIFO[51][3] )
         );
  DFE1 \FIFO_reg[51][2]  ( .D(n569), .E(N476), .C(inClock), .Q(\FIFO[51][2] )
         );
  DFE1 \FIFO_reg[51][1]  ( .D(n553), .E(N476), .C(inClock), .Q(\FIFO[51][1] )
         );
  DFE1 \FIFO_reg[51][0]  ( .D(n537), .E(N476), .C(inClock), .Q(\FIFO[51][0] )
         );
  DFE1 \FIFO_reg[49][3]  ( .D(n585), .E(N478), .C(inClock), .Q(\FIFO[49][3] )
         );
  DFE1 \FIFO_reg[49][2]  ( .D(n569), .E(N478), .C(inClock), .Q(\FIFO[49][2] )
         );
  DFE1 \FIFO_reg[49][1]  ( .D(n553), .E(N478), .C(inClock), .Q(\FIFO[49][1] )
         );
  DFE1 \FIFO_reg[49][0]  ( .D(n537), .E(N478), .C(inClock), .Q(\FIFO[49][0] )
         );
  DFE1 \FIFO_reg[48][3]  ( .D(n585), .E(N479), .C(inClock), .Q(\FIFO[48][3] )
         );
  DFE1 \FIFO_reg[48][2]  ( .D(n569), .E(N479), .C(inClock), .Q(\FIFO[48][2] )
         );
  DFE1 \FIFO_reg[48][1]  ( .D(n553), .E(N479), .C(inClock), .Q(\FIFO[48][1] )
         );
  DFE1 \FIFO_reg[48][0]  ( .D(n537), .E(N479), .C(inClock), .Q(\FIFO[48][0] )
         );
  DFE1 \FIFO_reg[47][3]  ( .D(n586), .E(N480), .C(inClock), .Q(\FIFO[47][3] )
         );
  DFE1 \FIFO_reg[47][2]  ( .D(n570), .E(N480), .C(inClock), .Q(\FIFO[47][2] )
         );
  DFE1 \FIFO_reg[47][1]  ( .D(n554), .E(N480), .C(inClock), .Q(\FIFO[47][1] )
         );
  DFE1 \FIFO_reg[47][0]  ( .D(n538), .E(N480), .C(inClock), .Q(\FIFO[47][0] )
         );
  DFE1 \FIFO_reg[45][3]  ( .D(n586), .E(N482), .C(inClock), .Q(\FIFO[45][3] )
         );
  DFE1 \FIFO_reg[45][2]  ( .D(n570), .E(N482), .C(inClock), .Q(\FIFO[45][2] )
         );
  DFE1 \FIFO_reg[45][1]  ( .D(n554), .E(N482), .C(inClock), .Q(\FIFO[45][1] )
         );
  DFE1 \FIFO_reg[45][0]  ( .D(n538), .E(N482), .C(inClock), .Q(\FIFO[45][0] )
         );
  DFE1 \FIFO_reg[44][3]  ( .D(n586), .E(N483), .C(inClock), .Q(\FIFO[44][3] )
         );
  DFE1 \FIFO_reg[44][2]  ( .D(n570), .E(N483), .C(inClock), .Q(\FIFO[44][2] )
         );
  DFE1 \FIFO_reg[44][1]  ( .D(n554), .E(N483), .C(inClock), .Q(\FIFO[44][1] )
         );
  DFE1 \FIFO_reg[44][0]  ( .D(n538), .E(N483), .C(inClock), .Q(\FIFO[44][0] )
         );
  DFE1 \FIFO_reg[43][3]  ( .D(n586), .E(N484), .C(inClock), .Q(\FIFO[43][3] )
         );
  DFE1 \FIFO_reg[43][2]  ( .D(n570), .E(N484), .C(inClock), .Q(\FIFO[43][2] )
         );
  DFE1 \FIFO_reg[43][1]  ( .D(n554), .E(N484), .C(inClock), .Q(\FIFO[43][1] )
         );
  DFE1 \FIFO_reg[43][0]  ( .D(n538), .E(N484), .C(inClock), .Q(\FIFO[43][0] )
         );
  DFE1 \FIFO_reg[41][3]  ( .D(n586), .E(N486), .C(inClock), .Q(\FIFO[41][3] )
         );
  DFE1 \FIFO_reg[41][2]  ( .D(n570), .E(N486), .C(inClock), .Q(\FIFO[41][2] )
         );
  DFE1 \FIFO_reg[41][1]  ( .D(n554), .E(N486), .C(inClock), .Q(\FIFO[41][1] )
         );
  DFE1 \FIFO_reg[41][0]  ( .D(n538), .E(N486), .C(inClock), .Q(\FIFO[41][0] )
         );
  DFE1 \FIFO_reg[40][3]  ( .D(n586), .E(N487), .C(inClock), .Q(\FIFO[40][3] )
         );
  DFE1 \FIFO_reg[40][2]  ( .D(n570), .E(N487), .C(inClock), .Q(\FIFO[40][2] )
         );
  DFE1 \FIFO_reg[40][1]  ( .D(n554), .E(N487), .C(inClock), .Q(\FIFO[40][1] )
         );
  DFE1 \FIFO_reg[40][0]  ( .D(n538), .E(N487), .C(inClock), .Q(\FIFO[40][0] )
         );
  DFE1 \FIFO_reg[39][3]  ( .D(n587), .E(N488), .C(inClock), .Q(\FIFO[39][3] )
         );
  DFE1 \FIFO_reg[39][2]  ( .D(n571), .E(N488), .C(inClock), .Q(\FIFO[39][2] )
         );
  DFE1 \FIFO_reg[39][1]  ( .D(n555), .E(N488), .C(inClock), .Q(\FIFO[39][1] )
         );
  DFE1 \FIFO_reg[39][0]  ( .D(n539), .E(N488), .C(inClock), .Q(\FIFO[39][0] )
         );
  DFE1 \FIFO_reg[37][3]  ( .D(n587), .E(N490), .C(inClock), .Q(\FIFO[37][3] )
         );
  DFE1 \FIFO_reg[37][2]  ( .D(n571), .E(N490), .C(inClock), .Q(\FIFO[37][2] )
         );
  DFE1 \FIFO_reg[37][1]  ( .D(n555), .E(N490), .C(inClock), .Q(\FIFO[37][1] )
         );
  DFE1 \FIFO_reg[37][0]  ( .D(n539), .E(N490), .C(inClock), .Q(\FIFO[37][0] )
         );
  DFE1 \FIFO_reg[36][3]  ( .D(n587), .E(N491), .C(inClock), .Q(\FIFO[36][3] )
         );
  DFE1 \FIFO_reg[36][2]  ( .D(n571), .E(N491), .C(inClock), .Q(\FIFO[36][2] )
         );
  DFE1 \FIFO_reg[36][1]  ( .D(n555), .E(N491), .C(inClock), .Q(\FIFO[36][1] )
         );
  DFE1 \FIFO_reg[36][0]  ( .D(n539), .E(N491), .C(inClock), .Q(\FIFO[36][0] )
         );
  DFE1 \FIFO_reg[35][3]  ( .D(n587), .E(N492), .C(inClock), .Q(\FIFO[35][3] )
         );
  DFE1 \FIFO_reg[35][2]  ( .D(n571), .E(N492), .C(inClock), .Q(\FIFO[35][2] )
         );
  DFE1 \FIFO_reg[35][1]  ( .D(n555), .E(N492), .C(inClock), .Q(\FIFO[35][1] )
         );
  DFE1 \FIFO_reg[35][0]  ( .D(n539), .E(N492), .C(inClock), .Q(\FIFO[35][0] )
         );
  DFE1 \FIFO_reg[33][3]  ( .D(n587), .E(N494), .C(inClock), .Q(\FIFO[33][3] )
         );
  DFE1 \FIFO_reg[33][2]  ( .D(n571), .E(N494), .C(inClock), .Q(\FIFO[33][2] )
         );
  DFE1 \FIFO_reg[33][1]  ( .D(n555), .E(N494), .C(inClock), .Q(\FIFO[33][1] )
         );
  DFE1 \FIFO_reg[33][0]  ( .D(n539), .E(N494), .C(inClock), .Q(\FIFO[33][0] )
         );
  DFE1 \FIFO_reg[32][3]  ( .D(n587), .E(N495), .C(inClock), .Q(\FIFO[32][3] )
         );
  DFE1 \FIFO_reg[32][2]  ( .D(n571), .E(N495), .C(inClock), .Q(\FIFO[32][2] )
         );
  DFE1 \FIFO_reg[32][1]  ( .D(n555), .E(N495), .C(inClock), .Q(\FIFO[32][1] )
         );
  DFE1 \FIFO_reg[32][0]  ( .D(n539), .E(N495), .C(inClock), .Q(\FIFO[32][0] )
         );
  DFE1 \FIFO_reg[31][3]  ( .D(n588), .E(N496), .C(inClock), .Q(\FIFO[31][3] )
         );
  DFE1 \FIFO_reg[31][2]  ( .D(n572), .E(N496), .C(inClock), .Q(\FIFO[31][2] )
         );
  DFE1 \FIFO_reg[31][1]  ( .D(n556), .E(N496), .C(inClock), .Q(\FIFO[31][1] )
         );
  DFE1 \FIFO_reg[31][0]  ( .D(n540), .E(N496), .C(inClock), .Q(\FIFO[31][0] )
         );
  DFE1 \FIFO_reg[29][3]  ( .D(n588), .E(N498), .C(inClock), .Q(\FIFO[29][3] )
         );
  DFE1 \FIFO_reg[29][2]  ( .D(n572), .E(N498), .C(inClock), .Q(\FIFO[29][2] )
         );
  DFE1 \FIFO_reg[29][1]  ( .D(n556), .E(N498), .C(inClock), .Q(\FIFO[29][1] )
         );
  DFE1 \FIFO_reg[29][0]  ( .D(n540), .E(N498), .C(inClock), .Q(\FIFO[29][0] )
         );
  DFE1 \FIFO_reg[28][3]  ( .D(n588), .E(N499), .C(inClock), .Q(\FIFO[28][3] )
         );
  DFE1 \FIFO_reg[28][2]  ( .D(n572), .E(N499), .C(inClock), .Q(\FIFO[28][2] )
         );
  DFE1 \FIFO_reg[28][1]  ( .D(n556), .E(N499), .C(inClock), .Q(\FIFO[28][1] )
         );
  DFE1 \FIFO_reg[28][0]  ( .D(n540), .E(N499), .C(inClock), .Q(\FIFO[28][0] )
         );
  DFE1 \FIFO_reg[27][3]  ( .D(n588), .E(N500), .C(inClock), .Q(\FIFO[27][3] )
         );
  DFE1 \FIFO_reg[27][2]  ( .D(n572), .E(N500), .C(inClock), .Q(\FIFO[27][2] )
         );
  DFE1 \FIFO_reg[27][1]  ( .D(n556), .E(N500), .C(inClock), .Q(\FIFO[27][1] )
         );
  DFE1 \FIFO_reg[27][0]  ( .D(n540), .E(N500), .C(inClock), .Q(\FIFO[27][0] )
         );
  DFE1 \FIFO_reg[25][3]  ( .D(n588), .E(N502), .C(inClock), .Q(\FIFO[25][3] )
         );
  DFE1 \FIFO_reg[25][2]  ( .D(n572), .E(N502), .C(inClock), .Q(\FIFO[25][2] )
         );
  DFE1 \FIFO_reg[25][1]  ( .D(n556), .E(N502), .C(inClock), .Q(\FIFO[25][1] )
         );
  DFE1 \FIFO_reg[25][0]  ( .D(n540), .E(N502), .C(inClock), .Q(\FIFO[25][0] )
         );
  DFE1 \FIFO_reg[24][3]  ( .D(n588), .E(N503), .C(inClock), .Q(\FIFO[24][3] )
         );
  DFE1 \FIFO_reg[24][2]  ( .D(n572), .E(N503), .C(inClock), .Q(\FIFO[24][2] )
         );
  DFE1 \FIFO_reg[24][1]  ( .D(n556), .E(N503), .C(inClock), .Q(\FIFO[24][1] )
         );
  DFE1 \FIFO_reg[24][0]  ( .D(n540), .E(N503), .C(inClock), .Q(\FIFO[24][0] )
         );
  DFE1 \FIFO_reg[23][3]  ( .D(n589), .E(N504), .C(inClock), .Q(\FIFO[23][3] )
         );
  DFE1 \FIFO_reg[23][2]  ( .D(n573), .E(N504), .C(inClock), .Q(\FIFO[23][2] )
         );
  DFE1 \FIFO_reg[23][1]  ( .D(n557), .E(N504), .C(inClock), .Q(\FIFO[23][1] )
         );
  DFE1 \FIFO_reg[23][0]  ( .D(n541), .E(N504), .C(inClock), .Q(\FIFO[23][0] )
         );
  DFE1 \FIFO_reg[21][3]  ( .D(n589), .E(N506), .C(inClock), .Q(\FIFO[21][3] )
         );
  DFE1 \FIFO_reg[21][2]  ( .D(n573), .E(N506), .C(inClock), .Q(\FIFO[21][2] )
         );
  DFE1 \FIFO_reg[21][1]  ( .D(n557), .E(N506), .C(inClock), .Q(\FIFO[21][1] )
         );
  DFE1 \FIFO_reg[21][0]  ( .D(n541), .E(N506), .C(inClock), .Q(\FIFO[21][0] )
         );
  DFE1 \FIFO_reg[20][3]  ( .D(n589), .E(N507), .C(inClock), .Q(\FIFO[20][3] )
         );
  DFE1 \FIFO_reg[20][2]  ( .D(n573), .E(N507), .C(inClock), .Q(\FIFO[20][2] )
         );
  DFE1 \FIFO_reg[20][1]  ( .D(n557), .E(N507), .C(inClock), .Q(\FIFO[20][1] )
         );
  DFE1 \FIFO_reg[20][0]  ( .D(n541), .E(N507), .C(inClock), .Q(\FIFO[20][0] )
         );
  DFE1 \FIFO_reg[19][3]  ( .D(n589), .E(N508), .C(inClock), .Q(\FIFO[19][3] )
         );
  DFE1 \FIFO_reg[19][2]  ( .D(n573), .E(N508), .C(inClock), .Q(\FIFO[19][2] )
         );
  DFE1 \FIFO_reg[19][1]  ( .D(n557), .E(N508), .C(inClock), .Q(\FIFO[19][1] )
         );
  DFE1 \FIFO_reg[19][0]  ( .D(n541), .E(N508), .C(inClock), .Q(\FIFO[19][0] )
         );
  DFE1 \FIFO_reg[17][3]  ( .D(n589), .E(N510), .C(inClock), .Q(\FIFO[17][3] )
         );
  DFE1 \FIFO_reg[17][2]  ( .D(n573), .E(N510), .C(inClock), .Q(\FIFO[17][2] )
         );
  DFE1 \FIFO_reg[17][1]  ( .D(n557), .E(N510), .C(inClock), .Q(\FIFO[17][1] )
         );
  DFE1 \FIFO_reg[17][0]  ( .D(n541), .E(N510), .C(inClock), .Q(\FIFO[17][0] )
         );
  DFE1 \FIFO_reg[16][3]  ( .D(n589), .E(N511), .C(inClock), .Q(\FIFO[16][3] )
         );
  DFE1 \FIFO_reg[16][2]  ( .D(n573), .E(N511), .C(inClock), .Q(\FIFO[16][2] )
         );
  DFE1 \FIFO_reg[16][1]  ( .D(n557), .E(N511), .C(inClock), .Q(\FIFO[16][1] )
         );
  DFE1 \FIFO_reg[16][0]  ( .D(n541), .E(N511), .C(inClock), .Q(\FIFO[16][0] )
         );
  DFE1 \FIFO_reg[15][3]  ( .D(n590), .E(N512), .C(inClock), .Q(\FIFO[15][3] )
         );
  DFE1 \FIFO_reg[15][2]  ( .D(n574), .E(N512), .C(inClock), .Q(\FIFO[15][2] )
         );
  DFE1 \FIFO_reg[15][1]  ( .D(n558), .E(N512), .C(inClock), .Q(\FIFO[15][1] )
         );
  DFE1 \FIFO_reg[15][0]  ( .D(n542), .E(N512), .C(inClock), .Q(\FIFO[15][0] )
         );
  DFE1 \FIFO_reg[13][3]  ( .D(n590), .E(N514), .C(inClock), .Q(\FIFO[13][3] )
         );
  DFE1 \FIFO_reg[13][2]  ( .D(n574), .E(N514), .C(inClock), .Q(\FIFO[13][2] )
         );
  DFE1 \FIFO_reg[13][1]  ( .D(n558), .E(N514), .C(inClock), .Q(\FIFO[13][1] )
         );
  DFE1 \FIFO_reg[13][0]  ( .D(n542), .E(N514), .C(inClock), .Q(\FIFO[13][0] )
         );
  DFE1 \FIFO_reg[12][3]  ( .D(n590), .E(N515), .C(inClock), .Q(\FIFO[12][3] )
         );
  DFE1 \FIFO_reg[12][2]  ( .D(n574), .E(N515), .C(inClock), .Q(\FIFO[12][2] )
         );
  DFE1 \FIFO_reg[12][1]  ( .D(n558), .E(N515), .C(inClock), .Q(\FIFO[12][1] )
         );
  DFE1 \FIFO_reg[12][0]  ( .D(n542), .E(N515), .C(inClock), .Q(\FIFO[12][0] )
         );
  DFE1 \FIFO_reg[11][3]  ( .D(n590), .E(N516), .C(inClock), .Q(\FIFO[11][3] )
         );
  DFE1 \FIFO_reg[11][2]  ( .D(n574), .E(N516), .C(inClock), .Q(\FIFO[11][2] )
         );
  DFE1 \FIFO_reg[11][1]  ( .D(n558), .E(N516), .C(inClock), .Q(\FIFO[11][1] )
         );
  DFE1 \FIFO_reg[11][0]  ( .D(n542), .E(N516), .C(inClock), .Q(\FIFO[11][0] )
         );
  DFE1 \FIFO_reg[9][3]  ( .D(n590), .E(N518), .C(inClock), .Q(\FIFO[9][3] ) );
  DFE1 \FIFO_reg[9][2]  ( .D(n574), .E(N518), .C(inClock), .Q(\FIFO[9][2] ) );
  DFE1 \FIFO_reg[9][1]  ( .D(n558), .E(N518), .C(inClock), .Q(\FIFO[9][1] ) );
  DFE1 \FIFO_reg[9][0]  ( .D(n542), .E(N518), .C(inClock), .Q(\FIFO[9][0] ) );
  DFE1 \FIFO_reg[8][3]  ( .D(n590), .E(N519), .C(inClock), .Q(\FIFO[8][3] ) );
  DFE1 \FIFO_reg[8][2]  ( .D(n574), .E(N519), .C(inClock), .Q(\FIFO[8][2] ) );
  DFE1 \FIFO_reg[8][1]  ( .D(n558), .E(N519), .C(inClock), .Q(\FIFO[8][1] ) );
  DFE1 \FIFO_reg[8][0]  ( .D(n542), .E(N519), .C(inClock), .Q(\FIFO[8][0] ) );
  DFE1 \FIFO_reg[7][3]  ( .D(n591), .E(N520), .C(inClock), .Q(\FIFO[7][3] ) );
  DFE1 \FIFO_reg[7][2]  ( .D(n575), .E(N520), .C(inClock), .Q(\FIFO[7][2] ) );
  DFE1 \FIFO_reg[7][1]  ( .D(n559), .E(N520), .C(inClock), .Q(\FIFO[7][1] ) );
  DFE1 \FIFO_reg[7][0]  ( .D(n543), .E(N520), .C(inClock), .Q(\FIFO[7][0] ) );
  DFE1 \FIFO_reg[5][3]  ( .D(n591), .E(N522), .C(inClock), .Q(\FIFO[5][3] ) );
  DFE1 \FIFO_reg[5][2]  ( .D(n575), .E(N522), .C(inClock), .Q(\FIFO[5][2] ) );
  DFE1 \FIFO_reg[5][1]  ( .D(n559), .E(N522), .C(inClock), .Q(\FIFO[5][1] ) );
  DFE1 \FIFO_reg[5][0]  ( .D(n543), .E(N522), .C(inClock), .Q(\FIFO[5][0] ) );
  DFE1 \FIFO_reg[4][3]  ( .D(n591), .E(N524), .C(inClock), .Q(\FIFO[4][3] ) );
  DFE1 \FIFO_reg[4][2]  ( .D(n575), .E(N524), .C(inClock), .Q(\FIFO[4][2] ) );
  DFE1 \FIFO_reg[4][1]  ( .D(n559), .E(N524), .C(inClock), .Q(\FIFO[4][1] ) );
  DFE1 \FIFO_reg[4][0]  ( .D(n543), .E(N524), .C(inClock), .Q(\FIFO[4][0] ) );
  DFE1 \FIFO_reg[3][3]  ( .D(n591), .E(N525), .C(inClock), .Q(\FIFO[3][3] ) );
  DFE1 \FIFO_reg[3][2]  ( .D(n575), .E(N525), .C(inClock), .Q(\FIFO[3][2] ) );
  DFE1 \FIFO_reg[3][1]  ( .D(n559), .E(N525), .C(inClock), .Q(\FIFO[3][1] ) );
  DFE1 \FIFO_reg[3][0]  ( .D(n543), .E(N525), .C(inClock), .Q(\FIFO[3][0] ) );
  DFE1 \FIFO_reg[1][3]  ( .D(n591), .E(N527), .C(inClock), .Q(\FIFO[1][3] ) );
  DFE1 \FIFO_reg[1][2]  ( .D(n575), .E(N527), .C(inClock), .Q(\FIFO[1][2] ) );
  DFE1 \FIFO_reg[1][1]  ( .D(n559), .E(N527), .C(inClock), .Q(\FIFO[1][1] ) );
  DFE1 \FIFO_reg[1][0]  ( .D(n543), .E(N527), .C(inClock), .Q(\FIFO[1][0] ) );
  DFE1 \FIFO_reg[0][3]  ( .D(n591), .E(N528), .C(inClock), .Q(\FIFO[0][3] ) );
  DFE1 \FIFO_reg[0][2]  ( .D(n575), .E(N528), .C(inClock), .Q(\FIFO[0][2] ) );
  DFE1 \FIFO_reg[0][1]  ( .D(n559), .E(N528), .C(inClock), .Q(\FIFO[0][1] ) );
  DFE1 \FIFO_reg[0][0]  ( .D(n543), .E(N528), .C(inClock), .Q(\FIFO[0][0] ) );
  DFE1 \i_FIFO_reg[4]  ( .D(n645), .E(N396), .C(inClock), .Q(N41) );
  DFE1 \i_FIFO_reg[5]  ( .D(n646), .E(N396), .C(inClock), .Q(N42) );
  DFE1 \i_FIFO_reg[3]  ( .D(n644), .E(N396), .C(inClock), .Q(N40) );
  DFE1 \j_FIFO_reg[2]  ( .D(N227), .E(n600), .C(inClock), .Q(j_FIFO[2]), .QN(
        n491) );
  DFE1 \j_FIFO_reg[3]  ( .D(N228), .E(n600), .C(inClock), .Q(j_FIFO[3]), .QN(
        n512) );
  DFE1 \sigWRCOUNT_reg[7]  ( .D(n629), .E(N392), .C(inClock), .Q(
        outWriteCount[7]), .QN(n504) );
  DFE1 \sigWRCOUNT_reg[6]  ( .D(n628), .E(N392), .C(inClock), .Q(
        outWriteCount[6]), .QN(n506) );
  DFE1 \j_FIFO_reg[4]  ( .D(N229), .E(n600), .C(inClock), .Q(j_FIFO[4]), .QN(
        n486) );
  DFE1 \j_FIFO_reg[5]  ( .D(N230), .E(n600), .C(inClock), .Q(j_FIFO[5]), .QN(
        n488) );
  DFE1 \i_FIFO_reg[6]  ( .D(n647), .E(N396), .C(inClock), .Q(N43) );
  DFE1 \j_FIFO_reg[6]  ( .D(N231), .E(n600), .C(inClock), .Q(j_FIFO[6]), .QN(
        n485) );
  DFE1 \i_FIFO_reg[1]  ( .D(n642), .E(N396), .C(inClock), .Q(N38) );
  DFE1 \i_FIFO_reg[2]  ( .D(n643), .E(N396), .C(inClock), .Q(n487), .QN(n503)
         );
  DFE1 \sigRDCOUNT_reg[4]  ( .D(n634), .E(N393), .C(inClock), .Q(
        outReadCount[4]), .QN(n496) );
  DFE1 \sigRDCOUNT_reg[5]  ( .D(n635), .E(N393), .C(inClock), .Q(
        outReadCount[5]), .QN(n497) );
  DFE1 \sigRDCOUNT_reg[6]  ( .D(n636), .E(N393), .C(inClock), .Q(
        outReadCount[6]), .QN(n501) );
  DFE1 \j_FIFO_reg[1]  ( .D(N226), .E(n600), .C(inClock), .Q(j_FIFO[1]), .QN(
        n511) );
  DFE1 \sigWRCOUNT_reg[5]  ( .D(n627), .E(N392), .C(inClock), .Q(
        outWriteCount[5]), .QN(n508) );
  DFE1 \j_FIFO_reg[0]  ( .D(N225), .E(n600), .C(inClock), .Q(j_FIFO[0]), .QN(
        n490) );
  DFE1 \sigWRCOUNT_reg[4]  ( .D(n626), .E(N392), .C(inClock), .Q(
        outWriteCount[4]), .QN(n509) );
  DFE1 \sigRDCOUNT_reg[1]  ( .D(n631), .E(N393), .C(inClock), .Q(
        outReadCount[1]), .QN(n493) );
  DFE1 \sigRDCOUNT_reg[2]  ( .D(n632), .E(N393), .C(inClock), .Q(
        outReadCount[2]), .QN(n495) );
  DFE1 \sigRDCOUNT_reg[3]  ( .D(n633), .E(N393), .C(inClock), .Q(
        outReadCount[3]), .QN(n498) );
  DFE1 \sigWRCOUNT_reg[2]  ( .D(n624), .E(N392), .C(inClock), .Q(
        outWriteCount[2]), .QN(n500) );
  DFE1 \sigWRCOUNT_reg[3]  ( .D(n625), .E(N392), .C(inClock), .Q(
        outWriteCount[3]), .QN(n507) );
  DFE1 \sigWRCOUNT_reg[1]  ( .D(n623), .E(N392), .C(inClock), .Q(
        outWriteCount[1]) );
  DFE1 \sigRDCOUNT_reg[0]  ( .D(n630), .E(N393), .C(inClock), .Q(
        outReadCount[0]), .QN(n494) );
  DFE1 \sigWRCOUNT_reg[0]  ( .D(n622), .E(N392), .C(inClock), .Q(
        outWriteCount[0]), .QN(n499) );
  IMUX21 U464 ( .A(n357), .B(n358), .S(N43), .Q(N203) );
  MUX41 U628 ( .A(N203), .B(N201), .C(N202), .D(N200), .S0(N45), .S1(N44), .Q(
        N204) );
  IMUX40 U471 ( .A(n390), .B(n391), .C(n392), .D(n393), .S0(n605), .S1(n522), 
        .Q(n389) );
  IMUX40 U542 ( .A(n374), .B(n364), .C(n369), .D(n359), .S0(n520), .S1(n521), 
        .Q(n400) );
  IMUX40 U559 ( .A(n394), .B(n384), .C(n389), .D(n379), .S0(n520), .S1(n521), 
        .Q(n399) );
  IMUX21 U473 ( .A(n399), .B(n400), .S(N43), .Q(N202) );
  IMUX40 U480 ( .A(n432), .B(n433), .C(n434), .D(n435), .S0(n604), .S1(n522), 
        .Q(n431) );
  IMUX40 U576 ( .A(n416), .B(n406), .C(n411), .D(n401), .S0(n520), .S1(n521), 
        .Q(n442) );
  IMUX40 U593 ( .A(n436), .B(n426), .C(n431), .D(n421), .S0(n520), .S1(n521), 
        .Q(n441) );
  IMUX21 U482 ( .A(n441), .B(n442), .S(N43), .Q(N201) );
  IMUX40 U498 ( .A(\FIFO[100][0] ), .B(\FIFO[101][0] ), .C(\FIFO[102][0] ), 
        .D(\FIFO[103][0] ), .S0(n620), .S1(n606), .Q(n325) );
  IMUX40 U494 ( .A(\FIFO[116][0] ), .B(\FIFO[117][0] ), .C(\FIFO[118][0] ), 
        .D(\FIFO[119][0] ), .S0(n620), .S1(n606), .Q(n320) );
  IMUX40 U519 ( .A(\FIFO[20][0] ), .B(\FIFO[21][0] ), .C(\FIFO[22][0] ), .D(
        \FIFO[23][0] ), .S0(n616), .S1(n523), .Q(n350) );
  IMUX40 U515 ( .A(\FIFO[36][0] ), .B(\FIFO[37][0] ), .C(\FIFO[38][0] ), .D(
        \FIFO[39][0] ), .S0(n616), .S1(N38), .Q(n345) );
  IMUX40 U523 ( .A(\FIFO[4][0] ), .B(\FIFO[5][0] ), .C(\FIFO[6][0] ), .D(
        \FIFO[7][0] ), .S0(n614), .S1(n610), .Q(n355) );
  IMUX40 U502 ( .A(\FIFO[84][0] ), .B(\FIFO[85][0] ), .C(\FIFO[86][0] ), .D(
        \FIFO[87][0] ), .S0(n619), .S1(N38), .Q(n330) );
  IMUX40 U553 ( .A(\FIFO[20][1] ), .B(\FIFO[21][1] ), .C(\FIFO[22][1] ), .D(
        \FIFO[23][1] ), .S0(n616), .S1(n606), .Q(n392) );
  IMUX40 U587 ( .A(\FIFO[20][2] ), .B(\FIFO[21][2] ), .C(\FIFO[22][2] ), .D(
        \FIFO[23][2] ), .S0(n614), .S1(n607), .Q(n434) );
  IMUX40 U621 ( .A(\FIFO[20][3] ), .B(\FIFO[21][3] ), .C(\FIFO[22][3] ), .D(
        \FIFO[23][3] ), .S0(n611), .S1(n609), .Q(n476) );
  IMUX40 U535 ( .A(\FIFO[88][1] ), .B(\FIFO[89][1] ), .C(\FIFO[90][1] ), .D(
        \FIFO[91][1] ), .S0(n618), .S1(n606), .Q(n371) );
  IMUX40 U534 ( .A(\FIFO[92][1] ), .B(\FIFO[93][1] ), .C(\FIFO[94][1] ), .D(
        \FIFO[95][1] ), .S0(n618), .S1(n606), .Q(n373) );
  IMUX40 U536 ( .A(\FIFO[84][1] ), .B(\FIFO[85][1] ), .C(\FIFO[86][1] ), .D(
        \FIFO[87][1] ), .S0(n618), .S1(n606), .Q(n372) );
  IMUX40 U467 ( .A(n370), .B(n371), .C(n372), .D(n373), .S0(n605), .S1(n522), 
        .Q(n369) );
  IMUX40 U569 ( .A(\FIFO[88][2] ), .B(\FIFO[89][2] ), .C(\FIFO[90][2] ), .D(
        \FIFO[91][2] ), .S0(n615), .S1(N38), .Q(n413) );
  IMUX40 U568 ( .A(\FIFO[92][2] ), .B(\FIFO[93][2] ), .C(\FIFO[94][2] ), .D(
        \FIFO[95][2] ), .S0(n615), .S1(n608), .Q(n415) );
  IMUX40 U570 ( .A(\FIFO[84][2] ), .B(\FIFO[85][2] ), .C(\FIFO[86][2] ), .D(
        \FIFO[87][2] ), .S0(n615), .S1(n523), .Q(n414) );
  IMUX40 U476 ( .A(n412), .B(n413), .C(n414), .D(n415), .S0(N40), .S1(n522), 
        .Q(n411) );
  IMUX40 U603 ( .A(\FIFO[88][3] ), .B(\FIFO[89][3] ), .C(\FIFO[90][3] ), .D(
        \FIFO[91][3] ), .S0(n612), .S1(n608), .Q(n455) );
  IMUX40 U602 ( .A(\FIFO[92][3] ), .B(\FIFO[93][3] ), .C(\FIFO[94][3] ), .D(
        \FIFO[95][3] ), .S0(n612), .S1(n608), .Q(n457) );
  IMUX40 U604 ( .A(\FIFO[84][3] ), .B(\FIFO[85][3] ), .C(\FIFO[86][3] ), .D(
        \FIFO[87][3] ), .S0(n612), .S1(n608), .Q(n456) );
  IMUX40 U485 ( .A(n454), .B(n455), .C(n456), .D(n457), .S0(n604), .S1(n522), 
        .Q(n453) );
  IMUX40 U496 ( .A(\FIFO[108][0] ), .B(\FIFO[109][0] ), .C(\FIFO[110][0] ), 
        .D(\FIFO[111][0] ), .S0(n620), .S1(n606), .Q(n326) );
  IMUX40 U497 ( .A(\FIFO[104][0] ), .B(\FIFO[105][0] ), .C(\FIFO[106][0] ), 
        .D(\FIFO[107][0] ), .S0(n620), .S1(n607), .Q(n324) );
  IMUX40 U499 ( .A(\FIFO[96][0] ), .B(\FIFO[97][0] ), .C(\FIFO[98][0] ), .D(
        \FIFO[99][0] ), .S0(n620), .S1(N38), .Q(n323) );
  IMUX40 U492 ( .A(\FIFO[124][0] ), .B(\FIFO[125][0] ), .C(\FIFO[126][0] ), 
        .D(\FIFO[127][0] ), .S0(n620), .S1(n609), .Q(n321) );
  IMUX40 U493 ( .A(\FIFO[120][0] ), .B(\FIFO[121][0] ), .C(\FIFO[122][0] ), 
        .D(\FIFO[123][0] ), .S0(n620), .S1(N38), .Q(n319) );
  IMUX40 U495 ( .A(\FIFO[112][0] ), .B(\FIFO[113][0] ), .C(\FIFO[114][0] ), 
        .D(\FIFO[115][0] ), .S0(n620), .S1(N38), .Q(n318) );
  IMUX40 U517 ( .A(\FIFO[28][0] ), .B(\FIFO[29][0] ), .C(\FIFO[30][0] ), .D(
        \FIFO[31][0] ), .S0(n615), .S1(N38), .Q(n351) );
  IMUX40 U518 ( .A(\FIFO[24][0] ), .B(\FIFO[25][0] ), .C(\FIFO[26][0] ), .D(
        \FIFO[27][0] ), .S0(n615), .S1(n523), .Q(n349) );
  IMUX40 U520 ( .A(\FIFO[16][0] ), .B(\FIFO[17][0] ), .C(\FIFO[18][0] ), .D(
        \FIFO[19][0] ), .S0(n617), .S1(n606), .Q(n348) );
  IMUX40 U513 ( .A(\FIFO[44][0] ), .B(\FIFO[45][0] ), .C(\FIFO[46][0] ), .D(
        \FIFO[47][0] ), .S0(n614), .S1(n610), .Q(n346) );
  IMUX40 U514 ( .A(\FIFO[40][0] ), .B(\FIFO[41][0] ), .C(\FIFO[42][0] ), .D(
        \FIFO[43][0] ), .S0(n613), .S1(n523), .Q(n344) );
  IMUX40 U516 ( .A(\FIFO[32][0] ), .B(\FIFO[33][0] ), .C(\FIFO[34][0] ), .D(
        \FIFO[35][0] ), .S0(n613), .S1(n523), .Q(n343) );
  IMUX40 U521 ( .A(\FIFO[12][0] ), .B(\FIFO[13][0] ), .C(\FIFO[14][0] ), .D(
        \FIFO[15][0] ), .S0(n617), .S1(n610), .Q(n356) );
  IMUX40 U522 ( .A(\FIFO[8][0] ), .B(\FIFO[9][0] ), .C(\FIFO[10][0] ), .D(
        \FIFO[11][0] ), .S0(n617), .S1(n607), .Q(n354) );
  IMUX40 U524 ( .A(\FIFO[0][0] ), .B(\FIFO[1][0] ), .C(\FIFO[2][0] ), .D(
        \FIFO[3][0] ), .S0(n614), .S1(n609), .Q(n353) );
  IMUX40 U512 ( .A(\FIFO[48][0] ), .B(\FIFO[49][0] ), .C(\FIFO[50][0] ), .D(
        \FIFO[51][0] ), .S0(n619), .S1(n523), .Q(n338) );
  IMUX40 U500 ( .A(\FIFO[92][0] ), .B(\FIFO[93][0] ), .C(\FIFO[94][0] ), .D(
        \FIFO[95][0] ), .S0(n619), .S1(n609), .Q(n331) );
  IMUX40 U501 ( .A(\FIFO[88][0] ), .B(\FIFO[89][0] ), .C(\FIFO[90][0] ), .D(
        \FIFO[91][0] ), .S0(n619), .S1(N38), .Q(n329) );
  IMUX40 U503 ( .A(\FIFO[80][0] ), .B(\FIFO[81][0] ), .C(\FIFO[82][0] ), .D(
        \FIFO[83][0] ), .S0(n619), .S1(N38), .Q(n328) );
  IMUX40 U507 ( .A(\FIFO[64][0] ), .B(\FIFO[65][0] ), .C(\FIFO[66][0] ), .D(
        \FIFO[67][0] ), .S0(n619), .S1(n523), .Q(n333) );
  IMUX40 U551 ( .A(\FIFO[28][1] ), .B(\FIFO[29][1] ), .C(\FIFO[30][1] ), .D(
        \FIFO[31][1] ), .S0(n616), .S1(n608), .Q(n393) );
  IMUX40 U552 ( .A(\FIFO[24][1] ), .B(\FIFO[25][1] ), .C(\FIFO[26][1] ), .D(
        \FIFO[27][1] ), .S0(n616), .S1(N38), .Q(n391) );
  IMUX40 U554 ( .A(\FIFO[16][1] ), .B(\FIFO[17][1] ), .C(\FIFO[18][1] ), .D(
        \FIFO[19][1] ), .S0(n616), .S1(n607), .Q(n390) );
  IMUX40 U550 ( .A(\FIFO[32][1] ), .B(\FIFO[33][1] ), .C(\FIFO[34][1] ), .D(
        \FIFO[35][1] ), .S0(n617), .S1(n610), .Q(n385) );
  IMUX40 U558 ( .A(\FIFO[0][1] ), .B(\FIFO[1][1] ), .C(\FIFO[2][1] ), .D(
        \FIFO[3][1] ), .S0(n616), .S1(n608), .Q(n395) );
  IMUX40 U546 ( .A(\FIFO[48][1] ), .B(\FIFO[49][1] ), .C(\FIFO[50][1] ), .D(
        \FIFO[51][1] ), .S0(n617), .S1(n606), .Q(n380) );
  IMUX40 U537 ( .A(\FIFO[80][1] ), .B(\FIFO[81][1] ), .C(\FIFO[82][1] ), .D(
        \FIFO[83][1] ), .S0(n618), .S1(n606), .Q(n370) );
  IMUX40 U533 ( .A(\FIFO[96][1] ), .B(\FIFO[97][1] ), .C(\FIFO[98][1] ), .D(
        \FIFO[99][1] ), .S0(n618), .S1(n610), .Q(n365) );
  IMUX40 U541 ( .A(\FIFO[64][1] ), .B(\FIFO[65][1] ), .C(\FIFO[66][1] ), .D(
        \FIFO[67][1] ), .S0(n617), .S1(n606), .Q(n375) );
  IMUX40 U529 ( .A(\FIFO[112][1] ), .B(\FIFO[113][1] ), .C(\FIFO[114][1] ), 
        .D(\FIFO[115][1] ), .S0(n618), .S1(n610), .Q(n360) );
  IMUX40 U585 ( .A(\FIFO[28][2] ), .B(\FIFO[29][2] ), .C(\FIFO[30][2] ), .D(
        \FIFO[31][2] ), .S0(n614), .S1(n607), .Q(n435) );
  IMUX40 U586 ( .A(\FIFO[24][2] ), .B(\FIFO[25][2] ), .C(\FIFO[26][2] ), .D(
        \FIFO[27][2] ), .S0(n614), .S1(n607), .Q(n433) );
  IMUX40 U588 ( .A(\FIFO[16][2] ), .B(\FIFO[17][2] ), .C(\FIFO[18][2] ), .D(
        \FIFO[19][2] ), .S0(n614), .S1(n607), .Q(n432) );
  IMUX40 U584 ( .A(\FIFO[32][2] ), .B(\FIFO[33][2] ), .C(\FIFO[34][2] ), .D(
        \FIFO[35][2] ), .S0(n614), .S1(n607), .Q(n427) );
  IMUX40 U592 ( .A(\FIFO[0][2] ), .B(\FIFO[1][2] ), .C(\FIFO[2][2] ), .D(
        \FIFO[3][2] ), .S0(n613), .S1(n607), .Q(n437) );
  IMUX40 U580 ( .A(\FIFO[48][2] ), .B(\FIFO[49][2] ), .C(\FIFO[50][2] ), .D(
        \FIFO[51][2] ), .S0(n614), .S1(n607), .Q(n422) );
  IMUX40 U571 ( .A(\FIFO[80][2] ), .B(\FIFO[81][2] ), .C(\FIFO[82][2] ), .D(
        \FIFO[83][2] ), .S0(n615), .S1(N38), .Q(n412) );
  IMUX40 U567 ( .A(\FIFO[96][2] ), .B(\FIFO[97][2] ), .C(\FIFO[98][2] ), .D(
        \FIFO[99][2] ), .S0(n615), .S1(N38), .Q(n407) );
  IMUX40 U575 ( .A(\FIFO[64][2] ), .B(\FIFO[65][2] ), .C(\FIFO[66][2] ), .D(
        \FIFO[67][2] ), .S0(n615), .S1(N38), .Q(n417) );
  IMUX40 U563 ( .A(\FIFO[112][2] ), .B(\FIFO[113][2] ), .C(\FIFO[114][2] ), 
        .D(\FIFO[115][2] ), .S0(n616), .S1(n607), .Q(n402) );
  IMUX40 U619 ( .A(\FIFO[28][3] ), .B(\FIFO[29][3] ), .C(\FIFO[30][3] ), .D(
        \FIFO[31][3] ), .S0(n611), .S1(n609), .Q(n477) );
  IMUX40 U620 ( .A(\FIFO[24][3] ), .B(\FIFO[25][3] ), .C(\FIFO[26][3] ), .D(
        \FIFO[27][3] ), .S0(n611), .S1(n609), .Q(n475) );
  IMUX40 U622 ( .A(\FIFO[16][3] ), .B(\FIFO[17][3] ), .C(\FIFO[18][3] ), .D(
        \FIFO[19][3] ), .S0(n611), .S1(n609), .Q(n474) );
  IMUX40 U626 ( .A(\FIFO[0][3] ), .B(\FIFO[1][3] ), .C(\FIFO[2][3] ), .D(
        \FIFO[3][3] ), .S0(n611), .S1(n610), .Q(n479) );
  IMUX40 U618 ( .A(\FIFO[32][3] ), .B(\FIFO[33][3] ), .C(\FIFO[34][3] ), .D(
        \FIFO[35][3] ), .S0(n611), .S1(n609), .Q(n469) );
  IMUX40 U614 ( .A(\FIFO[48][3] ), .B(\FIFO[49][3] ), .C(\FIFO[50][3] ), .D(
        \FIFO[51][3] ), .S0(n612), .S1(n609), .Q(n464) );
  IMUX40 U605 ( .A(\FIFO[80][3] ), .B(\FIFO[81][3] ), .C(\FIFO[82][3] ), .D(
        \FIFO[83][3] ), .S0(n612), .S1(n608), .Q(n454) );
  IMUX40 U609 ( .A(\FIFO[64][3] ), .B(\FIFO[65][3] ), .C(\FIFO[66][3] ), .D(
        \FIFO[67][3] ), .S0(n612), .S1(n609), .Q(n459) );
  IMUX40 U601 ( .A(\FIFO[96][3] ), .B(\FIFO[97][3] ), .C(\FIFO[98][3] ), .D(
        \FIFO[99][3] ), .S0(n613), .S1(n608), .Q(n449) );
  IMUX40 U597 ( .A(\FIFO[112][3] ), .B(\FIFO[113][3] ), .C(\FIFO[114][3] ), 
        .D(\FIFO[115][3] ), .S0(n613), .S1(n608), .Q(n444) );
  IMUX40 U624 ( .A(\FIFO[8][3] ), .B(\FIFO[9][3] ), .C(\FIFO[10][3] ), .D(
        \FIFO[11][3] ), .S0(n611), .S1(n610), .Q(n480) );
  IMUX40 U623 ( .A(\FIFO[12][3] ), .B(\FIFO[13][3] ), .C(\FIFO[14][3] ), .D(
        \FIFO[15][3] ), .S0(n611), .S1(n610), .Q(n482) );
  IMUX40 U625 ( .A(\FIFO[4][3] ), .B(\FIFO[5][3] ), .C(\FIFO[6][3] ), .D(
        \FIFO[7][3] ), .S0(n611), .S1(n610), .Q(n481) );
  IMUX40 U490 ( .A(n479), .B(n480), .C(n481), .D(n482), .S0(n604), .S1(n522), 
        .Q(n478) );
  IMUX40 U510 ( .A(\FIFO[56][0] ), .B(\FIFO[57][0] ), .C(\FIFO[58][0] ), .D(
        \FIFO[59][0] ), .S0(n619), .S1(n523), .Q(n339) );
  IMUX40 U509 ( .A(\FIFO[60][0] ), .B(\FIFO[61][0] ), .C(\FIFO[62][0] ), .D(
        \FIFO[63][0] ), .S0(n619), .S1(n608), .Q(n341) );
  IMUX40 U511 ( .A(\FIFO[52][0] ), .B(\FIFO[53][0] ), .C(\FIFO[54][0] ), .D(
        \FIFO[55][0] ), .S0(n619), .S1(n523), .Q(n340) );
  IMUX40 U460 ( .A(n338), .B(n339), .C(n340), .D(n341), .S0(n605), .S1(n487), 
        .Q(n337) );
  IMUX40 U505 ( .A(\FIFO[72][0] ), .B(\FIFO[73][0] ), .C(\FIFO[74][0] ), .D(
        \FIFO[75][0] ), .S0(n619), .S1(N38), .Q(n334) );
  IMUX40 U504 ( .A(\FIFO[76][0] ), .B(\FIFO[77][0] ), .C(\FIFO[78][0] ), .D(
        \FIFO[79][0] ), .S0(n619), .S1(n609), .Q(n336) );
  IMUX40 U506 ( .A(\FIFO[68][0] ), .B(\FIFO[69][0] ), .C(\FIFO[70][0] ), .D(
        \FIFO[71][0] ), .S0(n619), .S1(n523), .Q(n335) );
  IMUX40 U459 ( .A(n333), .B(n334), .C(n335), .D(n336), .S0(n605), .S1(n522), 
        .Q(n332) );
  IMUX40 U548 ( .A(\FIFO[40][1] ), .B(\FIFO[41][1] ), .C(\FIFO[42][1] ), .D(
        \FIFO[43][1] ), .S0(n617), .S1(n606), .Q(n386) );
  IMUX40 U547 ( .A(\FIFO[44][1] ), .B(\FIFO[45][1] ), .C(\FIFO[46][1] ), .D(
        \FIFO[47][1] ), .S0(n617), .S1(n606), .Q(n388) );
  IMUX40 U549 ( .A(\FIFO[36][1] ), .B(\FIFO[37][1] ), .C(\FIFO[38][1] ), .D(
        \FIFO[39][1] ), .S0(n617), .S1(n610), .Q(n387) );
  IMUX40 U470 ( .A(n385), .B(n386), .C(n387), .D(n388), .S0(n604), .S1(n487), 
        .Q(n384) );
  IMUX40 U556 ( .A(\FIFO[8][1] ), .B(\FIFO[9][1] ), .C(\FIFO[10][1] ), .D(
        \FIFO[11][1] ), .S0(n616), .S1(n609), .Q(n396) );
  IMUX40 U555 ( .A(\FIFO[12][1] ), .B(\FIFO[13][1] ), .C(\FIFO[14][1] ), .D(
        \FIFO[15][1] ), .S0(n616), .S1(N38), .Q(n398) );
  IMUX40 U557 ( .A(\FIFO[4][1] ), .B(\FIFO[5][1] ), .C(\FIFO[6][1] ), .D(
        \FIFO[7][1] ), .S0(n616), .S1(n523), .Q(n397) );
  IMUX40 U472 ( .A(n395), .B(n396), .C(n397), .D(n398), .S0(N40), .S1(n522), 
        .Q(n394) );
  IMUX40 U544 ( .A(\FIFO[56][1] ), .B(\FIFO[57][1] ), .C(\FIFO[58][1] ), .D(
        \FIFO[59][1] ), .S0(n617), .S1(n606), .Q(n381) );
  IMUX40 U543 ( .A(\FIFO[60][1] ), .B(\FIFO[61][1] ), .C(\FIFO[62][1] ), .D(
        \FIFO[63][1] ), .S0(n617), .S1(n606), .Q(n383) );
  IMUX40 U545 ( .A(\FIFO[52][1] ), .B(\FIFO[53][1] ), .C(\FIFO[54][1] ), .D(
        \FIFO[55][1] ), .S0(n617), .S1(n606), .Q(n382) );
  IMUX40 U469 ( .A(n380), .B(n381), .C(n382), .D(n383), .S0(n605), .S1(n487), 
        .Q(n379) );
  IMUX40 U531 ( .A(\FIFO[104][1] ), .B(\FIFO[105][1] ), .C(\FIFO[106][1] ), 
        .D(\FIFO[107][1] ), .S0(n618), .S1(n610), .Q(n366) );
  IMUX40 U530 ( .A(\FIFO[108][1] ), .B(\FIFO[109][1] ), .C(\FIFO[110][1] ), 
        .D(\FIFO[111][1] ), .S0(n618), .S1(n610), .Q(n368) );
  IMUX40 U532 ( .A(\FIFO[100][1] ), .B(\FIFO[101][1] ), .C(\FIFO[102][1] ), 
        .D(\FIFO[103][1] ), .S0(n618), .S1(n610), .Q(n367) );
  IMUX40 U466 ( .A(n365), .B(n366), .C(n367), .D(n368), .S0(n604), .S1(n487), 
        .Q(n364) );
  IMUX40 U539 ( .A(\FIFO[72][1] ), .B(\FIFO[73][1] ), .C(\FIFO[74][1] ), .D(
        \FIFO[75][1] ), .S0(n617), .S1(n606), .Q(n376) );
  IMUX40 U538 ( .A(\FIFO[76][1] ), .B(\FIFO[77][1] ), .C(\FIFO[78][1] ), .D(
        \FIFO[79][1] ), .S0(n617), .S1(n606), .Q(n378) );
  IMUX40 U540 ( .A(\FIFO[68][1] ), .B(\FIFO[69][1] ), .C(\FIFO[70][1] ), .D(
        \FIFO[71][1] ), .S0(n617), .S1(n606), .Q(n377) );
  IMUX40 U468 ( .A(n375), .B(n376), .C(n377), .D(n378), .S0(N40), .S1(n522), 
        .Q(n374) );
  IMUX40 U527 ( .A(\FIFO[120][1] ), .B(\FIFO[121][1] ), .C(\FIFO[122][1] ), 
        .D(\FIFO[123][1] ), .S0(n618), .S1(n610), .Q(n361) );
  IMUX40 U526 ( .A(\FIFO[124][1] ), .B(\FIFO[125][1] ), .C(\FIFO[126][1] ), 
        .D(\FIFO[127][1] ), .S0(n618), .S1(n610), .Q(n363) );
  IMUX40 U528 ( .A(\FIFO[116][1] ), .B(\FIFO[117][1] ), .C(\FIFO[118][1] ), 
        .D(\FIFO[119][1] ), .S0(n618), .S1(n610), .Q(n362) );
  IMUX40 U465 ( .A(n360), .B(n361), .C(n362), .D(n363), .S0(n605), .S1(n487), 
        .Q(n359) );
  IMUX40 U582 ( .A(\FIFO[40][2] ), .B(\FIFO[41][2] ), .C(\FIFO[42][2] ), .D(
        \FIFO[43][2] ), .S0(n614), .S1(n607), .Q(n428) );
  IMUX40 U581 ( .A(\FIFO[44][2] ), .B(\FIFO[45][2] ), .C(\FIFO[46][2] ), .D(
        \FIFO[47][2] ), .S0(n614), .S1(n607), .Q(n430) );
  IMUX40 U583 ( .A(\FIFO[36][2] ), .B(\FIFO[37][2] ), .C(\FIFO[38][2] ), .D(
        \FIFO[39][2] ), .S0(n614), .S1(n607), .Q(n429) );
  IMUX40 U479 ( .A(n427), .B(n428), .C(n429), .D(n430), .S0(n604), .S1(n522), 
        .Q(n426) );
  IMUX40 U590 ( .A(\FIFO[8][2] ), .B(\FIFO[9][2] ), .C(\FIFO[10][2] ), .D(
        \FIFO[11][2] ), .S0(n613), .S1(n607), .Q(n438) );
  IMUX40 U589 ( .A(\FIFO[12][2] ), .B(\FIFO[13][2] ), .C(\FIFO[14][2] ), .D(
        \FIFO[15][2] ), .S0(n613), .S1(n607), .Q(n440) );
  IMUX40 U591 ( .A(\FIFO[4][2] ), .B(\FIFO[5][2] ), .C(\FIFO[6][2] ), .D(
        \FIFO[7][2] ), .S0(n613), .S1(n607), .Q(n439) );
  IMUX40 U481 ( .A(n437), .B(n438), .C(n439), .D(n440), .S0(n604), .S1(n522), 
        .Q(n436) );
  IMUX40 U578 ( .A(\FIFO[56][2] ), .B(\FIFO[57][2] ), .C(\FIFO[58][2] ), .D(
        \FIFO[59][2] ), .S0(n614), .S1(N38), .Q(n423) );
  IMUX40 U577 ( .A(\FIFO[60][2] ), .B(\FIFO[61][2] ), .C(\FIFO[62][2] ), .D(
        \FIFO[63][2] ), .S0(n614), .S1(n606), .Q(n425) );
  IMUX40 U579 ( .A(\FIFO[52][2] ), .B(\FIFO[53][2] ), .C(\FIFO[54][2] ), .D(
        \FIFO[55][2] ), .S0(n614), .S1(n607), .Q(n424) );
  IMUX40 U478 ( .A(n422), .B(n423), .C(n424), .D(n425), .S0(n604), .S1(n487), 
        .Q(n421) );
  IMUX40 U565 ( .A(\FIFO[104][2] ), .B(\FIFO[105][2] ), .C(\FIFO[106][2] ), 
        .D(\FIFO[107][2] ), .S0(n615), .S1(n610), .Q(n408) );
  IMUX40 U564 ( .A(\FIFO[108][2] ), .B(\FIFO[109][2] ), .C(\FIFO[110][2] ), 
        .D(\FIFO[111][2] ), .S0(n615), .S1(n607), .Q(n410) );
  IMUX40 U566 ( .A(\FIFO[100][2] ), .B(\FIFO[101][2] ), .C(\FIFO[102][2] ), 
        .D(\FIFO[103][2] ), .S0(n615), .S1(n607), .Q(n409) );
  IMUX40 U475 ( .A(n407), .B(n408), .C(n409), .D(n410), .S0(N40), .S1(n522), 
        .Q(n406) );
  IMUX40 U573 ( .A(\FIFO[72][2] ), .B(\FIFO[73][2] ), .C(\FIFO[74][2] ), .D(
        \FIFO[75][2] ), .S0(n615), .S1(n523), .Q(n418) );
  IMUX40 U572 ( .A(\FIFO[76][2] ), .B(\FIFO[77][2] ), .C(\FIFO[78][2] ), .D(
        \FIFO[79][2] ), .S0(n615), .S1(n608), .Q(n420) );
  IMUX40 U574 ( .A(\FIFO[68][2] ), .B(\FIFO[69][2] ), .C(\FIFO[70][2] ), .D(
        \FIFO[71][2] ), .S0(n615), .S1(n609), .Q(n419) );
  IMUX40 U477 ( .A(n417), .B(n418), .C(n419), .D(n420), .S0(N40), .S1(n522), 
        .Q(n416) );
  IMUX40 U561 ( .A(\FIFO[120][2] ), .B(\FIFO[121][2] ), .C(\FIFO[122][2] ), 
        .D(\FIFO[123][2] ), .S0(n616), .S1(n608), .Q(n403) );
  IMUX40 U560 ( .A(\FIFO[124][2] ), .B(\FIFO[125][2] ), .C(\FIFO[126][2] ), 
        .D(\FIFO[127][2] ), .S0(n616), .S1(n610), .Q(n405) );
  IMUX40 U562 ( .A(\FIFO[116][2] ), .B(\FIFO[117][2] ), .C(\FIFO[118][2] ), 
        .D(\FIFO[119][2] ), .S0(n616), .S1(n610), .Q(n404) );
  IMUX40 U474 ( .A(n402), .B(n403), .C(n404), .D(n405), .S0(n605), .S1(n487), 
        .Q(n401) );
  IMUX40 U616 ( .A(\FIFO[40][3] ), .B(\FIFO[41][3] ), .C(\FIFO[42][3] ), .D(
        \FIFO[43][3] ), .S0(n611), .S1(n609), .Q(n470) );
  IMUX40 U615 ( .A(\FIFO[44][3] ), .B(\FIFO[45][3] ), .C(\FIFO[46][3] ), .D(
        \FIFO[47][3] ), .S0(n611), .S1(n609), .Q(n472) );
  IMUX40 U617 ( .A(\FIFO[36][3] ), .B(\FIFO[37][3] ), .C(\FIFO[38][3] ), .D(
        \FIFO[39][3] ), .S0(n611), .S1(n609), .Q(n471) );
  IMUX40 U488 ( .A(n469), .B(n470), .C(n471), .D(n472), .S0(n604), .S1(n487), 
        .Q(n468) );
  IMUX40 U612 ( .A(\FIFO[56][3] ), .B(\FIFO[57][3] ), .C(\FIFO[58][3] ), .D(
        \FIFO[59][3] ), .S0(n612), .S1(n609), .Q(n465) );
  IMUX40 U611 ( .A(\FIFO[60][3] ), .B(\FIFO[61][3] ), .C(\FIFO[62][3] ), .D(
        \FIFO[63][3] ), .S0(n612), .S1(n609), .Q(n467) );
  IMUX40 U613 ( .A(\FIFO[52][3] ), .B(\FIFO[53][3] ), .C(\FIFO[54][3] ), .D(
        \FIFO[55][3] ), .S0(n612), .S1(n609), .Q(n466) );
  IMUX40 U487 ( .A(n464), .B(n465), .C(n466), .D(n467), .S0(n604), .S1(n487), 
        .Q(n463) );
  IMUX40 U607 ( .A(\FIFO[72][3] ), .B(\FIFO[73][3] ), .C(\FIFO[74][3] ), .D(
        \FIFO[75][3] ), .S0(n612), .S1(n608), .Q(n460) );
  IMUX40 U606 ( .A(\FIFO[76][3] ), .B(\FIFO[77][3] ), .C(\FIFO[78][3] ), .D(
        \FIFO[79][3] ), .S0(n612), .S1(n608), .Q(n462) );
  IMUX40 U608 ( .A(\FIFO[68][3] ), .B(\FIFO[69][3] ), .C(\FIFO[70][3] ), .D(
        \FIFO[71][3] ), .S0(n612), .S1(n609), .Q(n461) );
  IMUX40 U486 ( .A(n459), .B(n460), .C(n461), .D(n462), .S0(n604), .S1(n522), 
        .Q(n458) );
  IMUX40 U599 ( .A(\FIFO[104][3] ), .B(\FIFO[105][3] ), .C(\FIFO[106][3] ), 
        .D(\FIFO[107][3] ), .S0(n613), .S1(n608), .Q(n450) );
  IMUX40 U598 ( .A(\FIFO[108][3] ), .B(\FIFO[109][3] ), .C(\FIFO[110][3] ), 
        .D(\FIFO[111][3] ), .S0(n613), .S1(n608), .Q(n452) );
  IMUX40 U600 ( .A(\FIFO[100][3] ), .B(\FIFO[101][3] ), .C(\FIFO[102][3] ), 
        .D(\FIFO[103][3] ), .S0(n613), .S1(n608), .Q(n451) );
  IMUX40 U484 ( .A(n449), .B(n450), .C(n451), .D(n452), .S0(n604), .S1(n487), 
        .Q(n448) );
  IMUX40 U595 ( .A(\FIFO[120][3] ), .B(\FIFO[121][3] ), .C(\FIFO[122][3] ), 
        .D(\FIFO[123][3] ), .S0(n613), .S1(n608), .Q(n445) );
  IMUX40 U594 ( .A(\FIFO[124][3] ), .B(\FIFO[125][3] ), .C(\FIFO[126][3] ), 
        .D(\FIFO[127][3] ), .S0(n613), .S1(n608), .Q(n447) );
  IMUX40 U596 ( .A(\FIFO[116][3] ), .B(\FIFO[117][3] ), .C(\FIFO[118][3] ), 
        .D(\FIFO[119][3] ), .S0(n613), .S1(n608), .Q(n446) );
  IMUX40 U483 ( .A(n444), .B(n445), .C(n446), .D(n447), .S0(n604), .S1(n487), 
        .Q(n443) );
  IMUX40 U489 ( .A(n474), .B(n475), .C(n476), .D(n477), .S0(n604), .S1(n522), 
        .Q(n473) );
  IMUX40 U610 ( .A(n458), .B(n448), .C(n453), .D(n443), .S0(n520), .S1(n521), 
        .Q(n484) );
  IMUX40 U627 ( .A(n478), .B(n468), .C(n473), .D(n463), .S0(n520), .S1(n521), 
        .Q(n483) );
  IMUX21 U491 ( .A(n483), .B(n484), .S(N43), .Q(N200) );
  DFE1 sigOutData_reg ( .D(n649), .E(N199), .C(inClock), .Q(outData) );
  DFE1 sigWError_reg ( .D(N382), .E(N530), .C(inClock), .Q(outWriteError) );
  DFE1 sigRError_reg ( .D(N381), .E(N532), .C(inClock), .Q(outReadError) );
  IMUX40 U458 ( .A(n328), .B(n329), .C(n330), .D(n331), .S0(n605), .S1(n522), 
        .Q(n327) );
  IMUX40 U456 ( .A(n318), .B(n319), .C(n320), .D(n321), .S0(n605), .S1(n487), 
        .Q(n317) );
  IMUX40 U457 ( .A(n323), .B(n324), .C(n325), .D(n326), .S0(n605), .S1(n522), 
        .Q(n322) );
  IMUX40 U508 ( .A(n332), .B(n322), .C(n327), .D(n317), .S0(n520), .S1(n521), 
        .Q(n358) );
  IMUX40 U463 ( .A(n353), .B(n354), .C(n355), .D(n356), .S0(n605), .S1(n522), 
        .Q(n352) );
  IMUX40 U461 ( .A(n343), .B(n344), .C(n345), .D(n346), .S0(n605), .S1(n522), 
        .Q(n342) );
  IMUX40 U462 ( .A(n348), .B(n349), .C(n350), .D(n351), .S0(n605), .S1(n522), 
        .Q(n347) );
  IMUX40 U525 ( .A(n352), .B(n342), .C(n347), .D(n337), .S0(n520), .S1(n521), 
        .Q(n357) );
  DFE1 \i_FIFO_reg[0]  ( .D(n641), .E(N396), .C(inClock), .QN(n502) );
  NOR21 U629 ( .A(n286), .B(n516), .Q(N231) );
  NOR21 U630 ( .A(n601), .B(n99), .Q(n100) );
  INV3 U631 ( .A(n600), .Q(n593) );
  INV3 U632 ( .A(n600), .Q(n594) );
  INV3 U633 ( .A(n600), .Q(n595) );
  INV3 U634 ( .A(n600), .Q(n596) );
  INV3 U635 ( .A(n600), .Q(n597) );
  INV3 U636 ( .A(n600), .Q(n598) );
  INV3 U637 ( .A(n600), .Q(n599) );
  INV3 U638 ( .A(n600), .Q(n592) );
  INV3 U639 ( .A(n134), .Q(n665) );
  INV3 U640 ( .A(N375), .Q(n657) );
  NOR21 U641 ( .A(n280), .B(n281), .Q(N392) );
  INV3 U642 ( .A(n278), .Q(n676) );
  NAND22 U643 ( .A(n272), .B(n251), .Q(n278) );
  NAND22 U644 ( .A(n147), .B(n148), .Q(n134) );
  INV3 U645 ( .A(n100), .Q(n600) );
  INV3 U646 ( .A(n524), .Q(n525) );
  NOR40 U647 ( .A(n659), .B(n708), .C(N135), .D(N134), .Q(N375) );
  NAND22 U648 ( .A(N140), .B(n660), .Q(n708) );
  INV3 U649 ( .A(n707), .Q(n659) );
  INV3 U650 ( .A(N133), .Q(n660) );
  NOR40 U651 ( .A(N139), .B(N138), .C(N137), .D(N136), .Q(n707) );
  NOR21 U652 ( .A(n131), .B(n601), .Q(N50) );
  AOI211 U653 ( .A(n654), .B(n663), .C(n132), .Q(n131) );
  INV3 U654 ( .A(n706), .Q(n654) );
  AOI221 U655 ( .A(n134), .B(n657), .C(n663), .D(n706), .Q(n146) );
  INV3 U656 ( .A(n293), .Q(n628) );
  AOI221 U657 ( .A(N148), .B(n279), .C(N139), .D(n292), .Q(n293) );
  INV3 U658 ( .A(n502), .Q(n619) );
  INV3 U659 ( .A(n502), .Q(n615) );
  INV3 U660 ( .A(n502), .Q(n613) );
  INV3 U661 ( .A(n502), .Q(n614) );
  INV3 U662 ( .A(n502), .Q(n618) );
  INV3 U663 ( .A(n502), .Q(n617) );
  INV3 U664 ( .A(n502), .Q(n616) );
  INV3 U665 ( .A(n502), .Q(n612) );
  INV3 U666 ( .A(n502), .Q(n611) );
  INV3 U667 ( .A(n502), .Q(n620) );
  INV3 U668 ( .A(n503), .Q(n522) );
  NOR21 U669 ( .A(n286), .B(n667), .Q(N230) );
  INV3 U670 ( .A(N216), .Q(n667) );
  INV3 U671 ( .A(n295), .Q(n626) );
  AOI221 U672 ( .A(N146), .B(n279), .C(N137), .D(n292), .Q(n295) );
  INV3 U673 ( .A(n294), .Q(n627) );
  AOI221 U674 ( .A(N147), .B(n279), .C(N138), .D(n292), .Q(n294) );
  AOI211 U675 ( .A(n279), .B(n510), .C(n280), .Q(N393) );
  NOR21 U676 ( .A(n161), .B(n662), .Q(n279) );
  NOR21 U677 ( .A(n287), .B(n601), .Q(n292) );
  NOR21 U678 ( .A(n511), .B(n490), .Q(n251) );
  NAND31 U679 ( .A(n505), .B(n489), .C(n166), .Q(n148) );
  INV3 U680 ( .A(n240), .Q(n687) );
  NAND22 U681 ( .A(n241), .B(n242), .Q(n240) );
  INV3 U682 ( .A(n253), .Q(n686) );
  NAND22 U683 ( .A(n254), .B(n241), .Q(n253) );
  INV3 U684 ( .A(n244), .Q(n675) );
  NAND22 U685 ( .A(n245), .B(n242), .Q(n244) );
  INV3 U686 ( .A(n247), .Q(n683) );
  NAND22 U687 ( .A(n248), .B(n242), .Q(n247) );
  INV3 U688 ( .A(n250), .Q(n679) );
  NAND22 U689 ( .A(n251), .B(n242), .Q(n250) );
  INV3 U690 ( .A(n258), .Q(n682) );
  NAND22 U691 ( .A(n254), .B(n248), .Q(n258) );
  INV3 U692 ( .A(n262), .Q(n685) );
  NAND22 U693 ( .A(n263), .B(n241), .Q(n262) );
  INV3 U694 ( .A(n267), .Q(n681) );
  NAND22 U695 ( .A(n263), .B(n248), .Q(n267) );
  INV3 U696 ( .A(n271), .Q(n684) );
  NAND22 U697 ( .A(n272), .B(n241), .Q(n271) );
  INV3 U698 ( .A(n265), .Q(n673) );
  NAND22 U699 ( .A(n263), .B(n245), .Q(n265) );
  INV3 U700 ( .A(n274), .Q(n672) );
  NAND22 U701 ( .A(n272), .B(n245), .Q(n274) );
  INV3 U702 ( .A(n269), .Q(n677) );
  NAND22 U703 ( .A(n263), .B(n251), .Q(n269) );
  AOI211 U704 ( .A(n505), .B(n666), .C(n99), .Q(n96) );
  INV3 U705 ( .A(n276), .Q(n680) );
  NAND22 U706 ( .A(n272), .B(n248), .Q(n276) );
  INV3 U707 ( .A(n256), .Q(n674) );
  NAND22 U708 ( .A(n254), .B(n245), .Q(n256) );
  INV3 U709 ( .A(n260), .Q(n678) );
  NAND22 U710 ( .A(n254), .B(n251), .Q(n260) );
  NOR31 U711 ( .A(n99), .B(N396), .C(n662), .Q(n280) );
  NOR21 U712 ( .A(n512), .B(n491), .Q(n272) );
  NOR40 U713 ( .A(n601), .B(n162), .C(n514), .D(n492), .Q(N196) );
  NOR21 U714 ( .A(n592), .B(n103), .Q(N527) );
  AOI211 U715 ( .A(n675), .B(n527), .C(n601), .Q(n103) );
  NOR21 U716 ( .A(n592), .B(n104), .Q(N526) );
  AOI211 U717 ( .A(n683), .B(n527), .C(n601), .Q(n104) );
  NOR21 U718 ( .A(n592), .B(n105), .Q(N525) );
  AOI211 U719 ( .A(n679), .B(n527), .C(n602), .Q(n105) );
  NOR21 U720 ( .A(n592), .B(n107), .Q(N522) );
  AOI211 U721 ( .A(n674), .B(n527), .C(n602), .Q(n107) );
  NOR21 U722 ( .A(n592), .B(n108), .Q(N521) );
  AOI211 U723 ( .A(n682), .B(n527), .C(n601), .Q(n108) );
  NOR21 U724 ( .A(n592), .B(n109), .Q(N520) );
  AOI211 U725 ( .A(n678), .B(n527), .C(n602), .Q(n109) );
  NOR21 U726 ( .A(n592), .B(n110), .Q(N519) );
  AOI211 U727 ( .A(n685), .B(n527), .C(n602), .Q(n110) );
  NOR21 U728 ( .A(n592), .B(n111), .Q(N518) );
  AOI211 U729 ( .A(n673), .B(n102), .C(n602), .Q(n111) );
  NOR21 U730 ( .A(n592), .B(n112), .Q(N517) );
  AOI211 U731 ( .A(n681), .B(n527), .C(n602), .Q(n112) );
  NOR21 U732 ( .A(n592), .B(n113), .Q(N516) );
  AOI211 U733 ( .A(n677), .B(n102), .C(n602), .Q(n113) );
  NOR21 U734 ( .A(n592), .B(n114), .Q(N515) );
  AOI211 U735 ( .A(n684), .B(n527), .C(n602), .Q(n114) );
  NOR21 U736 ( .A(n592), .B(n115), .Q(N514) );
  AOI211 U737 ( .A(n672), .B(n102), .C(n602), .Q(n115) );
  NOR21 U738 ( .A(n592), .B(n277), .Q(N397) );
  AOI211 U739 ( .A(n525), .B(n676), .C(n601), .Q(n277) );
  BUF2 U740 ( .A(n523), .Q(n608) );
  BUF2 U741 ( .A(n523), .Q(n609) );
  BUF2 U742 ( .A(n523), .Q(n607) );
  BUF2 U743 ( .A(n523), .Q(n606) );
  NOR21 U744 ( .A(n596), .B(n101), .Q(N528) );
  AOI211 U745 ( .A(n527), .B(n687), .C(n603), .Q(n101) );
  NOR21 U746 ( .A(n593), .B(n116), .Q(N513) );
  AOI211 U747 ( .A(n680), .B(n527), .C(n602), .Q(n116) );
  NOR21 U748 ( .A(n593), .B(n117), .Q(N512) );
  AOI211 U749 ( .A(n676), .B(n102), .C(n602), .Q(n117) );
  NOR21 U750 ( .A(n593), .B(n118), .Q(N511) );
  AOI211 U751 ( .A(n119), .B(n687), .C(n602), .Q(n118) );
  NOR21 U752 ( .A(n593), .B(n120), .Q(N510) );
  AOI211 U753 ( .A(n119), .B(n675), .C(n602), .Q(n120) );
  NOR21 U754 ( .A(n593), .B(n121), .Q(N509) );
  AOI211 U755 ( .A(n119), .B(n683), .C(n602), .Q(n121) );
  NOR21 U756 ( .A(n593), .B(n122), .Q(N508) );
  AOI211 U757 ( .A(n119), .B(n679), .C(n602), .Q(n122) );
  NOR21 U758 ( .A(n593), .B(n123), .Q(N507) );
  AOI211 U759 ( .A(n119), .B(n686), .C(n602), .Q(n123) );
  NOR21 U760 ( .A(n593), .B(n124), .Q(N506) );
  AOI211 U761 ( .A(n119), .B(n674), .C(n602), .Q(n124) );
  NOR21 U762 ( .A(n593), .B(n125), .Q(N505) );
  AOI211 U763 ( .A(n119), .B(n682), .C(n602), .Q(n125) );
  NOR21 U764 ( .A(n593), .B(n126), .Q(N504) );
  AOI211 U765 ( .A(n119), .B(n678), .C(n603), .Q(n126) );
  NOR21 U766 ( .A(n593), .B(n127), .Q(N503) );
  AOI211 U767 ( .A(n119), .B(n685), .C(n602), .Q(n127) );
  NOR21 U768 ( .A(n593), .B(n128), .Q(N502) );
  AOI211 U769 ( .A(n119), .B(n673), .C(n603), .Q(n128) );
  NOR21 U770 ( .A(n593), .B(n129), .Q(N501) );
  AOI211 U771 ( .A(n119), .B(n681), .C(n603), .Q(n129) );
  NOR21 U772 ( .A(n594), .B(n130), .Q(N500) );
  AOI211 U773 ( .A(n119), .B(n677), .C(n603), .Q(n130) );
  NOR21 U774 ( .A(n594), .B(n135), .Q(N499) );
  AOI211 U775 ( .A(n119), .B(n684), .C(n603), .Q(n135) );
  NOR21 U776 ( .A(n594), .B(n136), .Q(N498) );
  AOI211 U777 ( .A(n119), .B(n672), .C(n603), .Q(n136) );
  NOR21 U778 ( .A(n594), .B(n137), .Q(N497) );
  AOI211 U779 ( .A(n119), .B(n680), .C(n603), .Q(n137) );
  NOR21 U780 ( .A(n594), .B(n138), .Q(N496) );
  AOI211 U781 ( .A(n119), .B(n676), .C(n603), .Q(n138) );
  NOR21 U782 ( .A(n594), .B(n139), .Q(N495) );
  AOI211 U783 ( .A(n140), .B(n687), .C(n603), .Q(n139) );
  NOR21 U784 ( .A(n594), .B(n141), .Q(N494) );
  AOI211 U785 ( .A(n140), .B(n675), .C(n603), .Q(n141) );
  NOR21 U786 ( .A(n594), .B(n142), .Q(N493) );
  AOI211 U787 ( .A(n140), .B(n683), .C(n603), .Q(n142) );
  NOR21 U788 ( .A(n594), .B(n143), .Q(N492) );
  AOI211 U789 ( .A(n140), .B(n679), .C(n603), .Q(n143) );
  NOR21 U790 ( .A(n594), .B(n144), .Q(N491) );
  AOI211 U791 ( .A(n140), .B(n686), .C(n602), .Q(n144) );
  NOR21 U792 ( .A(n594), .B(n145), .Q(N490) );
  AOI211 U793 ( .A(n140), .B(n674), .C(n603), .Q(n145) );
  NOR21 U794 ( .A(n594), .B(n149), .Q(N489) );
  AOI211 U795 ( .A(n140), .B(n682), .C(n603), .Q(n149) );
  NOR21 U796 ( .A(n594), .B(n150), .Q(N488) );
  AOI211 U797 ( .A(n140), .B(n678), .C(n603), .Q(n150) );
  NOR21 U798 ( .A(n595), .B(n151), .Q(N487) );
  AOI211 U799 ( .A(n140), .B(n685), .C(n603), .Q(n151) );
  NOR21 U800 ( .A(n595), .B(n152), .Q(N486) );
  AOI211 U801 ( .A(n140), .B(n673), .C(n603), .Q(n152) );
  NOR21 U802 ( .A(n595), .B(n153), .Q(N485) );
  AOI211 U803 ( .A(n140), .B(n681), .C(n603), .Q(n153) );
  NOR21 U804 ( .A(n595), .B(n154), .Q(N484) );
  AOI211 U805 ( .A(n140), .B(n677), .C(n603), .Q(n154) );
  NOR21 U806 ( .A(n595), .B(n155), .Q(N483) );
  AOI211 U807 ( .A(n140), .B(n684), .C(n601), .Q(n155) );
  NOR21 U808 ( .A(n595), .B(n156), .Q(N482) );
  AOI211 U809 ( .A(n140), .B(n672), .C(n602), .Q(n156) );
  NOR21 U810 ( .A(n595), .B(n157), .Q(N481) );
  AOI211 U811 ( .A(n140), .B(n680), .C(n603), .Q(n157) );
  NOR21 U812 ( .A(n595), .B(n158), .Q(N480) );
  AOI211 U813 ( .A(n140), .B(n676), .C(n603), .Q(n158) );
  NOR21 U814 ( .A(n595), .B(n167), .Q(N479) );
  AOI211 U815 ( .A(n168), .B(n687), .C(n601), .Q(n167) );
  NOR21 U816 ( .A(n595), .B(n169), .Q(N478) );
  AOI211 U817 ( .A(n168), .B(n675), .C(n602), .Q(n169) );
  NOR21 U818 ( .A(n595), .B(n170), .Q(N477) );
  AOI211 U819 ( .A(n168), .B(n683), .C(n603), .Q(n170) );
  NOR21 U820 ( .A(n595), .B(n171), .Q(N476) );
  AOI211 U821 ( .A(n168), .B(n679), .C(n601), .Q(n171) );
  NOR21 U822 ( .A(n595), .B(n172), .Q(N475) );
  AOI211 U823 ( .A(n168), .B(n686), .C(n601), .Q(n172) );
  NOR21 U824 ( .A(n596), .B(n174), .Q(N472) );
  AOI211 U825 ( .A(n168), .B(n682), .C(n602), .Q(n174) );
  NOR21 U826 ( .A(n596), .B(n175), .Q(N471) );
  AOI211 U827 ( .A(n168), .B(n678), .C(n603), .Q(n175) );
  NOR21 U828 ( .A(n596), .B(n176), .Q(N470) );
  AOI211 U829 ( .A(n168), .B(n685), .C(n602), .Q(n176) );
  NOR21 U830 ( .A(n596), .B(n180), .Q(N469) );
  AOI211 U831 ( .A(n168), .B(n673), .C(n601), .Q(n180) );
  NOR21 U832 ( .A(n596), .B(n181), .Q(N468) );
  AOI211 U833 ( .A(n168), .B(n681), .C(n602), .Q(n181) );
  NOR21 U834 ( .A(n596), .B(n182), .Q(N467) );
  AOI211 U835 ( .A(n168), .B(n677), .C(n603), .Q(n182) );
  NOR21 U836 ( .A(n596), .B(n183), .Q(N466) );
  AOI211 U837 ( .A(n168), .B(n684), .C(n603), .Q(n183) );
  NOR21 U838 ( .A(n596), .B(n184), .Q(N465) );
  AOI211 U839 ( .A(n168), .B(n672), .C(n601), .Q(n184) );
  NOR21 U840 ( .A(n596), .B(n185), .Q(N464) );
  AOI211 U841 ( .A(n168), .B(n680), .C(n602), .Q(n185) );
  NOR21 U842 ( .A(n596), .B(n186), .Q(N463) );
  AOI211 U843 ( .A(n168), .B(n676), .C(n601), .Q(n186) );
  NOR21 U844 ( .A(n596), .B(n187), .Q(N462) );
  AOI211 U845 ( .A(n188), .B(n687), .C(n602), .Q(n187) );
  NOR21 U846 ( .A(n596), .B(n189), .Q(N461) );
  AOI211 U847 ( .A(n188), .B(n675), .C(n603), .Q(n189) );
  NOR21 U848 ( .A(n597), .B(n190), .Q(N460) );
  AOI211 U849 ( .A(n188), .B(n683), .C(n603), .Q(n190) );
  NOR21 U850 ( .A(n597), .B(n191), .Q(N459) );
  AOI211 U851 ( .A(n188), .B(n679), .C(n603), .Q(n191) );
  NOR21 U852 ( .A(n597), .B(n192), .Q(N458) );
  AOI211 U853 ( .A(n188), .B(n686), .C(n601), .Q(n192) );
  NOR21 U854 ( .A(n597), .B(n193), .Q(N457) );
  AOI211 U855 ( .A(n188), .B(n674), .C(n602), .Q(n193) );
  NOR21 U856 ( .A(n597), .B(n194), .Q(N456) );
  AOI211 U857 ( .A(n188), .B(n682), .C(n603), .Q(n194) );
  NOR21 U858 ( .A(n597), .B(n195), .Q(N455) );
  AOI211 U859 ( .A(n188), .B(n678), .C(n601), .Q(n195) );
  NOR21 U860 ( .A(n597), .B(n196), .Q(N454) );
  AOI211 U861 ( .A(n188), .B(n685), .C(n601), .Q(n196) );
  NOR21 U862 ( .A(n597), .B(n197), .Q(N453) );
  AOI211 U863 ( .A(n188), .B(n673), .C(n601), .Q(n197) );
  NOR21 U864 ( .A(n597), .B(n198), .Q(N452) );
  AOI211 U865 ( .A(n188), .B(n681), .C(n602), .Q(n198) );
  NOR21 U866 ( .A(n597), .B(n199), .Q(N451) );
  AOI211 U867 ( .A(n188), .B(n677), .C(n603), .Q(n199) );
  NOR21 U868 ( .A(n597), .B(n200), .Q(N450) );
  AOI211 U869 ( .A(n188), .B(n684), .C(n602), .Q(n200) );
  NOR21 U870 ( .A(n597), .B(n201), .Q(N449) );
  AOI211 U871 ( .A(n188), .B(n672), .C(n602), .Q(n201) );
  NOR21 U872 ( .A(n597), .B(n203), .Q(N446) );
  AOI211 U873 ( .A(n188), .B(n676), .C(n601), .Q(n203) );
  NOR21 U874 ( .A(n593), .B(n204), .Q(N445) );
  AOI211 U875 ( .A(n205), .B(n687), .C(n601), .Q(n204) );
  NOR21 U876 ( .A(n596), .B(n206), .Q(N444) );
  AOI211 U877 ( .A(n205), .B(n675), .C(n602), .Q(n206) );
  NOR21 U878 ( .A(n597), .B(n207), .Q(N443) );
  AOI211 U879 ( .A(n205), .B(n683), .C(n603), .Q(n207) );
  NOR21 U880 ( .A(n593), .B(n208), .Q(N442) );
  AOI211 U881 ( .A(n205), .B(n679), .C(n601), .Q(n208) );
  NOR21 U882 ( .A(n596), .B(n209), .Q(N441) );
  AOI211 U883 ( .A(n205), .B(n686), .C(n602), .Q(n209) );
  NOR21 U884 ( .A(n597), .B(n210), .Q(N440) );
  AOI211 U885 ( .A(n205), .B(n674), .C(n603), .Q(n210) );
  NOR21 U886 ( .A(n595), .B(n211), .Q(N439) );
  AOI211 U887 ( .A(n205), .B(n682), .C(n601), .Q(n211) );
  NOR21 U888 ( .A(n593), .B(n212), .Q(N438) );
  AOI211 U889 ( .A(n205), .B(n678), .C(n602), .Q(n212) );
  NOR21 U890 ( .A(n596), .B(n213), .Q(N437) );
  AOI211 U891 ( .A(n205), .B(n685), .C(n603), .Q(n213) );
  NOR21 U892 ( .A(n597), .B(n214), .Q(N436) );
  AOI211 U893 ( .A(n205), .B(n673), .C(n601), .Q(n214) );
  NOR21 U894 ( .A(n595), .B(n215), .Q(N435) );
  AOI211 U895 ( .A(n205), .B(n681), .C(n602), .Q(n215) );
  NOR21 U896 ( .A(n593), .B(n216), .Q(N434) );
  AOI211 U897 ( .A(n205), .B(n677), .C(n603), .Q(n216) );
  NOR21 U898 ( .A(n596), .B(n217), .Q(N433) );
  AOI211 U899 ( .A(n205), .B(n684), .C(n601), .Q(n217) );
  NOR21 U900 ( .A(n598), .B(n218), .Q(N432) );
  AOI211 U901 ( .A(n205), .B(n672), .C(n602), .Q(n218) );
  NOR21 U902 ( .A(n598), .B(n219), .Q(N431) );
  AOI211 U903 ( .A(n205), .B(n680), .C(n603), .Q(n219) );
  NOR21 U904 ( .A(n598), .B(n220), .Q(N430) );
  AOI211 U905 ( .A(n205), .B(n676), .C(n601), .Q(n220) );
  NOR21 U906 ( .A(n598), .B(n221), .Q(N429) );
  AOI211 U907 ( .A(n222), .B(n687), .C(n602), .Q(n221) );
  NOR21 U908 ( .A(n598), .B(n223), .Q(N428) );
  AOI211 U909 ( .A(n222), .B(n675), .C(n603), .Q(n223) );
  NOR21 U910 ( .A(n598), .B(n224), .Q(N427) );
  AOI211 U911 ( .A(n222), .B(n683), .C(n601), .Q(n224) );
  NOR21 U912 ( .A(n598), .B(n225), .Q(N426) );
  AOI211 U913 ( .A(n222), .B(n679), .C(n603), .Q(n225) );
  NOR21 U914 ( .A(n598), .B(n226), .Q(N425) );
  AOI211 U915 ( .A(n222), .B(n686), .C(n601), .Q(n226) );
  NOR21 U916 ( .A(n598), .B(n227), .Q(N424) );
  AOI211 U917 ( .A(n222), .B(n674), .C(n603), .Q(n227) );
  NOR21 U918 ( .A(n598), .B(n228), .Q(N423) );
  AOI211 U919 ( .A(n222), .B(n682), .C(n601), .Q(n228) );
  NOR21 U920 ( .A(n598), .B(n230), .Q(N420) );
  AOI211 U921 ( .A(n222), .B(n685), .C(n602), .Q(n230) );
  NOR21 U922 ( .A(n598), .B(n231), .Q(N419) );
  AOI211 U923 ( .A(n222), .B(n673), .C(n603), .Q(n231) );
  NOR21 U924 ( .A(n599), .B(n232), .Q(N418) );
  AOI211 U925 ( .A(n222), .B(n681), .C(n601), .Q(n232) );
  NOR21 U926 ( .A(n598), .B(n233), .Q(N417) );
  AOI211 U927 ( .A(n222), .B(n677), .C(n601), .Q(n233) );
  NOR21 U928 ( .A(n599), .B(n234), .Q(N416) );
  AOI211 U929 ( .A(n222), .B(n684), .C(n601), .Q(n234) );
  NOR21 U930 ( .A(n599), .B(n235), .Q(N415) );
  AOI211 U931 ( .A(n222), .B(n672), .C(n601), .Q(n235) );
  NOR21 U932 ( .A(n599), .B(n236), .Q(N414) );
  AOI211 U933 ( .A(n222), .B(n680), .C(n602), .Q(n236) );
  NOR21 U934 ( .A(n599), .B(n237), .Q(N413) );
  AOI211 U935 ( .A(n222), .B(n676), .C(n603), .Q(n237) );
  NOR21 U936 ( .A(n599), .B(n238), .Q(N412) );
  AOI211 U937 ( .A(n525), .B(n687), .C(n601), .Q(n238) );
  NOR21 U938 ( .A(n599), .B(n243), .Q(N411) );
  AOI211 U939 ( .A(n525), .B(n675), .C(n602), .Q(n243) );
  NOR21 U940 ( .A(n599), .B(n246), .Q(N410) );
  AOI211 U941 ( .A(n239), .B(n683), .C(n602), .Q(n246) );
  NOR21 U942 ( .A(n599), .B(n249), .Q(N409) );
  AOI211 U943 ( .A(n525), .B(n679), .C(n601), .Q(n249) );
  NOR21 U944 ( .A(n599), .B(n252), .Q(N408) );
  AOI211 U945 ( .A(n525), .B(n686), .C(n602), .Q(n252) );
  NOR21 U946 ( .A(n599), .B(n255), .Q(N407) );
  AOI211 U947 ( .A(n525), .B(n674), .C(n603), .Q(n255) );
  NOR21 U948 ( .A(n599), .B(n257), .Q(N406) );
  AOI211 U949 ( .A(n239), .B(n682), .C(n601), .Q(n257) );
  NOR21 U950 ( .A(n599), .B(n259), .Q(N405) );
  AOI211 U951 ( .A(n525), .B(n678), .C(n602), .Q(n259) );
  NOR21 U952 ( .A(n106), .B(n592), .Q(N524) );
  AOI211 U953 ( .A(n102), .B(n686), .C(n601), .Q(n106) );
  NOR21 U954 ( .A(n173), .B(n594), .Q(N474) );
  AOI211 U955 ( .A(n674), .B(n168), .C(n602), .Q(n173) );
  NOR21 U956 ( .A(n202), .B(n598), .Q(N448) );
  AOI211 U957 ( .A(n680), .B(n188), .C(n602), .Q(n202) );
  NOR21 U958 ( .A(n229), .B(n599), .Q(N422) );
  AOI211 U959 ( .A(n678), .B(n222), .C(n602), .Q(n229) );
  NOR21 U960 ( .A(n594), .B(n261), .Q(N404) );
  AOI211 U961 ( .A(n239), .B(n685), .C(n603), .Q(n261) );
  NOR21 U962 ( .A(n598), .B(n264), .Q(N403) );
  AOI211 U963 ( .A(n525), .B(n673), .C(n603), .Q(n264) );
  NOR21 U964 ( .A(n599), .B(n266), .Q(N402) );
  AOI211 U965 ( .A(n239), .B(n681), .C(n603), .Q(n266) );
  NOR21 U966 ( .A(n594), .B(n268), .Q(N401) );
  AOI211 U967 ( .A(n525), .B(n677), .C(n603), .Q(n268) );
  NOR21 U968 ( .A(n598), .B(n270), .Q(N400) );
  AOI211 U969 ( .A(n239), .B(n684), .C(n603), .Q(n270) );
  NOR21 U970 ( .A(n599), .B(n273), .Q(N399) );
  AOI211 U971 ( .A(n525), .B(n672), .C(n601), .Q(n273) );
  NOR21 U972 ( .A(n595), .B(n275), .Q(N398) );
  AOI211 U973 ( .A(n525), .B(n680), .C(n602), .Q(n275) );
  NOR21 U974 ( .A(n286), .B(n668), .Q(N229) );
  INV3 U975 ( .A(N215), .Q(n668) );
  NOR21 U976 ( .A(n286), .B(n669), .Q(N228) );
  INV3 U977 ( .A(N214), .Q(n669) );
  NOR21 U978 ( .A(n286), .B(n670), .Q(N227) );
  INV3 U979 ( .A(N213), .Q(n670) );
  NOR21 U980 ( .A(n286), .B(n671), .Q(N226) );
  INV3 U981 ( .A(N212), .Q(n671) );
  INV3 U982 ( .A(n526), .Q(n527) );
  INV3 U983 ( .A(n287), .Q(n662) );
  INV3 U984 ( .A(n239), .Q(n524) );
  NOR31 U985 ( .A(n488), .B(n486), .C(n485), .Q(n239) );
  INV3 U986 ( .A(n133), .Q(n666) );
  INV3 U987 ( .A(n298), .Q(n623) );
  AOI221 U988 ( .A(N143), .B(n279), .C(N134), .D(n292), .Q(n298) );
  INV3 U989 ( .A(n297), .Q(n624) );
  AOI221 U990 ( .A(N144), .B(n279), .C(N135), .D(n292), .Q(n297) );
  INV3 U991 ( .A(n296), .Q(n625) );
  AOI221 U992 ( .A(N145), .B(n279), .C(N136), .D(n292), .Q(n296) );
  INV3 U993 ( .A(n299), .Q(n622) );
  AOI221 U994 ( .A(n499), .B(n279), .C(N133), .D(n292), .Q(n299) );
  BUF2 U995 ( .A(n523), .Q(n610) );
  INV3 U996 ( .A(n310), .Q(n635) );
  NAND22 U997 ( .A(n281), .B(N123), .Q(n310) );
  INV3 U998 ( .A(n311), .Q(n634) );
  NAND22 U999 ( .A(n281), .B(N122), .Q(n311) );
  INV3 U1000 ( .A(n312), .Q(n633) );
  NAND22 U1001 ( .A(n281), .B(N121), .Q(n312) );
  NOR21 U1002 ( .A(n510), .B(n601), .Q(n281) );
  NAND22 U1003 ( .A(n179), .B(n489), .Q(n147) );
  NOR21 U1004 ( .A(n601), .B(n97), .Q(N381) );
  NOR21 U1005 ( .A(n601), .B(n98), .Q(N382) );
  INV3 U1006 ( .A(n313), .Q(n632) );
  NAND22 U1007 ( .A(n281), .B(N120), .Q(n313) );
  INV3 U1008 ( .A(n314), .Q(n631) );
  NAND22 U1009 ( .A(n281), .B(N119), .Q(n314) );
  INV3 U1010 ( .A(n315), .Q(n630) );
  NAND22 U1011 ( .A(n281), .B(n494), .Q(n315) );
  INV3 U1012 ( .A(n289), .Q(n648) );
  AOI2111 U1013 ( .A(N138), .B(n712), .C(N140), .D(N139), .Q(N390) );
  NAND22 U1014 ( .A(n711), .B(n710), .Q(n712) );
  NOR21 U1015 ( .A(N134), .B(N133), .Q(n711) );
  NOR31 U1016 ( .A(N135), .B(N137), .C(N136), .Q(n710) );
  BUF2 U1017 ( .A(n650), .Q(n543) );
  BUF2 U1018 ( .A(n651), .Q(n559) );
  BUF2 U1019 ( .A(n652), .Q(n575) );
  BUF2 U1020 ( .A(n653), .Q(n591) );
  BUF2 U1021 ( .A(n650), .Q(n542) );
  BUF2 U1022 ( .A(n651), .Q(n558) );
  BUF2 U1023 ( .A(n652), .Q(n574) );
  BUF2 U1024 ( .A(n653), .Q(n590) );
  BUF2 U1025 ( .A(n650), .Q(n541) );
  BUF2 U1026 ( .A(n651), .Q(n557) );
  BUF2 U1027 ( .A(n652), .Q(n573) );
  BUF2 U1028 ( .A(n653), .Q(n589) );
  BUF2 U1029 ( .A(n650), .Q(n540) );
  BUF2 U1030 ( .A(n651), .Q(n556) );
  BUF2 U1031 ( .A(n652), .Q(n572) );
  BUF2 U1032 ( .A(n653), .Q(n588) );
  BUF2 U1033 ( .A(n650), .Q(n539) );
  BUF2 U1034 ( .A(n651), .Q(n555) );
  BUF2 U1035 ( .A(n652), .Q(n571) );
  BUF2 U1036 ( .A(n653), .Q(n587) );
  BUF2 U1037 ( .A(n650), .Q(n538) );
  BUF2 U1038 ( .A(n651), .Q(n554) );
  BUF2 U1039 ( .A(n652), .Q(n570) );
  BUF2 U1040 ( .A(n653), .Q(n586) );
  BUF2 U1041 ( .A(n650), .Q(n537) );
  BUF2 U1042 ( .A(n651), .Q(n553) );
  BUF2 U1043 ( .A(n652), .Q(n569) );
  BUF2 U1044 ( .A(n653), .Q(n585) );
  BUF2 U1045 ( .A(n650), .Q(n536) );
  BUF2 U1046 ( .A(n651), .Q(n552) );
  BUF2 U1047 ( .A(n652), .Q(n568) );
  BUF2 U1048 ( .A(n653), .Q(n584) );
  BUF2 U1049 ( .A(n650), .Q(n535) );
  BUF2 U1050 ( .A(n651), .Q(n551) );
  BUF2 U1051 ( .A(n652), .Q(n567) );
  BUF2 U1052 ( .A(n653), .Q(n583) );
  BUF2 U1053 ( .A(n650), .Q(n534) );
  BUF2 U1054 ( .A(n651), .Q(n550) );
  BUF2 U1055 ( .A(n652), .Q(n566) );
  BUF2 U1056 ( .A(n653), .Q(n582) );
  BUF2 U1057 ( .A(n650), .Q(n533) );
  BUF2 U1058 ( .A(n651), .Q(n549) );
  BUF2 U1059 ( .A(n652), .Q(n565) );
  BUF2 U1060 ( .A(n653), .Q(n581) );
  BUF2 U1061 ( .A(n650), .Q(n532) );
  BUF2 U1062 ( .A(n651), .Q(n548) );
  BUF2 U1063 ( .A(n652), .Q(n564) );
  BUF2 U1064 ( .A(n653), .Q(n580) );
  BUF2 U1065 ( .A(n650), .Q(n531) );
  BUF2 U1066 ( .A(n651), .Q(n547) );
  BUF2 U1067 ( .A(n652), .Q(n563) );
  BUF2 U1068 ( .A(n653), .Q(n579) );
  BUF2 U1069 ( .A(n650), .Q(n530) );
  BUF2 U1070 ( .A(n651), .Q(n546) );
  BUF2 U1071 ( .A(n652), .Q(n562) );
  BUF2 U1072 ( .A(n653), .Q(n578) );
  BUF2 U1073 ( .A(n650), .Q(n529) );
  BUF2 U1074 ( .A(n651), .Q(n545) );
  BUF2 U1075 ( .A(n652), .Q(n561) );
  BUF2 U1076 ( .A(n653), .Q(n577) );
  BUF2 U1077 ( .A(n650), .Q(n528) );
  BUF2 U1078 ( .A(n651), .Q(n544) );
  BUF2 U1079 ( .A(n652), .Q(n560) );
  BUF2 U1080 ( .A(n653), .Q(n576) );
  INV3 U1081 ( .A(n702), .Q(n656) );
  NAND22 U1082 ( .A(n493), .B(n703), .Q(n702) );
  INV3 U1083 ( .A(n709), .Q(outAlmostFull) );
  AOI211 U1084 ( .A(N139), .B(N138), .C(N140), .Q(n709) );
  INV3 U1085 ( .A(n519), .Q(\r96/carry [1]) );
  NOR21 U1086 ( .A(n494), .B(outWriteCount[0]), .Q(n519) );
  XNR21 U1087 ( .A(\r96/carry [7]), .B(outWriteCount[7]), .Q(N140) );
  AOI311 U1088 ( .A(n162), .B(n148), .C(n177), .D(n601), .Q(N47) );
  AOI221 U1089 ( .A(n178), .B(n163), .C(n664), .D(N375), .Q(n177) );
  NOR21 U1090 ( .A(currentState[2]), .B(n517), .Q(n178) );
  INV3 U1091 ( .A(n147), .Q(n664) );
  INV3 U1092 ( .A(n291), .Q(n629) );
  AOI221 U1093 ( .A(N149), .B(n279), .C(N140), .D(n292), .Q(n291) );
  XOR21 U1094 ( .A(\add_263/carry [7]), .B(outWriteCount[7]), .Q(N149) );
  BUF2 U1095 ( .A(N38), .Q(n523) );
  XNR21 U1096 ( .A(\add_357/carry [6]), .B(j_FIFO[6]), .Q(n516) );
  INV3 U1097 ( .A(n309), .Q(n636) );
  NAND22 U1098 ( .A(n281), .B(N124), .Q(n309) );
  XOR21 U1099 ( .A(\add_252/carry [6]), .B(outReadCount[6]), .Q(N124) );
  INV3 U1100 ( .A(n302), .Q(n647) );
  NAND22 U1101 ( .A(N131), .B(inReset), .Q(n302) );
  XOR21 U1102 ( .A(\add_253/carry [6]), .B(N43), .Q(N131) );
  INV3 U1103 ( .A(n288), .Q(n649) );
  NAND22 U1104 ( .A(N204), .B(inReset), .Q(n288) );
  INV3 U1105 ( .A(n303), .Q(n646) );
  NAND22 U1106 ( .A(N130), .B(inReset), .Q(n303) );
  INV3 U1107 ( .A(n304), .Q(n645) );
  NAND22 U1108 ( .A(N129), .B(inReset), .Q(n304) );
  NAND22 U1109 ( .A(inReset), .B(n287), .Q(n286) );
  NAND31 U1110 ( .A(currentState[1]), .B(n505), .C(n666), .Q(n162) );
  AOI311 U1111 ( .A(n701), .B(n699), .C(n698), .D(outWriteCount[7]), .Q(n700)
         );
  OAI2111 U1112 ( .A(outReadCount[5]), .B(n508), .C(n697), .D(n696), .Q(n698)
         );
  NAND22 U1113 ( .A(outWriteCount[4]), .B(n496), .Q(n696) );
  XNR21 U1114 ( .A(outWriteCount[0]), .B(n494), .Q(N133) );
  NOR21 U1115 ( .A(j_FIFO[3]), .B(j_FIFO[2]), .Q(n242) );
  NOR21 U1116 ( .A(j_FIFO[1]), .B(j_FIFO[0]), .Q(n241) );
  NOR21 U1117 ( .A(n511), .B(j_FIFO[0]), .Q(n248) );
  NOR21 U1118 ( .A(n490), .B(j_FIFO[1]), .Q(n245) );
  NOR21 U1119 ( .A(n133), .B(currentState[1]), .Q(n99) );
  NAND22 U1120 ( .A(n300), .B(n301), .Q(n287) );
  NOR40 U1121 ( .A(outWriteCount[2]), .B(outWriteCount[1]), .C(
        outWriteCount[0]), .D(n504), .Q(n300) );
  NOR40 U1122 ( .A(outWriteCount[6]), .B(outWriteCount[5]), .C(
        outWriteCount[4]), .D(outWriteCount[3]), .Q(n301) );
  BUF2 U1123 ( .A(N40), .Q(n604) );
  OAI2111 U1124 ( .A(n695), .B(n694), .C(n693), .D(n692), .Q(n697) );
  NOR21 U1125 ( .A(outReadCount[3]), .B(n507), .Q(n695) );
  OAI2111 U1126 ( .A(n690), .B(n493), .C(n655), .D(n689), .Q(n691) );
  NAND22 U1127 ( .A(currentState[2]), .B(n489), .Q(n133) );
  NOR21 U1128 ( .A(n491), .B(j_FIFO[3]), .Q(n254) );
  NOR21 U1129 ( .A(n512), .B(j_FIFO[2]), .Q(n263) );
  NOR21 U1130 ( .A(n513), .B(currentState[2]), .Q(n166) );
  BUF2 U1131 ( .A(N40), .Q(n605) );
  BUF2 U1132 ( .A(N42), .Q(n520) );
  NAND22 U1133 ( .A(outReadCount[6]), .B(n506), .Q(n701) );
  NOR31 U1134 ( .A(n486), .B(j_FIFO[6]), .C(n488), .Q(n168) );
  AOI211 U1135 ( .A(n163), .B(n164), .C(n663), .Q(n159) );
  XNR21 U1136 ( .A(n517), .B(sig_fsm_start_W), .Q(n164) );
  NOR21 U1137 ( .A(\os2/sigQout2 ), .B(n515), .Q(sig_fsm_start_W) );
  NAND22 U1138 ( .A(n99), .B(inReset), .Q(n161) );
  NAND22 U1139 ( .A(outReadCount[3]), .B(n507), .Q(n692) );
  NAND31 U1140 ( .A(n96), .B(n97), .C(inReset), .Q(N532) );
  NAND31 U1141 ( .A(n96), .B(n98), .C(inReset), .Q(N530) );
  NAND22 U1142 ( .A(outReadCount[2]), .B(n500), .Q(n689) );
  NOR21 U1143 ( .A(n499), .B(outReadCount[0]), .Q(n690) );
  NAND22 U1144 ( .A(inReset), .B(n162), .Q(N199) );
  NAND22 U1145 ( .A(outReadCount[4]), .B(n509), .Q(n693) );
  NOR21 U1146 ( .A(n286), .B(j_FIFO[0]), .Q(N225) );
  INV3 U1147 ( .A(n102), .Q(n526) );
  NOR31 U1148 ( .A(j_FIFO[5]), .B(j_FIFO[6]), .C(j_FIFO[4]), .Q(n102) );
  NOR31 U1149 ( .A(j_FIFO[5]), .B(j_FIFO[6]), .C(n486), .Q(n119) );
  NOR31 U1150 ( .A(j_FIFO[4]), .B(j_FIFO[6]), .C(n488), .Q(n140) );
  NOR31 U1151 ( .A(j_FIFO[4]), .B(j_FIFO[5]), .C(n485), .Q(n188) );
  BUF2 U1152 ( .A(N41), .Q(n521) );
  NOR31 U1153 ( .A(n486), .B(j_FIFO[5]), .C(n485), .Q(n205) );
  NOR31 U1154 ( .A(n488), .B(j_FIFO[4]), .C(n485), .Q(n222) );
  INV3 U1155 ( .A(n160), .Q(n621) );
  INV3 U1156 ( .A(n688), .Q(n655) );
  AOI211 U1157 ( .A(n493), .B(n690), .C(outWriteCount[1]), .Q(n688) );
  INV3 U1158 ( .A(n305), .Q(n644) );
  NAND22 U1159 ( .A(N128), .B(inReset), .Q(n305) );
  INV3 U1160 ( .A(n306), .Q(n643) );
  NAND22 U1161 ( .A(N127), .B(inReset), .Q(n306) );
  INV3 U1162 ( .A(n307), .Q(n642) );
  NAND22 U1163 ( .A(N126), .B(inReset), .Q(n307) );
  NAND22 U1164 ( .A(inReset), .B(n510), .Q(N396) );
  NAND31 U1165 ( .A(currentState[3]), .B(n505), .C(n166), .Q(n97) );
  NOR31 U1166 ( .A(currentState[1]), .B(currentState[2]), .C(n505), .Q(n179)
         );
  NOR31 U1167 ( .A(currentState[1]), .B(currentState[3]), .C(currentState[0]), 
        .Q(n163) );
  NAND22 U1168 ( .A(n179), .B(currentState[3]), .Q(n98) );
  NAND22 U1169 ( .A(outReadCount[5]), .B(n508), .Q(n699) );
  AOI221 U1170 ( .A(n289), .B(n290), .C(n514), .D(n492), .Q(N190) );
  NAND22 U1171 ( .A(inReset), .B(n492), .Q(n290) );
  NAND22 U1172 ( .A(inReset), .B(n514), .Q(n289) );
  INV3 U1173 ( .A(n165), .Q(n663) );
  NAND31 U1174 ( .A(n166), .B(n489), .C(currentState[0]), .Q(n165) );
  NAND22 U1175 ( .A(n518), .B(\os1/sigQout1 ), .Q(n517) );
  INV3 U1176 ( .A(n308), .Q(n641) );
  NAND22 U1177 ( .A(n502), .B(inReset), .Q(n308) );
  INV3 U1178 ( .A(n713), .Q(n637) );
  NAND22 U1179 ( .A(inReset), .B(\os1/sigQout1 ), .Q(n713) );
  INV3 U1180 ( .A(n715), .Q(n639) );
  NAND22 U1181 ( .A(inReset), .B(\os2/sigQout1 ), .Q(n715) );
  INV3 U1182 ( .A(n285), .Q(n650) );
  NAND22 U1183 ( .A(inData[0]), .B(inReset), .Q(n285) );
  INV3 U1184 ( .A(n284), .Q(n651) );
  NAND22 U1185 ( .A(inData[1]), .B(inReset), .Q(n284) );
  INV3 U1186 ( .A(n283), .Q(n652) );
  NAND22 U1187 ( .A(inData[2]), .B(inReset), .Q(n283) );
  INV3 U1188 ( .A(n282), .Q(n653) );
  NAND22 U1189 ( .A(inData[3]), .B(inReset), .Q(n282) );
  INV3 U1190 ( .A(inReset), .Q(n602) );
  INV3 U1191 ( .A(inReset), .Q(n603) );
  INV3 U1192 ( .A(inReset), .Q(n601) );
  NOR40 U1193 ( .A(currentState[2]), .B(currentState[1]), .C(currentState[0]), 
        .D(n489), .Q(outDone) );
  NOR40 U1194 ( .A(n705), .B(n706), .C(n661), .D(n704), .Q(N391) );
  INV3 U1195 ( .A(n701), .Q(n661) );
  AOI211 U1196 ( .A(outWriteCount[1]), .B(n703), .C(n656), .Q(n704) );
  NAND41 U1197 ( .A(n699), .B(n693), .C(n692), .D(n689), .Q(n705) );
  NAND22 U1198 ( .A(outReadCount[0]), .B(n499), .Q(n703) );
  INV3 U1199 ( .A(n714), .Q(n638) );
  NAND22 U1200 ( .A(inReset), .B(inWriteEnable), .Q(n714) );
  INV3 U1201 ( .A(\os1/dff1/n2 ), .Q(n640) );
  NAND22 U1202 ( .A(inReset), .B(inReadEnable), .Q(\os1/dff1/n2 ) );
  OAI212 U1203 ( .A(outReadCount[2]), .B(n500), .C(n691), .Q(n694) );
  OAI212 U1204 ( .A(outReadCount[6]), .B(n506), .C(n700), .Q(n706) );
endmodule

