`timescale 1ns / 1ps

 
module tb_MUX();

parameter	CLK_PERIOD = 20 ; 

reg	[1  : 0]	inData211	;
reg	    	    inSel211	;
reg	    	    outData211	;

reg [15 : 0]    inData414	;
reg	[1  : 0]	inSel414	;
reg	[3  : 0] 	outData414	;

reg	[7  : 0]	inData811	;
reg	[2  : 0]	inSel811	;
reg	        	outData811	;


MUX211 u_mux211 (
	.inData			(inData211	), 
	.inSel			(inSel211	),
	.outData		(outData211	)
);

MUX414 u_mux414 (
	.inData			(inData414	), 
	.inSel			(inSel414	),
	.outData		(outData414	)
);

MUX811 u_mux811 (
	.inData			(inData811	), 
	.inSel			(inSel811	),
	.outData		(outData811	)
);

initial begin 
	inData211 = 2'b0;
	inSel211  = 1'b0;

	inData414 = 16'b0;
	inSel414  = 2'b0;

	inData811 = 8'b0;
	inSel811  = 3'b0;
end


always begin : SEL

    inSel211  = 1'b0; inSel414  = 2'b00; inSel811  = 3'b000;
	#CLK_PERIOD ; #CLK_PERIOD ; #CLK_PERIOD ; #CLK_PERIOD ;
	#CLK_PERIOD ; #CLK_PERIOD ; #CLK_PERIOD ; #CLK_PERIOD ;
	#CLK_PERIOD ; #CLK_PERIOD ; #CLK_PERIOD ; #CLK_PERIOD ;
	#CLK_PERIOD ; #CLK_PERIOD ; #CLK_PERIOD ; #CLK_PERIOD ;
	#CLK_PERIOD ; #CLK_PERIOD ; #CLK_PERIOD ; #CLK_PERIOD ;
	#CLK_PERIOD ; #CLK_PERIOD ; #CLK_PERIOD ; #CLK_PERIOD ;
	#CLK_PERIOD ; #CLK_PERIOD ; #CLK_PERIOD ; #CLK_PERIOD ;
	#CLK_PERIOD ; #CLK_PERIOD ; #CLK_PERIOD ; #CLK_PERIOD ;

    inSel211  = 1'b1; inSel414  = 2'b01; inSel811  = 3'b001;
	#CLK_PERIOD ; #CLK_PERIOD ; #CLK_PERIOD ; #CLK_PERIOD ;
	#CLK_PERIOD ; #CLK_PERIOD ; #CLK_PERIOD ; #CLK_PERIOD ;
	#CLK_PERIOD ; #CLK_PERIOD ; #CLK_PERIOD ; #CLK_PERIOD ;
	#CLK_PERIOD ; #CLK_PERIOD ; #CLK_PERIOD ; #CLK_PERIOD ;
	#CLK_PERIOD ; #CLK_PERIOD ; #CLK_PERIOD ; #CLK_PERIOD ;
	#CLK_PERIOD ; #CLK_PERIOD ; #CLK_PERIOD ; #CLK_PERIOD ;
	#CLK_PERIOD ; #CLK_PERIOD ; #CLK_PERIOD ; #CLK_PERIOD ;
	#CLK_PERIOD ; #CLK_PERIOD ; #CLK_PERIOD ; #CLK_PERIOD ;
    
    inSel211  = 1'b0; inSel414  = 2'b10; inSel811  = 3'b010;
	#CLK_PERIOD ; #CLK_PERIOD ; #CLK_PERIOD ; #CLK_PERIOD ;
	#CLK_PERIOD ; #CLK_PERIOD ; #CLK_PERIOD ; #CLK_PERIOD ;
	#CLK_PERIOD ; #CLK_PERIOD ; #CLK_PERIOD ; #CLK_PERIOD ;
	#CLK_PERIOD ; #CLK_PERIOD ; #CLK_PERIOD ; #CLK_PERIOD ;
	#CLK_PERIOD ; #CLK_PERIOD ; #CLK_PERIOD ; #CLK_PERIOD ;
	#CLK_PERIOD ; #CLK_PERIOD ; #CLK_PERIOD ; #CLK_PERIOD ;
	#CLK_PERIOD ; #CLK_PERIOD ; #CLK_PERIOD ; #CLK_PERIOD ;
	#CLK_PERIOD ; #CLK_PERIOD ; #CLK_PERIOD ; #CLK_PERIOD ;
    
    inSel211  = 1'b1; inSel414  = 2'b11; inSel811  = 3'b011;
	#CLK_PERIOD ; #CLK_PERIOD ; #CLK_PERIOD ; #CLK_PERIOD ;
	#CLK_PERIOD ; #CLK_PERIOD ; #CLK_PERIOD ; #CLK_PERIOD ;
	#CLK_PERIOD ; #CLK_PERIOD ; #CLK_PERIOD ; #CLK_PERIOD ;
	#CLK_PERIOD ; #CLK_PERIOD ; #CLK_PERIOD ; #CLK_PERIOD ;
	#CLK_PERIOD ; #CLK_PERIOD ; #CLK_PERIOD ; #CLK_PERIOD ;
	#CLK_PERIOD ; #CLK_PERIOD ; #CLK_PERIOD ; #CLK_PERIOD ;
	#CLK_PERIOD ; #CLK_PERIOD ; #CLK_PERIOD ; #CLK_PERIOD ;
	#CLK_PERIOD ; #CLK_PERIOD ; #CLK_PERIOD ; #CLK_PERIOD ;
    
    inSel211  = 1'b0; inSel414  = 2'b00; inSel811  = 3'b100;
	#CLK_PERIOD ; #CLK_PERIOD ; #CLK_PERIOD ; #CLK_PERIOD ;
	#CLK_PERIOD ; #CLK_PERIOD ; #CLK_PERIOD ; #CLK_PERIOD ;
	#CLK_PERIOD ; #CLK_PERIOD ; #CLK_PERIOD ; #CLK_PERIOD ;
	#CLK_PERIOD ; #CLK_PERIOD ; #CLK_PERIOD ; #CLK_PERIOD ;
	#CLK_PERIOD ; #CLK_PERIOD ; #CLK_PERIOD ; #CLK_PERIOD ;
	#CLK_PERIOD ; #CLK_PERIOD ; #CLK_PERIOD ; #CLK_PERIOD ;
	#CLK_PERIOD ; #CLK_PERIOD ; #CLK_PERIOD ; #CLK_PERIOD ;
	#CLK_PERIOD ; #CLK_PERIOD ; #CLK_PERIOD ; #CLK_PERIOD ;
    
    inSel211  = 1'b1; inSel414  = 2'b01; inSel811  = 3'b101;
	#CLK_PERIOD ; #CLK_PERIOD ; #CLK_PERIOD ; #CLK_PERIOD ;
	#CLK_PERIOD ; #CLK_PERIOD ; #CLK_PERIOD ; #CLK_PERIOD ;
	#CLK_PERIOD ; #CLK_PERIOD ; #CLK_PERIOD ; #CLK_PERIOD ;
	#CLK_PERIOD ; #CLK_PERIOD ; #CLK_PERIOD ; #CLK_PERIOD ;
	#CLK_PERIOD ; #CLK_PERIOD ; #CLK_PERIOD ; #CLK_PERIOD ;
	#CLK_PERIOD ; #CLK_PERIOD ; #CLK_PERIOD ; #CLK_PERIOD ;
	#CLK_PERIOD ; #CLK_PERIOD ; #CLK_PERIOD ; #CLK_PERIOD ;
	#CLK_PERIOD ; #CLK_PERIOD ; #CLK_PERIOD ; #CLK_PERIOD ;
    
    inSel211  = 1'b0; inSel414  = 2'b10; inSel811  = 3'b110;
	#CLK_PERIOD ; #CLK_PERIOD ; #CLK_PERIOD ; #CLK_PERIOD ;
	#CLK_PERIOD ; #CLK_PERIOD ; #CLK_PERIOD ; #CLK_PERIOD ;
	#CLK_PERIOD ; #CLK_PERIOD ; #CLK_PERIOD ; #CLK_PERIOD ;
	#CLK_PERIOD ; #CLK_PERIOD ; #CLK_PERIOD ; #CLK_PERIOD ;
	#CLK_PERIOD ; #CLK_PERIOD ; #CLK_PERIOD ; #CLK_PERIOD ;
	#CLK_PERIOD ; #CLK_PERIOD ; #CLK_PERIOD ; #CLK_PERIOD ;
	#CLK_PERIOD ; #CLK_PERIOD ; #CLK_PERIOD ; #CLK_PERIOD ;
	#CLK_PERIOD ; #CLK_PERIOD ; #CLK_PERIOD ; #CLK_PERIOD ;
    
    inSel211  = 1'b1; inSel414  = 2'b11; inSel811  = 3'b111;
	#CLK_PERIOD ; #CLK_PERIOD ; #CLK_PERIOD ; #CLK_PERIOD ;
	#CLK_PERIOD ; #CLK_PERIOD ; #CLK_PERIOD ; #CLK_PERIOD ;
	#CLK_PERIOD ; #CLK_PERIOD ; #CLK_PERIOD ; #CLK_PERIOD ;
	#CLK_PERIOD ; #CLK_PERIOD ; #CLK_PERIOD ; #CLK_PERIOD ;
	#CLK_PERIOD ; #CLK_PERIOD ; #CLK_PERIOD ; #CLK_PERIOD ;
	#CLK_PERIOD ; #CLK_PERIOD ; #CLK_PERIOD ; #CLK_PERIOD ;
	#CLK_PERIOD ; #CLK_PERIOD ; #CLK_PERIOD ; #CLK_PERIOD ;
	#CLK_PERIOD ; #CLK_PERIOD ; #CLK_PERIOD ; #CLK_PERIOD ;
    
end

always begin : DATA211

    inData211 = 2'b00;
    #CLK_PERIOD;

    inData211 = 2'b01;
    #CLK_PERIOD;

    inData211 = 2'b10;
    #CLK_PERIOD;

    inData211 = 2'b11;
    #CLK_PERIOD;

end

always begin : DATA414
    
    inData414 = 16'h00;
    #CLK_PERIOD;
    inData414 = 16'h01;
    #CLK_PERIOD;
    inData414 = 16'h02;
    #CLK_PERIOD;
    inData414 = 16'h03;
    #CLK_PERIOD;
    inData414 = 16'h04;
    #CLK_PERIOD;
    inData414 = 16'h05;
    #CLK_PERIOD;
    inData414 = 16'h06;
    #CLK_PERIOD;
    inData414 = 16'h07;
    #CLK_PERIOD;
    inData414 = 16'h08;
    #CLK_PERIOD;
    inData414 = 16'h09;
    #CLK_PERIOD;
    inData414 = 16'h0A;
    #CLK_PERIOD;
    inData414 = 16'h0B;
    #CLK_PERIOD;
    inData414 = 16'h0C;
    #CLK_PERIOD;
    inData414 = 16'h0D;
    #CLK_PERIOD;
    inData414 = 16'h0E;
    #CLK_PERIOD;
    inData414 = 16'h0F;
    #CLK_PERIOD;
    inData414 = 16'h00;
    #CLK_PERIOD;
    inData414 = 16'h10;
    #CLK_PERIOD;
    inData414 = 16'h20;
    #CLK_PERIOD;
    inData414 = 16'h30;
    #CLK_PERIOD;
    inData414 = 16'h40;
    #CLK_PERIOD;
    inData414 = 16'h50;
    #CLK_PERIOD;
    inData414 = 16'h60;
    #CLK_PERIOD;
    inData414 = 16'h70;
    #CLK_PERIOD;
    inData414 = 16'h80;
    #CLK_PERIOD;
    inData414 = 16'h90;
    #CLK_PERIOD;
    inData414 = 16'hA0;
    #CLK_PERIOD;
    inData414 = 16'hB0;
    #CLK_PERIOD;
    inData414 = 16'hC0;
    #CLK_PERIOD;
    inData414 = 16'hD0;
    #CLK_PERIOD;
    inData414 = 16'hE0;
    #CLK_PERIOD;
    inData414 = 16'hF0;
    #CLK_PERIOD;

end

always begin : DATA811
    
    inData811 = 8'h00;
    #CLK_PERIOD;

    inData811 = 8'h01;
    #CLK_PERIOD;

    inData811 = 8'h02;
    #CLK_PERIOD;

    inData811 = 8'h03;
    #CLK_PERIOD;

    inData811 = 8'h04;
    #CLK_PERIOD;

    inData811 = 8'h05;
    #CLK_PERIOD;

    inData811 = 8'h06;
    #CLK_PERIOD;

    inData811 = 8'h07;
    #CLK_PERIOD;

    inData811 = 8'h08;
    #CLK_PERIOD;

    inData811 = 8'h09;
    #CLK_PERIOD;

    inData811 = 8'h0A;
    #CLK_PERIOD;

    inData811 = 8'h0B;
    #CLK_PERIOD;

    inData811 = 8'h0C;
    #CLK_PERIOD;

    inData811 = 8'h0D;
    #CLK_PERIOD;

    inData811 = 8'h0E;
    #CLK_PERIOD;

    inData811 = 8'h0F;
    #CLK_PERIOD;

    inData811 = 8'h00;
    #CLK_PERIOD;

    inData811 = 8'h10;
    #CLK_PERIOD;

    inData811 = 8'h20;
    #CLK_PERIOD;

    inData811 = 8'h30;
    #CLK_PERIOD;

    inData811 = 8'h40;
    #CLK_PERIOD;

    inData811 = 8'h50;
    #CLK_PERIOD;

    inData811 = 8'h60;
    #CLK_PERIOD;

    inData811 = 8'h70;
    #CLK_PERIOD;

    inData811 = 8'h80;
    #CLK_PERIOD;

    inData811 = 8'h90;
    #CLK_PERIOD;

    inData811 = 8'hA0;
    #CLK_PERIOD;

    inData811 = 8'hB0;
    #CLK_PERIOD;

    inData811 = 8'hC0;
    #CLK_PERIOD;

    inData811 = 8'hD0;
    #CLK_PERIOD;

    inData811 = 8'hE0;
    #CLK_PERIOD;

    inData811 = 8'hF0;
    #CLK_PERIOD;

end



endmodule

