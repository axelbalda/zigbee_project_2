
module MSK_MODULATOR ( clk, reset, i_empty, i_data, o_ready, o_sinI, o_sinQ, 
        o_sinI_four, o_sinQ_four );
  output [3:0] o_sinI;
  output [3:0] o_sinQ;
  output [3:0] o_sinI_four;
  output [3:0] o_sinQ_four;
  input clk, reset, i_empty, i_data;
  output o_ready;
  wire   clk_10M, N459, N460, N461, N462, N463, N464, N465, N466, N467, N468,
         N469, N470, N471, N472, N473, N474, N475, N476, \stateI[0] ,
         \stateQ[0] , IorQ, sin_was_positiveI, sin_was_positiveQ, isPositiveI,
         isPositiveQ, is9, old_i_data, N499, N501, N503, N504, N505, N506,
         N507, N508, N509, N510, N511, N512, N513, N514, N515, N516, N517,
         N518, N519, N520, N521, N522, N564, N651, N652, N655, N695, N696,
         N697, N698, N699, N700, N701, N702, N703, N704, N705, N706, N707,
         N708, N709, N710, N711, N712, N771, N772, N773, N774, N775, N776,
         N777, N778, N779, N780, N781, N782, N783, N784, N785, N786, N787,
         N788, N789, N790, N791, N793, N794, N795, N796, N797, N798, N799,
         N800, N936, N937, N942, N982, N983, N984, N985, N986, N987, N988,
         N989, N990, N991, N992, N993, N994, N995, N996, N997, N998, N999,
         N1059, N1060, N1061, N1062, N1063, N1064, N1065, N1066, N1067, N1068,
         N1069, N1070, N1071, N1072, N1073, N1074, N1075, N1076, N1077, N1078,
         N1079, N1081, N1082, N1083, N1084, N1085, N1086, N1087, N1088, N1090,
         N1091, N1092, N1093, N1094, N1095, N1102, N1103, N1108, N1109, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n191, n192, n193, n194, n195, n196, n197,
         n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208,
         n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, \o_sinQ_four[0] , n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414;
  wire   [19:0] c;
  wire   [19:0] i;
  wire   [19:0] j;
  wire   [19:2] \add_271/carry ;
  wire   [19:2] \add_198/carry ;
  wire   [19:2] \add_93/carry ;
  assign o_sinI_four[0] = \o_sinQ_four[0] ;
  assign o_sinQ_four[0] = \o_sinQ_four[0] ;

  OAI222 U13 ( .A(n129), .B(n130), .C(isPositiveQ), .D(n320), .Q(N937) );
  OAI222 U14 ( .A(n129), .B(n130), .C(n320), .D(n258), .Q(N936) );
  OAI222 U18 ( .A(n292), .B(n276), .C(n137), .D(n138), .Q(N797) );
  OAI222 U20 ( .A(n141), .B(n276), .C(n142), .D(n143), .Q(N796) );
  OAI222 U22 ( .A(n146), .B(n147), .C(n148), .D(n149), .Q(n145) );
  OAI222 U23 ( .A(n150), .B(n347), .C(n350), .D(n143), .Q(n144) );
  OAI222 U26 ( .A(n151), .B(n276), .C(n142), .D(n372), .Q(N795) );
  OAI222 U30 ( .A(n156), .B(n147), .C(n157), .D(n149), .Q(n153) );
  OAI222 U31 ( .A(n156), .B(n138), .C(n157), .D(n158), .Q(n152) );
  OAI212 U40 ( .A(n150), .B(n347), .C(n147), .Q(n140) );
  OAI212 U44 ( .A(n276), .B(n347), .C(n169), .Q(N793) );
  OAI222 U75 ( .A(isPositiveI), .B(n175), .C(n349), .D(n150), .Q(N652) );
  OAI222 U76 ( .A(n175), .B(n259), .C(n349), .D(n150), .Q(N651) );
  OAI212 U118 ( .A(n256), .B(n313), .C(n314), .Q(N1095) );
  OAI222 U139 ( .A(n290), .B(n316), .C(n201), .D(n205), .Q(N1086) );
  OAI212 U140 ( .A(n202), .B(n207), .C(n208), .Q(N1085) );
  OAI212 U141 ( .A(n209), .B(n210), .C(n202), .Q(n208) );
  OAI222 U142 ( .A(n343), .B(n211), .C(n342), .D(n212), .Q(n210) );
  OAI222 U143 ( .A(n214), .B(n207), .C(n130), .D(n215), .Q(n209) );
  OAI222 U146 ( .A(n202), .B(n340), .C(n217), .D(n316), .Q(N1084) );
  OAI222 U149 ( .A(n341), .B(n211), .C(n221), .D(n212), .Q(n219) );
  OAI222 U150 ( .A(n341), .B(n205), .C(n221), .D(n222), .Q(n218) );
  OAI212 U159 ( .A(n130), .B(n215), .C(n211), .Q(n206) );
  OAI212 U167 ( .A(n382), .B(n381), .C(n132), .Q(n234) );
  OAI212 U173 ( .A(n201), .B(n313), .C(n314), .Q(N1081) );
  ADD22 \add_271/U1_1_1  ( .A(j[1]), .B(n270), .CO(\add_271/carry [2]), .S(
        N982) );
  ADD22 \add_271/U1_1_2  ( .A(j[2]), .B(\add_271/carry [2]), .CO(
        \add_271/carry [3]), .S(N983) );
  ADD22 \add_271/U1_1_3  ( .A(j[3]), .B(\add_271/carry [3]), .CO(
        \add_271/carry [4]), .S(N984) );
  ADD22 \add_271/U1_1_4  ( .A(j[4]), .B(\add_271/carry [4]), .CO(
        \add_271/carry [5]), .S(N985) );
  ADD22 \add_271/U1_1_5  ( .A(j[5]), .B(\add_271/carry [5]), .CO(
        \add_271/carry [6]), .S(N986) );
  ADD22 \add_271/U1_1_6  ( .A(j[6]), .B(\add_271/carry [6]), .CO(
        \add_271/carry [7]), .S(N987) );
  ADD22 \add_271/U1_1_7  ( .A(j[7]), .B(\add_271/carry [7]), .CO(
        \add_271/carry [8]), .S(N988) );
  ADD22 \add_271/U1_1_8  ( .A(j[8]), .B(\add_271/carry [8]), .CO(
        \add_271/carry [9]), .S(N989) );
  ADD22 \add_271/U1_1_9  ( .A(j[9]), .B(\add_271/carry [9]), .CO(
        \add_271/carry [10]), .S(N990) );
  ADD22 \add_271/U1_1_10  ( .A(j[10]), .B(\add_271/carry [10]), .CO(
        \add_271/carry [11]), .S(N991) );
  ADD22 \add_271/U1_1_11  ( .A(j[11]), .B(\add_271/carry [11]), .CO(
        \add_271/carry [12]), .S(N992) );
  ADD22 \add_271/U1_1_12  ( .A(j[12]), .B(\add_271/carry [12]), .CO(
        \add_271/carry [13]), .S(N993) );
  ADD22 \add_271/U1_1_13  ( .A(j[13]), .B(\add_271/carry [13]), .CO(
        \add_271/carry [14]), .S(N994) );
  ADD22 \add_271/U1_1_14  ( .A(j[14]), .B(\add_271/carry [14]), .CO(
        \add_271/carry [15]), .S(N995) );
  ADD22 \add_271/U1_1_15  ( .A(j[15]), .B(\add_271/carry [15]), .CO(
        \add_271/carry [16]), .S(N996) );
  ADD22 \add_271/U1_1_16  ( .A(j[16]), .B(\add_271/carry [16]), .CO(
        \add_271/carry [17]), .S(N997) );
  ADD22 \add_271/U1_1_17  ( .A(j[17]), .B(\add_271/carry [17]), .CO(
        \add_271/carry [18]), .S(N998) );
  ADD22 \add_271/U1_1_18  ( .A(j[18]), .B(\add_271/carry [18]), .CO(
        \add_271/carry [19]), .S(N999) );
  ADD22 \add_198/U1_1_1  ( .A(n268), .B(n269), .CO(\add_198/carry [2]), .S(
        N695) );
  ADD22 \add_198/U1_1_2  ( .A(i[2]), .B(\add_198/carry [2]), .CO(
        \add_198/carry [3]), .S(N696) );
  ADD22 \add_198/U1_1_3  ( .A(i[3]), .B(\add_198/carry [3]), .CO(
        \add_198/carry [4]), .S(N697) );
  ADD22 \add_198/U1_1_4  ( .A(i[4]), .B(\add_198/carry [4]), .CO(
        \add_198/carry [5]), .S(N698) );
  ADD22 \add_198/U1_1_5  ( .A(i[5]), .B(\add_198/carry [5]), .CO(
        \add_198/carry [6]), .S(N699) );
  ADD22 \add_198/U1_1_6  ( .A(i[6]), .B(\add_198/carry [6]), .CO(
        \add_198/carry [7]), .S(N700) );
  ADD22 \add_198/U1_1_7  ( .A(i[7]), .B(\add_198/carry [7]), .CO(
        \add_198/carry [8]), .S(N701) );
  ADD22 \add_198/U1_1_8  ( .A(i[8]), .B(\add_198/carry [8]), .CO(
        \add_198/carry [9]), .S(N702) );
  ADD22 \add_198/U1_1_9  ( .A(i[9]), .B(\add_198/carry [9]), .CO(
        \add_198/carry [10]), .S(N703) );
  ADD22 \add_198/U1_1_10  ( .A(i[10]), .B(\add_198/carry [10]), .CO(
        \add_198/carry [11]), .S(N704) );
  ADD22 \add_198/U1_1_11  ( .A(i[11]), .B(\add_198/carry [11]), .CO(
        \add_198/carry [12]), .S(N705) );
  ADD22 \add_198/U1_1_12  ( .A(i[12]), .B(\add_198/carry [12]), .CO(
        \add_198/carry [13]), .S(N706) );
  ADD22 \add_198/U1_1_13  ( .A(i[13]), .B(\add_198/carry [13]), .CO(
        \add_198/carry [14]), .S(N707) );
  ADD22 \add_198/U1_1_14  ( .A(i[14]), .B(\add_198/carry [14]), .CO(
        \add_198/carry [15]), .S(N708) );
  ADD22 \add_198/U1_1_15  ( .A(i[15]), .B(\add_198/carry [15]), .CO(
        \add_198/carry [16]), .S(N709) );
  ADD22 \add_198/U1_1_16  ( .A(i[16]), .B(\add_198/carry [16]), .CO(
        \add_198/carry [17]), .S(N710) );
  ADD22 \add_198/U1_1_17  ( .A(i[17]), .B(\add_198/carry [17]), .CO(
        \add_198/carry [18]), .S(N711) );
  ADD22 \add_198/U1_1_18  ( .A(i[18]), .B(\add_198/carry [18]), .CO(
        \add_198/carry [19]), .S(N712) );
  ADD22 \add_93/U1_1_1  ( .A(c[1]), .B(c[0]), .CO(\add_93/carry [2]), .S(N459)
         );
  ADD22 \add_93/U1_1_2  ( .A(c[2]), .B(\add_93/carry [2]), .CO(
        \add_93/carry [3]), .S(N460) );
  ADD22 \add_93/U1_1_3  ( .A(c[3]), .B(\add_93/carry [3]), .CO(
        \add_93/carry [4]), .S(N461) );
  ADD22 \add_93/U1_1_4  ( .A(c[4]), .B(\add_93/carry [4]), .CO(
        \add_93/carry [5]), .S(N462) );
  ADD22 \add_93/U1_1_5  ( .A(c[5]), .B(\add_93/carry [5]), .CO(
        \add_93/carry [6]), .S(N463) );
  ADD22 \add_93/U1_1_6  ( .A(c[6]), .B(\add_93/carry [6]), .CO(
        \add_93/carry [7]), .S(N464) );
  ADD22 \add_93/U1_1_7  ( .A(c[7]), .B(\add_93/carry [7]), .CO(
        \add_93/carry [8]), .S(N465) );
  ADD22 \add_93/U1_1_8  ( .A(c[8]), .B(\add_93/carry [8]), .CO(
        \add_93/carry [9]), .S(N466) );
  ADD22 \add_93/U1_1_9  ( .A(c[9]), .B(\add_93/carry [9]), .CO(
        \add_93/carry [10]), .S(N467) );
  ADD22 \add_93/U1_1_10  ( .A(c[10]), .B(\add_93/carry [10]), .CO(
        \add_93/carry [11]), .S(N468) );
  ADD22 \add_93/U1_1_11  ( .A(c[11]), .B(\add_93/carry [11]), .CO(
        \add_93/carry [12]), .S(N469) );
  ADD22 \add_93/U1_1_12  ( .A(c[12]), .B(\add_93/carry [12]), .CO(
        \add_93/carry [13]), .S(N470) );
  ADD22 \add_93/U1_1_13  ( .A(c[13]), .B(\add_93/carry [13]), .CO(
        \add_93/carry [14]), .S(N471) );
  ADD22 \add_93/U1_1_14  ( .A(c[14]), .B(\add_93/carry [14]), .CO(
        \add_93/carry [15]), .S(N472) );
  ADD22 \add_93/U1_1_15  ( .A(c[15]), .B(\add_93/carry [15]), .CO(
        \add_93/carry [16]), .S(N473) );
  ADD22 \add_93/U1_1_16  ( .A(c[16]), .B(\add_93/carry [16]), .CO(
        \add_93/carry [17]), .S(N474) );
  ADD22 \add_93/U1_1_17  ( .A(c[17]), .B(\add_93/carry [17]), .CO(
        \add_93/carry [18]), .S(N475) );
  ADD22 \add_93/U1_1_18  ( .A(c[18]), .B(\add_93/carry [18]), .CO(
        \add_93/carry [19]), .S(N476) );
  DF3 \c_reg[0]  ( .D(N503), .C(clk), .Q(c[0]), .QN(n262) );
  DF3 \c_reg[1]  ( .D(N504), .C(clk), .Q(c[1]) );
  DF3 \c_reg[2]  ( .D(N505), .C(clk), .Q(c[2]) );
  DF3 \c_reg[3]  ( .D(N506), .C(clk), .Q(c[3]) );
  DF3 \c_reg[4]  ( .D(N507), .C(clk), .Q(c[4]) );
  DF3 \c_reg[5]  ( .D(N508), .C(clk), .Q(c[5]) );
  DF3 \c_reg[6]  ( .D(N509), .C(clk), .Q(c[6]) );
  DF3 \c_reg[7]  ( .D(N510), .C(clk), .Q(c[7]) );
  DF3 \c_reg[8]  ( .D(N511), .C(clk), .Q(c[8]) );
  DF3 \c_reg[9]  ( .D(N512), .C(clk), .Q(c[9]) );
  DF3 \c_reg[10]  ( .D(N513), .C(clk), .Q(c[10]) );
  DF3 \c_reg[11]  ( .D(N514), .C(clk), .Q(c[11]) );
  DF3 \c_reg[12]  ( .D(N515), .C(clk), .Q(c[12]) );
  DF3 \c_reg[13]  ( .D(N516), .C(clk), .Q(c[13]) );
  DF3 \c_reg[14]  ( .D(N517), .C(clk), .Q(c[14]) );
  DF3 \c_reg[15]  ( .D(N518), .C(clk), .Q(c[15]) );
  DF3 \c_reg[16]  ( .D(N519), .C(clk), .Q(c[16]) );
  DF3 \c_reg[17]  ( .D(N520), .C(clk), .Q(c[17]) );
  DF3 \c_reg[18]  ( .D(N521), .C(clk), .Q(c[18]) );
  DF3 \c_reg[19]  ( .D(N522), .C(clk), .Q(c[19]) );
  DF3 clk_10M_reg ( .D(n311), .C(clk), .Q(clk_10M) );
  DF3 \stateQ_reg[0]  ( .D(N501), .C(clk), .Q(\stateQ[0] ), .QN(n256) );
  DF3 \stateI_reg[0]  ( .D(N499), .C(clk), .Q(\stateI[0] ), .QN(n260) );
  DFE1 \next_stateQ_reg[0]  ( .D(N1108), .E(N1109), .C(clk), .QN(n264) );
  DFE1 \next_stateI_reg[0]  ( .D(N1102), .E(N1103), .C(clk), .QN(n263) );
  DFE1 sin_was_positiveI_reg ( .D(N564), .E(n283), .C(clk), .Q(
        sin_was_positiveI) );
  DFE1 my_clk_10M_reg ( .D(clk_10M), .E(reset), .C(clk), .QN(n251) );
  DFE1 sin_was_positiveQ_reg ( .D(n287), .E(n284), .C(clk), .Q(
        sin_was_positiveQ) );
  DFE1 old_i_data_reg ( .D(N1091), .E(N1090), .C(clk), .Q(old_i_data) );
  DFE1 is9_reg ( .D(N1095), .E(N1094), .C(clk), .Q(is9) );
  DFE1 isPositiveI_reg ( .D(N800), .E(N799), .C(clk), .Q(isPositiveI), .QN(
        n259) );
  DFE1 \j_reg[16]  ( .D(N1076), .E(N1059), .C(clk), .Q(j[16]) );
  DFE1 \i_reg[16]  ( .D(N788), .E(N771), .C(clk), .Q(i[16]) );
  DFE1 \j_reg[15]  ( .D(N1075), .E(n275), .C(clk), .Q(j[15]) );
  DFE1 \i_reg[15]  ( .D(N787), .E(n282), .C(clk), .Q(i[15]) );
  DFE1 \j_reg[17]  ( .D(N1077), .E(n275), .C(clk), .Q(j[17]) );
  DFE1 \i_reg[17]  ( .D(N789), .E(n282), .C(clk), .Q(i[17]) );
  DFE1 \j_reg[18]  ( .D(N1078), .E(N1059), .C(clk), .Q(j[18]) );
  DFE1 \i_reg[18]  ( .D(N790), .E(N771), .C(clk), .Q(i[18]) );
  DFE1 IorQ_reg ( .D(N1093), .E(N1092), .C(clk), .Q(IorQ), .QN(n261) );
  DFE1 \j_reg[19]  ( .D(N1079), .E(n275), .C(clk), .Q(j[19]) );
  DFE1 \i_reg[19]  ( .D(N791), .E(n282), .C(clk), .Q(i[19]) );
  DFE1 isPositiveQ_reg ( .D(n291), .E(N1088), .C(clk), .Q(isPositiveQ), .QN(
        n258) );
  DFE1 \j_reg[12]  ( .D(N1072), .E(N1059), .C(clk), .Q(j[12]) );
  DFE1 \i_reg[12]  ( .D(N784), .E(N771), .C(clk), .Q(i[12]) );
  DFE1 \j_reg[14]  ( .D(N1074), .E(N1059), .C(clk), .Q(j[14]) );
  DFE1 \i_reg[14]  ( .D(N786), .E(N771), .C(clk), .Q(i[14]) );
  DFE1 \j_reg[13]  ( .D(N1073), .E(n275), .C(clk), .Q(j[13]) );
  DFE1 \i_reg[13]  ( .D(N785), .E(n282), .C(clk), .Q(i[13]) );
  DFE1 \j_reg[10]  ( .D(N1070), .E(N1059), .C(clk), .Q(j[10]) );
  DFE1 \j_reg[11]  ( .D(N1071), .E(n275), .C(clk), .Q(j[11]) );
  DFE1 \i_reg[10]  ( .D(N782), .E(N771), .C(clk), .Q(i[10]) );
  DFE1 \i_reg[11]  ( .D(N783), .E(n282), .C(clk), .Q(i[11]) );
  DFE1 \j_reg[9]  ( .D(N1069), .E(n275), .C(clk), .Q(j[9]) );
  DFE1 \i_reg[9]  ( .D(N781), .E(n282), .C(clk), .Q(i[9]) );
  DFE1 \j_reg[7]  ( .D(N1067), .E(n275), .C(clk), .Q(j[7]) );
  DFE1 \j_reg[8]  ( .D(N1068), .E(N1059), .C(clk), .Q(j[8]) );
  DFE1 \i_reg[7]  ( .D(N779), .E(n282), .C(clk), .Q(i[7]) );
  DFE1 \i_reg[8]  ( .D(N780), .E(N771), .C(clk), .Q(i[8]) );
  DFE1 \j_reg[4]  ( .D(N1064), .E(N1059), .C(clk), .Q(j[4]) );
  DFE1 \j_reg[5]  ( .D(N1065), .E(n275), .C(clk), .Q(j[5]) );
  DFE1 \i_reg[4]  ( .D(N776), .E(N771), .C(clk), .Q(i[4]) );
  DFE1 \i_reg[5]  ( .D(N777), .E(n282), .C(clk), .Q(i[5]) );
  DFE1 \j_reg[6]  ( .D(N1066), .E(N1059), .C(clk), .Q(j[6]) );
  DFE1 \i_reg[6]  ( .D(N778), .E(N771), .C(clk), .Q(i[6]) );
  DFE1 \i_reg[1]  ( .D(N773), .E(n282), .C(clk), .Q(i[1]) );
  DFE1 \j_reg[0]  ( .D(N1060), .E(N1059), .C(clk), .Q(j[0]), .QN(n252) );
  DFE1 \i_reg[3]  ( .D(N775), .E(n282), .C(clk), .Q(i[3]) );
  DFE1 \j_reg[1]  ( .D(N1061), .E(n275), .C(clk), .Q(j[1]), .QN(n250) );
  DFE1 \j_reg[3]  ( .D(N1063), .E(n275), .C(clk), .Q(j[3]), .QN(n255) );
  DFE1 \j_reg[2]  ( .D(N1062), .E(N1059), .C(clk), .Q(j[2]), .QN(n254) );
  DFE1 \i_reg[2]  ( .D(N774), .E(N771), .C(clk), .Q(i[2]), .QN(n257) );
  DFE1 \i_reg[0]  ( .D(N772), .E(N771), .C(clk), .Q(i[0]), .QN(n253) );
  DFE1 \o_sinI_four_reg[3]  ( .D(N652), .E(N798), .C(clk), .Q(o_sinI_four[3])
         );
  DFE1 \o_sinI_reg[0]  ( .D(N794), .E(N793), .C(clk), .Q(o_sinI[0]) );
  DFE1 \o_sinQ_four_reg[3]  ( .D(N937), .E(N1087), .C(clk), .Q(o_sinQ_four[3])
         );
  DFE1 \o_sinQ_reg[0]  ( .D(N1083), .E(N1082), .C(clk), .Q(o_sinQ[0]) );
  DFE1 \o_sinI_four_reg[1]  ( .D(N651), .E(N798), .C(clk), .Q(o_sinI_four[1])
         );
  DFE1 \o_sinI_four_reg[2]  ( .D(N651), .E(N798), .C(clk), .Q(o_sinI_four[2])
         );
  DFE1 \o_sinI_reg[1]  ( .D(N795), .E(N793), .C(clk), .Q(o_sinI[1]) );
  DFE1 \o_sinI_reg[2]  ( .D(N796), .E(N793), .C(clk), .Q(o_sinI[2]) );
  DFE1 \o_sinI_reg[3]  ( .D(N797), .E(N793), .C(clk), .Q(o_sinI[3]) );
  DFE1 \o_sinQ_four_reg[1]  ( .D(N936), .E(N1087), .C(clk), .Q(o_sinQ_four[1])
         );
  DFE1 \o_sinQ_four_reg[2]  ( .D(N936), .E(N1087), .C(clk), .Q(o_sinQ_four[2])
         );
  DFE1 o_ready_reg ( .D(N1081), .E(n286), .C(clk), .Q(o_ready) );
  DFE1 \o_sinQ_reg[2]  ( .D(N1085), .E(N1082), .C(clk), .Q(o_sinQ[2]) );
  DFE1 \o_sinQ_reg[1]  ( .D(N1084), .E(N1082), .C(clk), .Q(o_sinQ[1]) );
  DFE1 \o_sinQ_reg[3]  ( .D(N1086), .E(N1082), .C(clk), .Q(o_sinQ[3]) );
  LOGIC1 U344 ( .Q(\o_sinQ_four[0] ) );
  NOR21 U345 ( .A(n279), .B(n265), .Q(N791) );
  NOR21 U346 ( .A(n272), .B(n266), .Q(N1079) );
  NOR21 U347 ( .A(n177), .B(n267), .Q(N522) );
  INV3 U348 ( .A(n201), .Q(n315) );
  INV3 U349 ( .A(n237), .Q(n313) );
  NOR21 U350 ( .A(n316), .B(n319), .Q(n201) );
  NAND22 U351 ( .A(n142), .B(n350), .Q(n135) );
  INV3 U352 ( .A(n139), .Q(n350) );
  NOR21 U353 ( .A(n188), .B(n276), .Q(n237) );
  NAND22 U354 ( .A(n315), .B(n192), .Q(N1087) );
  NAND22 U355 ( .A(n135), .B(n136), .Q(N798) );
  NAND22 U356 ( .A(n162), .B(n351), .Q(n139) );
  NAND22 U357 ( .A(n317), .B(n214), .Q(n215) );
  INV3 U358 ( .A(n172), .Q(n347) );
  NOR21 U359 ( .A(n170), .B(n139), .Q(n172) );
  INV3 U360 ( .A(n214), .Q(n319) );
  INV3 U361 ( .A(n216), .Q(n342) );
  AOI221 U362 ( .A(n375), .B(n380), .C(n374), .D(n379), .Q(n143) );
  INV3 U363 ( .A(n146), .Q(n375) );
  AOI221 U364 ( .A(n213), .B(n382), .C(n216), .D(n381), .Q(n207) );
  INV3 U365 ( .A(n202), .Q(n316) );
  NAND22 U366 ( .A(n202), .B(n129), .Q(n192) );
  NAND22 U367 ( .A(n279), .B(n174), .Q(N771) );
  NAND22 U368 ( .A(n278), .B(n174), .Q(n282) );
  NAND22 U369 ( .A(n272), .B(n133), .Q(N1059) );
  NAND22 U370 ( .A(n271), .B(n133), .Q(n275) );
  NAND22 U371 ( .A(n349), .B(n142), .Q(n136) );
  NAND22 U372 ( .A(n198), .B(i[3]), .Q(n188) );
  NOR21 U373 ( .A(n352), .B(i[3]), .Q(n196) );
  INV3 U374 ( .A(n198), .Q(n352) );
  INV3 U375 ( .A(n236), .Q(n314) );
  INV3 U376 ( .A(n129), .Q(n320) );
  NOR21 U377 ( .A(n279), .B(n369), .Q(N775) );
  INV3 U378 ( .A(N697), .Q(n369) );
  NOR21 U379 ( .A(n281), .B(n371), .Q(N773) );
  INV3 U380 ( .A(N695), .Q(n371) );
  INV3 U381 ( .A(n213), .Q(n343) );
  INV3 U382 ( .A(n133), .Q(n284) );
  INV3 U383 ( .A(n174), .Q(n283) );
  NOR21 U384 ( .A(n177), .B(n294), .Q(N520) );
  INV3 U385 ( .A(N475), .Q(n294) );
  NOR21 U386 ( .A(n271), .B(n322), .Q(N1078) );
  INV3 U387 ( .A(N999), .Q(n322) );
  NOR21 U388 ( .A(n274), .B(n323), .Q(N1077) );
  INV3 U389 ( .A(N998), .Q(n323) );
  NOR21 U390 ( .A(n273), .B(n324), .Q(N1076) );
  INV3 U391 ( .A(N997), .Q(n324) );
  NOR21 U392 ( .A(n281), .B(n355), .Q(N789) );
  INV3 U393 ( .A(N711), .Q(n355) );
  NOR21 U394 ( .A(n280), .B(n356), .Q(N788) );
  INV3 U395 ( .A(N710), .Q(n356) );
  NOR21 U396 ( .A(n278), .B(n354), .Q(N790) );
  INV3 U397 ( .A(N712), .Q(n354) );
  NOR21 U398 ( .A(n277), .B(n293), .Q(N521) );
  INV3 U399 ( .A(N476), .Q(n293) );
  NOR21 U400 ( .A(n277), .B(n295), .Q(N519) );
  INV3 U401 ( .A(N474), .Q(n295) );
  NOR21 U402 ( .A(n277), .B(n297), .Q(N517) );
  INV3 U403 ( .A(N472), .Q(n297) );
  NOR21 U404 ( .A(n274), .B(n325), .Q(N1075) );
  INV3 U405 ( .A(N996), .Q(n325) );
  NOR21 U406 ( .A(n273), .B(n326), .Q(N1074) );
  INV3 U407 ( .A(N995), .Q(n326) );
  NOR21 U408 ( .A(n280), .B(n358), .Q(N786) );
  INV3 U409 ( .A(N708), .Q(n358) );
  NOR21 U410 ( .A(n281), .B(n357), .Q(N787) );
  INV3 U411 ( .A(N709), .Q(n357) );
  NOR21 U412 ( .A(n279), .B(n359), .Q(N785) );
  INV3 U413 ( .A(N707), .Q(n359) );
  NOR21 U414 ( .A(n177), .B(n296), .Q(N518) );
  INV3 U415 ( .A(N473), .Q(n296) );
  NOR21 U416 ( .A(n177), .B(n298), .Q(N516) );
  INV3 U417 ( .A(N471), .Q(n298) );
  NOR21 U418 ( .A(n272), .B(n327), .Q(N1073) );
  INV3 U419 ( .A(N994), .Q(n327) );
  NOR21 U420 ( .A(n271), .B(n328), .Q(N1072) );
  INV3 U421 ( .A(N993), .Q(n328) );
  NOR21 U422 ( .A(n279), .B(n361), .Q(N783) );
  INV3 U423 ( .A(N705), .Q(n361) );
  NOR21 U424 ( .A(n272), .B(n329), .Q(N1071) );
  INV3 U425 ( .A(N992), .Q(n329) );
  NOR21 U426 ( .A(n278), .B(n360), .Q(N784) );
  INV3 U427 ( .A(N706), .Q(n360) );
  NOR21 U428 ( .A(n277), .B(n299), .Q(N515) );
  INV3 U429 ( .A(N470), .Q(n299) );
  NOR21 U430 ( .A(n177), .B(n302), .Q(N512) );
  INV3 U431 ( .A(N467), .Q(n302) );
  NOR21 U432 ( .A(n271), .B(n330), .Q(N1070) );
  INV3 U433 ( .A(N991), .Q(n330) );
  NOR21 U434 ( .A(n273), .B(n332), .Q(N1068) );
  INV3 U435 ( .A(N989), .Q(n332) );
  NOR21 U436 ( .A(n280), .B(n364), .Q(N780) );
  INV3 U437 ( .A(N702), .Q(n364) );
  NOR21 U438 ( .A(n278), .B(n362), .Q(N782) );
  INV3 U439 ( .A(N704), .Q(n362) );
  NOR21 U440 ( .A(n281), .B(n363), .Q(N781) );
  INV3 U441 ( .A(N703), .Q(n363) );
  NOR21 U442 ( .A(n274), .B(n331), .Q(N1069) );
  INV3 U443 ( .A(N990), .Q(n331) );
  NOR21 U444 ( .A(n177), .B(n300), .Q(N514) );
  INV3 U445 ( .A(N469), .Q(n300) );
  NOR21 U446 ( .A(n277), .B(n301), .Q(N513) );
  INV3 U447 ( .A(N468), .Q(n301) );
  AOI211 U448 ( .A(n142), .B(n170), .C(n171), .Q(n169) );
  AOI211 U449 ( .A(n158), .B(n138), .C(n288), .Q(n171) );
  NAND22 U450 ( .A(n254), .B(n250), .Q(n216) );
  NAND31 U451 ( .A(n252), .B(n255), .C(n342), .Q(n227) );
  NAND22 U452 ( .A(N655), .B(n259), .Q(n147) );
  NAND22 U453 ( .A(N942), .B(n258), .Q(n211) );
  NOR21 U454 ( .A(n227), .B(n203), .Q(n214) );
  NOR21 U455 ( .A(n139), .B(n276), .Q(n137) );
  INV3 U456 ( .A(n140), .Q(n292) );
  NOR21 U457 ( .A(n144), .B(n145), .Q(n141) );
  NAND22 U458 ( .A(n149), .B(n147), .Q(n170) );
  NOR21 U459 ( .A(n277), .B(n303), .Q(N511) );
  INV3 U460 ( .A(N466), .Q(n303) );
  NOR21 U461 ( .A(n177), .B(n304), .Q(N510) );
  INV3 U462 ( .A(N465), .Q(n304) );
  INV3 U463 ( .A(n239), .Q(n351) );
  NAND22 U464 ( .A(n149), .B(n347), .Q(n167) );
  NOR21 U465 ( .A(n272), .B(n335), .Q(N1065) );
  INV3 U466 ( .A(N986), .Q(n335) );
  NOR21 U467 ( .A(n279), .B(n367), .Q(N777) );
  INV3 U468 ( .A(N699), .Q(n367) );
  NOR21 U469 ( .A(n274), .B(n333), .Q(N1067) );
  INV3 U470 ( .A(N988), .Q(n333) );
  NOR21 U471 ( .A(n273), .B(n334), .Q(N1066) );
  INV3 U472 ( .A(N987), .Q(n334) );
  INV3 U473 ( .A(n235), .Q(n317) );
  NAND22 U474 ( .A(n212), .B(n211), .Q(n235) );
  NOR21 U475 ( .A(n281), .B(n365), .Q(N779) );
  INV3 U476 ( .A(N701), .Q(n365) );
  INV3 U477 ( .A(n238), .Q(n286) );
  NOR40 U478 ( .A(n201), .B(n236), .C(n237), .D(N799), .Q(n238) );
  NOR21 U479 ( .A(n280), .B(n366), .Q(N778) );
  INV3 U480 ( .A(N700), .Q(n366) );
  NOR21 U481 ( .A(n277), .B(n305), .Q(N509) );
  INV3 U482 ( .A(N464), .Q(n305) );
  OAI2111 U483 ( .A(n317), .B(n316), .C(n315), .D(n234), .Q(N1082) );
  NOR21 U484 ( .A(n256), .B(n251), .Q(n202) );
  NOR31 U485 ( .A(n254), .B(n203), .C(n204), .Q(n129) );
  NAND31 U486 ( .A(n252), .B(n255), .C(n250), .Q(n204) );
  AOI2111 U487 ( .A(n253), .B(i[3]), .C(n159), .D(n373), .Q(n157) );
  AOI211 U488 ( .A(n269), .B(n268), .C(n257), .Q(n159) );
  INV3 U489 ( .A(n160), .Q(n373) );
  AOI311 U490 ( .A(n269), .B(n257), .C(n268), .D(n161), .Q(n160) );
  AOI2111 U491 ( .A(n269), .B(i[3]), .C(n162), .D(n268), .Q(n156) );
  NOR31 U492 ( .A(n216), .B(n203), .C(n252), .Q(n199) );
  INV3 U493 ( .A(n206), .Q(n290) );
  INV3 U494 ( .A(n218), .Q(n340) );
  AOI2111 U495 ( .A(n218), .B(n319), .C(n219), .D(n220), .Q(n217) );
  NOR31 U496 ( .A(n239), .B(n374), .C(n253), .Q(n198) );
  INV3 U497 ( .A(n152), .Q(n372) );
  AOI2111 U498 ( .A(n152), .B(n139), .C(n153), .D(n154), .Q(n151) );
  NOR31 U499 ( .A(n269), .B(i[3]), .C(n374), .Q(n162) );
  NOR21 U500 ( .A(n316), .B(n187), .Q(n236) );
  NAND22 U501 ( .A(n199), .B(n255), .Q(n194) );
  NOR21 U502 ( .A(n130), .B(n215), .Q(n220) );
  NAND22 U503 ( .A(n216), .B(n255), .Q(n213) );
  NOR21 U504 ( .A(n148), .B(i[3]), .Q(n146) );
  INV3 U505 ( .A(n148), .Q(n374) );
  BUF2 U506 ( .A(n248), .Q(n271) );
  BUF2 U507 ( .A(n248), .Q(n272) );
  BUF2 U508 ( .A(n173), .Q(n278) );
  BUF2 U509 ( .A(n173), .Q(n279) );
  NOR31 U510 ( .A(n253), .B(i[3]), .C(n268), .Q(n161) );
  NOR21 U511 ( .A(n177), .B(n306), .Q(N508) );
  INV3 U512 ( .A(N463), .Q(n306) );
  NOR21 U513 ( .A(n277), .B(n307), .Q(N507) );
  INV3 U514 ( .A(N462), .Q(n307) );
  NOR21 U515 ( .A(n177), .B(n308), .Q(N506) );
  INV3 U516 ( .A(N461), .Q(n308) );
  NOR21 U517 ( .A(n277), .B(n309), .Q(N505) );
  INV3 U518 ( .A(N460), .Q(n309) );
  NOR21 U519 ( .A(n177), .B(n310), .Q(N504) );
  INV3 U520 ( .A(N459), .Q(n310) );
  INV3 U521 ( .A(n175), .Q(n349) );
  BUF2 U522 ( .A(n248), .Q(n274) );
  BUF2 U523 ( .A(n248), .Q(n273) );
  BUF2 U524 ( .A(n173), .Q(n281) );
  BUF2 U525 ( .A(n173), .Q(n280) );
  INV3 U526 ( .A(n222), .Q(n381) );
  INV3 U527 ( .A(n205), .Q(n382) );
  INV3 U528 ( .A(n176), .Q(n288) );
  NOR21 U529 ( .A(n150), .B(n347), .Q(n154) );
  INV3 U530 ( .A(n142), .Q(n276) );
  NOR21 U531 ( .A(n251), .B(n260), .Q(n142) );
  NAND22 U532 ( .A(n212), .B(n215), .Q(n232) );
  NOR21 U533 ( .A(n134), .B(n135), .Q(N800) );
  INV3 U534 ( .A(n138), .Q(n380) );
  INV3 U535 ( .A(n226), .Q(n341) );
  OAI2111 U536 ( .A(n252), .B(n255), .C(n227), .D(n250), .Q(n226) );
  NOR21 U537 ( .A(n271), .B(n336), .Q(N1064) );
  INV3 U538 ( .A(N985), .Q(n336) );
  NOR21 U539 ( .A(n272), .B(n337), .Q(N1063) );
  INV3 U540 ( .A(N984), .Q(n337) );
  NOR21 U541 ( .A(n271), .B(n338), .Q(N1062) );
  INV3 U542 ( .A(N983), .Q(n338) );
  NOR21 U543 ( .A(n278), .B(n368), .Q(N776) );
  INV3 U544 ( .A(N698), .Q(n368) );
  NOR21 U545 ( .A(n278), .B(n370), .Q(N774) );
  INV3 U546 ( .A(N696), .Q(n370) );
  NOR21 U547 ( .A(n274), .B(n339), .Q(N1061) );
  INV3 U548 ( .A(N982), .Q(n339) );
  INV3 U549 ( .A(n200), .Q(n291) );
  NAND22 U550 ( .A(n130), .B(n201), .Q(n200) );
  NOR21 U551 ( .A(n285), .B(n132), .Q(n133) );
  NOR21 U552 ( .A(n285), .B(n176), .Q(n174) );
  INV3 U553 ( .A(n158), .Q(n379) );
  NOR21 U554 ( .A(n259), .B(n288), .Q(N564) );
  INV3 U555 ( .A(n128), .Q(n311) );
  BUF2 U556 ( .A(i[0]), .Q(n269) );
  XNR21 U557 ( .A(\add_198/carry [19]), .B(i[19]), .Q(n265) );
  BUF2 U558 ( .A(i[1]), .Q(n268) );
  BUF2 U559 ( .A(j[0]), .Q(n270) );
  XNR21 U560 ( .A(\add_271/carry [19]), .B(j[19]), .Q(n266) );
  XNR21 U561 ( .A(\add_93/carry [19]), .B(c[19]), .Q(n267) );
  NAND41 U562 ( .A(n240), .B(n241), .C(n242), .D(n243), .Q(n239) );
  NOR40 U563 ( .A(i[9]), .B(i[8]), .C(i[7]), .D(i[6]), .Q(n243) );
  NOR40 U564 ( .A(i[5]), .B(i[4]), .C(i[19]), .D(i[18]), .Q(n242) );
  NOR40 U565 ( .A(i[17]), .B(i[16]), .C(i[15]), .D(i[14]), .Q(n241) );
  NAND41 U566 ( .A(n400), .B(n399), .C(n398), .D(n397), .Q(N942) );
  NOR31 U567 ( .A(j[11]), .B(j[13]), .C(j[12]), .Q(n399) );
  NOR21 U568 ( .A(j[10]), .B(n270), .Q(n400) );
  NOR40 U569 ( .A(j[16]), .B(n346), .C(j[15]), .D(j[14]), .Q(n398) );
  NAND41 U570 ( .A(n391), .B(n390), .C(n389), .D(n388), .Q(N655) );
  NOR31 U571 ( .A(i[11]), .B(i[13]), .C(i[12]), .Q(n390) );
  NOR21 U572 ( .A(i[10]), .B(n269), .Q(n391) );
  NOR40 U573 ( .A(i[16]), .B(n378), .C(i[15]), .D(i[14]), .Q(n389) );
  NOR40 U574 ( .A(i[13]), .B(i[12]), .C(i[11]), .D(i[10]), .Q(n240) );
  NAND22 U575 ( .A(N942), .B(isPositiveQ), .Q(n212) );
  NAND22 U576 ( .A(N655), .B(isPositiveI), .Q(n149) );
  NOR40 U577 ( .A(n396), .B(n344), .C(j[1]), .D(j[19]), .Q(n397) );
  NAND22 U578 ( .A(n394), .B(n393), .Q(n396) );
  INV3 U579 ( .A(n395), .Q(n344) );
  NOR21 U580 ( .A(j[6]), .B(j[5]), .Q(n394) );
  NOR40 U581 ( .A(n387), .B(n376), .C(n268), .D(i[19]), .Q(n388) );
  NAND22 U582 ( .A(n385), .B(n384), .Q(n387) );
  INV3 U583 ( .A(n386), .Q(n376) );
  NOR21 U584 ( .A(i[6]), .B(i[5]), .Q(n385) );
  OAI311 U585 ( .A(n251), .B(n163), .C(n260), .D(n165), .Q(N794) );
  AOI221 U586 ( .A(n380), .B(n166), .C(n379), .D(n166), .Q(n165) );
  AOI221 U587 ( .A(n167), .B(n166), .C(n166), .D(n140), .Q(n163) );
  OAI2111 U588 ( .A(n269), .B(i[2]), .C(n268), .D(n168), .Q(n166) );
  OAI311 U589 ( .A(n256), .B(n229), .C(n251), .D(n230), .Q(N1083) );
  AOI221 U590 ( .A(n382), .B(n231), .C(n381), .D(n231), .Q(n230) );
  AOI221 U591 ( .A(n232), .B(n231), .C(n231), .D(n206), .Q(n229) );
  OAI2111 U592 ( .A(n270), .B(j[2]), .C(j[1]), .D(n233), .Q(n231) );
  NOR31 U593 ( .A(i[2]), .B(i[4]), .C(i[3]), .Q(n386) );
  NOR31 U594 ( .A(j[2]), .B(j[4]), .C(j[3]), .Q(n395) );
  NOR31 U595 ( .A(j[7]), .B(j[9]), .C(j[8]), .Q(n393) );
  NOR31 U596 ( .A(i[7]), .B(i[9]), .C(i[8]), .Q(n384) );
  NAND22 U597 ( .A(reset), .B(n135), .Q(N799) );
  XOR21 U598 ( .A(sin_was_positiveQ), .B(n155), .Q(n130) );
  NAND22 U599 ( .A(reset), .B(n128), .Q(n177) );
  NAND22 U600 ( .A(reset), .B(n128), .Q(n277) );
  NAND41 U601 ( .A(n178), .B(n179), .C(n180), .D(n181), .Q(n128) );
  NOR21 U602 ( .A(c[14]), .B(c[13]), .Q(n178) );
  NOR31 U603 ( .A(c[15]), .B(c[17]), .C(c[16]), .Q(n179) );
  NOR40 U604 ( .A(n186), .B(c[10]), .C(c[12]), .D(c[11]), .Q(n180) );
  NAND41 U605 ( .A(n244), .B(n245), .C(n246), .D(n247), .Q(n203) );
  NOR40 U606 ( .A(j[9]), .B(j[8]), .C(j[7]), .D(j[6]), .Q(n247) );
  NOR40 U607 ( .A(j[5]), .B(j[4]), .C(j[19]), .D(j[18]), .Q(n246) );
  NOR40 U608 ( .A(j[17]), .B(j[16]), .C(j[15]), .D(j[14]), .Q(n245) );
  XNR21 U609 ( .A(old_i_data), .B(i_data), .Q(n155) );
  XNR21 U610 ( .A(sin_was_positiveI), .B(n155), .Q(n134) );
  NAND31 U611 ( .A(i[2]), .B(n351), .C(n193), .Q(n175) );
  NOR31 U612 ( .A(n269), .B(i[3]), .C(n268), .Q(n193) );
  NOR40 U613 ( .A(j[13]), .B(j[12]), .C(j[11]), .D(j[10]), .Q(n244) );
  NOR40 U614 ( .A(i[12]), .B(i[11]), .C(i[10]), .D(n353), .Q(n406) );
  INV3 U615 ( .A(n401), .Q(n353) );
  OAI311 U616 ( .A(n269), .B(i[2]), .C(n268), .D(i[3]), .Q(n401) );
  NOR40 U617 ( .A(j[12]), .B(j[11]), .C(j[10]), .D(n321), .Q(n413) );
  INV3 U618 ( .A(n408), .Q(n321) );
  OAI311 U619 ( .A(n270), .B(j[2]), .C(j[1]), .D(j[3]), .Q(n408) );
  XOR21 U620 ( .A(sin_was_positiveI), .B(n155), .Q(n150) );
  NAND22 U621 ( .A(isPositiveI), .B(is9), .Q(n158) );
  NOR40 U622 ( .A(i[16]), .B(i[15]), .C(i[14]), .D(i[13]), .Q(n405) );
  NOR40 U623 ( .A(j[16]), .B(j[15]), .C(j[14]), .D(j[13]), .Q(n412) );
  NAND22 U624 ( .A(is9), .B(n158), .Q(n138) );
  NOR40 U625 ( .A(i[7]), .B(n377), .C(i[6]), .D(i[5]), .Q(n403) );
  INV3 U626 ( .A(n402), .Q(n377) );
  NOR21 U627 ( .A(i[9]), .B(i[8]), .Q(n402) );
  NOR40 U628 ( .A(j[7]), .B(n345), .C(j[6]), .D(j[5]), .Q(n410) );
  INV3 U629 ( .A(n409), .Q(n345) );
  NOR21 U630 ( .A(j[9]), .B(j[8]), .Q(n409) );
  NOR31 U631 ( .A(\stateI[0] ), .B(i_empty), .C(n261), .Q(n176) );
  NAND41 U632 ( .A(n314), .B(n313), .C(\stateQ[0] ), .D(n191), .Q(N1094) );
  NOR21 U633 ( .A(n260), .B(n285), .Q(n191) );
  AOI2111 U634 ( .A(n252), .B(j[3]), .C(n223), .D(n224), .Q(n221) );
  AOI211 U635 ( .A(n270), .B(j[1]), .C(n254), .Q(n223) );
  OAI311 U636 ( .A(n252), .B(j[2]), .C(n250), .D(n225), .Q(n224) );
  NAND31 U637 ( .A(n270), .B(n255), .C(n250), .Q(n225) );
  OAI2111 U638 ( .A(n316), .B(n194), .C(n197), .D(reset), .Q(N1090) );
  NAND22 U639 ( .A(n196), .B(n142), .Q(n197) );
  NAND22 U640 ( .A(is9), .B(isPositiveQ), .Q(n222) );
  NOR21 U641 ( .A(i[2]), .B(n268), .Q(n148) );
  NOR40 U642 ( .A(n182), .B(n312), .C(c[19]), .D(c[18]), .Q(n181) );
  INV3 U643 ( .A(n183), .Q(n312) );
  NAND22 U644 ( .A(n184), .B(n185), .Q(n182) );
  NOR31 U645 ( .A(c[1]), .B(c[4]), .C(c[3]), .Q(n183) );
  NAND22 U646 ( .A(is9), .B(n222), .Q(n205) );
  AOI211 U647 ( .A(i[2]), .B(n269), .C(i[3]), .Q(n168) );
  AOI211 U648 ( .A(j[2]), .B(n270), .C(j[3]), .Q(n233) );
  NAND22 U649 ( .A(j[3]), .B(n199), .Q(n187) );
  OAI311 U650 ( .A(n194), .B(n289), .C(n316), .D(n195), .Q(N1091) );
  INV3 U651 ( .A(i_data), .Q(n289) );
  NAND31 U652 ( .A(n142), .B(i_data), .C(n196), .Q(n195) );
  NOR31 U653 ( .A(c[7]), .B(c[9]), .C(c[8]), .Q(n185) );
  NAND31 U654 ( .A(n136), .B(n192), .C(reset), .Q(N1092) );
  NAND22 U655 ( .A(n318), .B(n202), .Q(n248) );
  INV3 U656 ( .A(n414), .Q(n318) );
  NAND41 U657 ( .A(n413), .B(n412), .C(n411), .D(n410), .Q(n414) );
  NOR40 U658 ( .A(j[4]), .B(j[19]), .C(j[18]), .D(j[17]), .Q(n411) );
  AOI211 U659 ( .A(n136), .B(n192), .C(IorQ), .Q(N1093) );
  NAND22 U660 ( .A(n348), .B(n142), .Q(n173) );
  INV3 U661 ( .A(n407), .Q(n348) );
  NAND41 U662 ( .A(n406), .B(n405), .C(n404), .D(n403), .Q(n407) );
  NOR40 U663 ( .A(i[4]), .B(i[19]), .C(i[18]), .D(i[17]), .Q(n404) );
  NOR21 U664 ( .A(n277), .B(c[0]), .Q(N503) );
  NAND22 U665 ( .A(c[2]), .B(n262), .Q(n186) );
  NAND22 U666 ( .A(reset), .B(n315), .Q(N1088) );
  NOR21 U667 ( .A(n273), .B(n270), .Q(N1060) );
  NOR21 U668 ( .A(n280), .B(n269), .Q(N772) );
  INV3 U669 ( .A(n392), .Q(n346) );
  NOR21 U670 ( .A(j[18]), .B(j[17]), .Q(n392) );
  INV3 U671 ( .A(n383), .Q(n378) );
  NOR21 U672 ( .A(i[18]), .B(i[17]), .Q(n383) );
  NOR31 U673 ( .A(IorQ), .B(i_empty), .C(\stateQ[0] ), .Q(n132) );
  NOR31 U674 ( .A(IorQ), .B(\stateQ[0] ), .C(i_empty), .Q(N1108) );
  NOR31 U675 ( .A(n261), .B(\stateI[0] ), .C(i_empty), .Q(N1102) );
  NOR21 U676 ( .A(c[6]), .B(c[5]), .Q(n184) );
  INV3 U677 ( .A(n131), .Q(n287) );
  NAND22 U678 ( .A(isPositiveQ), .B(n132), .Q(n131) );
  NOR21 U679 ( .A(n263), .B(n285), .Q(N499) );
  NOR21 U680 ( .A(n264), .B(n285), .Q(N501) );
  INV3 U681 ( .A(reset), .Q(n285) );
  OAI212 U682 ( .A(n187), .B(n251), .C(\stateQ[0] ), .Q(N1109) );
  OAI212 U683 ( .A(n188), .B(n251), .C(\stateI[0] ), .Q(N1103) );
endmodule

