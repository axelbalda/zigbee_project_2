
module TOP ( inClock, inReset, in_inFIFO_inData, in_outFIFO_inReadEnable, 
        in_DEMUX_inDEMUX1, in_DEMUX_inDEMUX2, in_DEMUX_inDEMUX17, 
        in_DEMUX_inDEMUX18, in_DEMUX_inSEL1, in_DEMUX_inSEL2, in_MUX_inSEL3, 
        in_MUX_inSEL6, in_MUX_inSEL9, in_MUX_inSEL11, in_MUX_inSEL12, 
        in_MUX_inSEL15, in_DEMUX_inSEL17, out_MUX_outMUX9, out_MUX_outMUX10, 
        out_MUX_outMUX15, out_MUX_outMUX16 );
  input [3:0] in_inFIFO_inData;
  input [3:0] in_DEMUX_inDEMUX17;
  input [3:0] in_DEMUX_inDEMUX18;
  input [2:0] in_DEMUX_inSEL1;
  input [2:0] in_DEMUX_inSEL2;
  input [1:0] in_MUX_inSEL6;
  input [1:0] in_MUX_inSEL9;
  input [1:0] in_MUX_inSEL15;
  output [3:0] out_MUX_outMUX9;
  output [3:0] out_MUX_outMUX10;
  input inClock, inReset, in_outFIFO_inReadEnable, in_DEMUX_inDEMUX1,
         in_DEMUX_inDEMUX2, in_MUX_inSEL3, in_MUX_inSEL11, in_MUX_inSEL12,
         in_DEMUX_inSEL17;
  output out_MUX_outMUX15, out_MUX_outMUX16;
  wire   \sig_MUX_inMUX3[0] , \sig_MUX_inMUX4[0] , \sig_MUX_inMUX5[0] ,
         \sig_MUX_inMUX8[0] , sig_MUX_outMUX8, \sig_MUX_inMUX11[0] ,
         \sig_MUX_inMUX14[0] , \sig_MUX_inMUX12[0] , \sig_MUX_inMUX13[0] ,
         \u_inFIFO/n294 , \u_inFIFO/n293 , \u_inFIFO/n292 , \u_inFIFO/n291 ,
         \u_inFIFO/n290 , \u_inFIFO/n289 , \u_inFIFO/n288 , \u_inFIFO/n287 ,
         \u_inFIFO/n286 , \u_inFIFO/n285 , \u_inFIFO/n284 , \u_inFIFO/n283 ,
         \u_inFIFO/n282 , \u_inFIFO/n281 , \u_inFIFO/n280 , \u_inFIFO/n279 ,
         \u_inFIFO/n278 , \u_inFIFO/n277 , \u_inFIFO/n276 , \u_inFIFO/n275 ,
         \u_inFIFO/n274 , \u_inFIFO/n273 , \u_inFIFO/n272 , \u_inFIFO/n271 ,
         \u_inFIFO/n270 , \u_inFIFO/n269 , \u_inFIFO/n268 , \u_inFIFO/n267 ,
         \u_inFIFO/n266 , \u_inFIFO/n265 , \u_inFIFO/n264 , \u_inFIFO/n263 ,
         \u_inFIFO/n262 , \u_inFIFO/n261 , \u_inFIFO/n260 , \u_inFIFO/n259 ,
         \u_inFIFO/n258 , \u_inFIFO/n257 , \u_inFIFO/n256 , \u_inFIFO/n255 ,
         \u_inFIFO/n253 , \u_inFIFO/n252 , \u_inFIFO/n251 , \u_inFIFO/n250 ,
         \u_inFIFO/n249 , \u_inFIFO/n248 , \u_inFIFO/n247 , \u_inFIFO/n246 ,
         \u_inFIFO/n245 , \u_inFIFO/n243 , \u_inFIFO/n242 , \u_inFIFO/n241 ,
         \u_inFIFO/n240 , \u_inFIFO/n239 , \u_inFIFO/n238 , \u_inFIFO/n237 ,
         \u_inFIFO/n236 , \u_inFIFO/n235 , \u_inFIFO/n234 , \u_inFIFO/n233 ,
         \u_inFIFO/n232 , \u_inFIFO/n231 , \u_inFIFO/n230 , \u_inFIFO/n229 ,
         \u_inFIFO/n228 , \u_inFIFO/n227 , \u_inFIFO/n226 , \u_inFIFO/n225 ,
         \u_inFIFO/n224 , \u_inFIFO/n223 , \u_inFIFO/n222 , \u_inFIFO/n221 ,
         \u_inFIFO/n220 , \u_inFIFO/n219 , \u_inFIFO/n218 , \u_inFIFO/n217 ,
         \u_inFIFO/n216 , \u_inFIFO/n215 , \u_inFIFO/n214 , \u_inFIFO/n213 ,
         \u_inFIFO/n212 , \u_inFIFO/n211 , \u_inFIFO/n210 , \u_inFIFO/n209 ,
         \u_inFIFO/n208 , \u_inFIFO/n207 , \u_inFIFO/n206 , \u_inFIFO/n205 ,
         \u_inFIFO/n204 , \u_inFIFO/n203 , \u_inFIFO/n202 , \u_inFIFO/n201 ,
         \u_inFIFO/n200 , \u_inFIFO/n199 , \u_inFIFO/n198 , \u_inFIFO/n197 ,
         \u_inFIFO/n196 , \u_inFIFO/n195 , \u_inFIFO/n194 , \u_inFIFO/n193 ,
         \u_inFIFO/n192 , \u_inFIFO/n191 , \u_inFIFO/n190 , \u_inFIFO/n189 ,
         \u_inFIFO/n188 , \u_inFIFO/n187 , \u_inFIFO/n186 , \u_inFIFO/n185 ,
         \u_inFIFO/n184 , \u_inFIFO/n183 , \u_inFIFO/n182 , \u_inFIFO/n181 ,
         \u_inFIFO/n180 , \u_inFIFO/n179 , \u_inFIFO/n178 , \u_inFIFO/n177 ,
         \u_inFIFO/n176 , \u_inFIFO/n175 , \u_inFIFO/n174 , \u_inFIFO/n173 ,
         \u_inFIFO/n172 , \u_inFIFO/n171 , \u_inFIFO/n170 , \u_inFIFO/n169 ,
         \u_inFIFO/n168 , \u_inFIFO/n167 , \u_inFIFO/n166 , \u_inFIFO/n165 ,
         \u_inFIFO/n164 , \u_inFIFO/n163 , \u_inFIFO/n162 , \u_inFIFO/n161 ,
         \u_inFIFO/n160 , \u_inFIFO/n159 , \u_inFIFO/n158 , \u_inFIFO/n157 ,
         \u_inFIFO/n156 , \u_inFIFO/n155 , \u_inFIFO/n154 , \u_inFIFO/n153 ,
         \u_inFIFO/n152 , \u_inFIFO/n151 , \u_inFIFO/n150 , \u_inFIFO/n149 ,
         \u_inFIFO/n148 , \u_inFIFO/n147 , \u_inFIFO/n146 , \u_inFIFO/n145 ,
         \u_inFIFO/n144 , \u_inFIFO/n143 , \u_inFIFO/n142 , \u_inFIFO/n141 ,
         \u_inFIFO/n140 , \u_inFIFO/n139 , \u_inFIFO/n138 , \u_inFIFO/n137 ,
         \u_inFIFO/n136 , \u_inFIFO/n135 , \u_inFIFO/n134 , \u_inFIFO/n133 ,
         \u_inFIFO/n132 , \u_inFIFO/n131 , \u_inFIFO/n130 , \u_inFIFO/n129 ,
         \u_inFIFO/n128 , \u_inFIFO/n127 , \u_inFIFO/n126 , \u_inFIFO/n125 ,
         \u_inFIFO/n124 , \u_inFIFO/n123 , \u_inFIFO/n122 , \u_inFIFO/n121 ,
         \u_inFIFO/n120 , \u_inFIFO/n119 , \u_inFIFO/n118 , \u_inFIFO/n117 ,
         \u_inFIFO/n116 , \u_inFIFO/n115 , \u_inFIFO/n114 , \u_inFIFO/n113 ,
         \u_inFIFO/n112 , \u_inFIFO/n111 , \u_inFIFO/n110 , \u_inFIFO/n109 ,
         \u_inFIFO/n106 , \u_inFIFO/n101 , \u_inFIFO/n100 , \u_inFIFO/n99 ,
         \u_inFIFO/n98 , \u_inFIFO/n97 , \u_inFIFO/n96 , \u_inFIFO/n94 ,
         \u_inFIFO/n93 , \u_inFIFO/n86 , \u_inFIFO/n85 , \u_inFIFO/n84 ,
         \u_inFIFO/n83 , \u_inFIFO/n82 , \u_inFIFO/n78 , \u_inFIFO/n77 ,
         \u_inFIFO/n76 , \u_inFIFO/n73 , \u_inFIFO/n26 , \u_inFIFO/N249 ,
         \u_inFIFO/N195 , \u_inFIFO/N194 , \u_inFIFO/N193 , \u_inFIFO/N192 ,
         \u_inFIFO/N183 , \u_inFIFO/N182 , \u_inFIFO/N181 , \u_inFIFO/N180 ,
         \u_inFIFO/FIFO[31][3] , \u_inFIFO/FIFO[31][2] ,
         \u_inFIFO/FIFO[31][1] , \u_inFIFO/FIFO[31][0] ,
         \u_inFIFO/FIFO[30][3] , \u_inFIFO/FIFO[30][2] ,
         \u_inFIFO/FIFO[30][1] , \u_inFIFO/FIFO[30][0] ,
         \u_inFIFO/FIFO[29][3] , \u_inFIFO/FIFO[29][2] ,
         \u_inFIFO/FIFO[29][1] , \u_inFIFO/FIFO[29][0] ,
         \u_inFIFO/FIFO[28][3] , \u_inFIFO/FIFO[28][2] ,
         \u_inFIFO/FIFO[28][1] , \u_inFIFO/FIFO[28][0] ,
         \u_inFIFO/FIFO[27][3] , \u_inFIFO/FIFO[27][2] ,
         \u_inFIFO/FIFO[27][1] , \u_inFIFO/FIFO[27][0] ,
         \u_inFIFO/FIFO[26][3] , \u_inFIFO/FIFO[26][2] ,
         \u_inFIFO/FIFO[26][1] , \u_inFIFO/FIFO[26][0] ,
         \u_inFIFO/FIFO[25][3] , \u_inFIFO/FIFO[25][2] ,
         \u_inFIFO/FIFO[25][1] , \u_inFIFO/FIFO[25][0] ,
         \u_inFIFO/FIFO[24][3] , \u_inFIFO/FIFO[24][2] ,
         \u_inFIFO/FIFO[24][1] , \u_inFIFO/FIFO[24][0] ,
         \u_inFIFO/FIFO[23][3] , \u_inFIFO/FIFO[23][2] ,
         \u_inFIFO/FIFO[23][1] , \u_inFIFO/FIFO[23][0] ,
         \u_inFIFO/FIFO[22][3] , \u_inFIFO/FIFO[22][2] ,
         \u_inFIFO/FIFO[22][1] , \u_inFIFO/FIFO[22][0] ,
         \u_inFIFO/FIFO[21][3] , \u_inFIFO/FIFO[21][2] ,
         \u_inFIFO/FIFO[21][1] , \u_inFIFO/FIFO[21][0] ,
         \u_inFIFO/FIFO[20][3] , \u_inFIFO/FIFO[20][2] ,
         \u_inFIFO/FIFO[20][1] , \u_inFIFO/FIFO[20][0] ,
         \u_inFIFO/FIFO[19][3] , \u_inFIFO/FIFO[19][2] ,
         \u_inFIFO/FIFO[19][1] , \u_inFIFO/FIFO[19][0] ,
         \u_inFIFO/FIFO[18][3] , \u_inFIFO/FIFO[18][2] ,
         \u_inFIFO/FIFO[18][1] , \u_inFIFO/FIFO[18][0] ,
         \u_inFIFO/FIFO[17][3] , \u_inFIFO/FIFO[17][2] ,
         \u_inFIFO/FIFO[17][1] , \u_inFIFO/FIFO[17][0] ,
         \u_inFIFO/FIFO[16][3] , \u_inFIFO/FIFO[16][2] ,
         \u_inFIFO/FIFO[16][1] , \u_inFIFO/FIFO[16][0] ,
         \u_inFIFO/FIFO[15][3] , \u_inFIFO/FIFO[15][2] ,
         \u_inFIFO/FIFO[15][1] , \u_inFIFO/FIFO[15][0] ,
         \u_inFIFO/FIFO[14][3] , \u_inFIFO/FIFO[14][2] ,
         \u_inFIFO/FIFO[14][1] , \u_inFIFO/FIFO[14][0] ,
         \u_inFIFO/FIFO[13][3] , \u_inFIFO/FIFO[13][2] ,
         \u_inFIFO/FIFO[13][1] , \u_inFIFO/FIFO[13][0] ,
         \u_inFIFO/FIFO[12][3] , \u_inFIFO/FIFO[12][2] ,
         \u_inFIFO/FIFO[12][1] , \u_inFIFO/FIFO[12][0] ,
         \u_inFIFO/FIFO[11][3] , \u_inFIFO/FIFO[11][2] ,
         \u_inFIFO/FIFO[11][1] , \u_inFIFO/FIFO[11][0] ,
         \u_inFIFO/FIFO[10][3] , \u_inFIFO/FIFO[10][2] ,
         \u_inFIFO/FIFO[10][1] , \u_inFIFO/FIFO[10][0] , \u_inFIFO/FIFO[9][3] ,
         \u_inFIFO/FIFO[9][2] , \u_inFIFO/FIFO[9][1] , \u_inFIFO/FIFO[9][0] ,
         \u_inFIFO/FIFO[8][3] , \u_inFIFO/FIFO[8][2] , \u_inFIFO/FIFO[8][1] ,
         \u_inFIFO/FIFO[8][0] , \u_inFIFO/FIFO[7][3] , \u_inFIFO/FIFO[7][2] ,
         \u_inFIFO/FIFO[7][1] , \u_inFIFO/FIFO[7][0] , \u_inFIFO/FIFO[6][3] ,
         \u_inFIFO/FIFO[6][2] , \u_inFIFO/FIFO[6][1] , \u_inFIFO/FIFO[6][0] ,
         \u_inFIFO/FIFO[5][3] , \u_inFIFO/FIFO[5][2] , \u_inFIFO/FIFO[5][1] ,
         \u_inFIFO/FIFO[5][0] , \u_inFIFO/FIFO[4][3] , \u_inFIFO/FIFO[4][2] ,
         \u_inFIFO/FIFO[4][1] , \u_inFIFO/FIFO[4][0] , \u_inFIFO/FIFO[3][3] ,
         \u_inFIFO/FIFO[3][2] , \u_inFIFO/FIFO[3][1] , \u_inFIFO/FIFO[3][0] ,
         \u_inFIFO/FIFO[2][3] , \u_inFIFO/FIFO[2][2] , \u_inFIFO/FIFO[2][1] ,
         \u_inFIFO/FIFO[2][0] , \u_inFIFO/FIFO[1][3] , \u_inFIFO/FIFO[1][2] ,
         \u_inFIFO/FIFO[1][1] , \u_inFIFO/FIFO[1][0] , \u_inFIFO/FIFO[0][3] ,
         \u_inFIFO/FIFO[0][2] , \u_inFIFO/FIFO[0][1] , \u_inFIFO/FIFO[0][0] ,
         \u_inFIFO/N176 , \u_inFIFO/N135 , \u_inFIFO/N134 , \u_inFIFO/N133 ,
         \u_inFIFO/N132 , \u_inFIFO/N131 , \u_inFIFO/N128 , \u_inFIFO/N127 ,
         \u_inFIFO/N126 , \u_inFIFO/N125 , \u_inFIFO/N124 , \u_inFIFO/N123 ,
         \u_inFIFO/N121 , \u_inFIFO/N120 , \u_inFIFO/N119 , \u_inFIFO/N118 ,
         \u_inFIFO/N116 , \u_inFIFO/N115 , \u_inFIFO/N114 , \u_inFIFO/N113 ,
         \u_inFIFO/sigEnableCounter , \u_inFIFO/N44 , \u_inFIFO/N43 ,
         \u_inFIFO/N42 , \u_inFIFO/N41 , \u_inFIFO/sig_fsm_start_W ,
         \u_inFIFO/sig_fsm_start_R , \u_inFIFO/outReadCount[0] ,
         \u_inFIFO/outReadCount[1] , \u_inFIFO/outReadCount[2] ,
         \u_inFIFO/outReadCount[3] , \u_inFIFO/outReadCount[4] ,
         \u_inFIFO/outWriteCount[0] , \u_inFIFO/outWriteCount[1] ,
         \u_inFIFO/outWriteCount[2] , \u_inFIFO/outWriteCount[3] ,
         \u_inFIFO/outWriteCount[4] , \u_inFIFO/outWriteCount[5] ,
         \u_inFIFO/N39 , \u_inFIFO/N38 , \u_inFIFO/N37 , \u_inFIFO/N36 ,
         \u_inFIFO/N35 , \u_inFIFO/N34 , \u_coder/n374 , \u_coder/n373 ,
         \u_coder/n372 , \u_coder/n371 , \u_coder/n370 , \u_coder/n369 ,
         \u_coder/n368 , \u_coder/n367 , \u_coder/n366 , \u_coder/n365 ,
         \u_coder/n364 , \u_coder/n363 , \u_coder/n362 , \u_coder/n361 ,
         \u_coder/n360 , \u_coder/n359 , \u_coder/n358 , \u_coder/n357 ,
         \u_coder/n356 , \u_coder/n355 , \u_coder/n354 , \u_coder/n353 ,
         \u_coder/n352 , \u_coder/n351 , \u_coder/n350 , \u_coder/n349 ,
         \u_coder/n348 , \u_coder/n347 , \u_coder/n346 , \u_coder/n345 ,
         \u_coder/n344 , \u_coder/n343 , \u_coder/n342 , \u_coder/n341 ,
         \u_coder/n340 , \u_coder/n339 , \u_coder/n338 , \u_coder/n337 ,
         \u_coder/n336 , \u_coder/n335 , \u_coder/n334 , \u_coder/n333 ,
         \u_coder/n332 , \u_coder/n331 , \u_coder/n330 , \u_coder/n329 ,
         \u_coder/n328 , \u_coder/n327 , \u_coder/n326 , \u_coder/n325 ,
         \u_coder/n324 , \u_coder/n323 , \u_coder/n322 , \u_coder/n321 ,
         \u_coder/n320 , \u_coder/n319 , \u_coder/n318 , \u_coder/n317 ,
         \u_coder/n316 , \u_coder/n315 , \u_coder/n314 , \u_coder/n313 ,
         \u_coder/n312 , \u_coder/n311 , \u_coder/n310 , \u_coder/n309 ,
         \u_coder/n308 , \u_coder/n307 , \u_coder/n306 , \u_coder/n305 ,
         \u_coder/n304 , \u_coder/n303 , \u_coder/n302 , \u_coder/n301 ,
         \u_coder/n300 , \u_coder/n299 , \u_coder/n298 , \u_coder/n297 ,
         \u_coder/n296 , \u_coder/n295 , \u_coder/n294 , \u_coder/n293 ,
         \u_coder/n292 , \u_coder/n291 , \u_coder/n290 , \u_coder/n289 ,
         \u_coder/n288 , \u_coder/n287 , \u_coder/n286 , \u_coder/n284 ,
         \u_coder/n283 , \u_coder/n282 , \u_coder/n281 , \u_coder/n280 ,
         \u_coder/n279 , \u_coder/n278 , \u_coder/n277 , \u_coder/n276 ,
         \u_coder/n275 , \u_coder/n274 , \u_coder/n273 , \u_coder/n272 ,
         \u_coder/n271 , \u_coder/n270 , \u_coder/n269 , \u_coder/n268 ,
         \u_coder/n267 , \u_coder/n266 , \u_coder/n265 , \u_coder/n264 ,
         \u_coder/n263 , \u_coder/n262 , \u_coder/n261 , \u_coder/n260 ,
         \u_coder/n259 , \u_coder/n258 , \u_coder/n257 , \u_coder/n256 ,
         \u_coder/n255 , \u_coder/n254 , \u_coder/n253 , \u_coder/n252 ,
         \u_coder/n251 , \u_coder/n250 , \u_coder/n249 , \u_coder/n248 ,
         \u_coder/n247 , \u_coder/n246 , \u_coder/n245 , \u_coder/n244 ,
         \u_coder/n243 , \u_coder/n242 , \u_coder/n241 , \u_coder/n240 ,
         \u_coder/n239 , \u_coder/n238 , \u_coder/n236 , \u_coder/n234 ,
         \u_coder/n233 , \u_coder/n232 , \u_coder/n231 , \u_coder/n230 ,
         \u_coder/n229 , \u_coder/n228 , \u_coder/n227 , \u_coder/n226 ,
         \u_coder/n225 , \u_coder/n224 , \u_coder/n223 , \u_coder/n222 ,
         \u_coder/n221 , \u_coder/n220 , \u_coder/n219 , \u_coder/n218 ,
         \u_coder/n217 , \u_coder/n216 , \u_coder/n215 , \u_coder/n214 ,
         \u_coder/n213 , \u_coder/n212 , \u_coder/n211 , \u_coder/n210 ,
         \u_coder/n209 , \u_coder/n208 , \u_coder/n207 , \u_coder/n206 ,
         \u_coder/n205 , \u_coder/n204 , \u_coder/n203 , \u_coder/n202 ,
         \u_coder/n201 , \u_coder/n200 , \u_coder/n199 , \u_coder/n198 ,
         \u_coder/n197 , \u_coder/n196 , \u_coder/n195 , \u_coder/n194 ,
         \u_coder/n193 , \u_coder/n192 , \u_coder/n189 , \u_coder/n188 ,
         \u_coder/n187 , \u_coder/n186 , \u_coder/n185 , \u_coder/n184 ,
         \u_coder/n183 , \u_coder/n182 , \u_coder/n181 , \u_coder/n180 ,
         \u_coder/n179 , \u_coder/n178 , \u_coder/n177 , \u_coder/n176 ,
         \u_coder/n175 , \u_coder/n174 , \u_coder/n173 , \u_coder/n172 ,
         \u_coder/n171 , \u_coder/n170 , \u_coder/n169 , \u_coder/n168 ,
         \u_coder/n167 , \u_coder/n166 , \u_coder/n165 , \u_coder/n164 ,
         \u_coder/n163 , \u_coder/n162 , \u_coder/n161 , \u_coder/n160 ,
         \u_coder/n159 , \u_coder/n158 , \u_coder/n157 , \u_coder/n156 ,
         \u_coder/n155 , \u_coder/n154 , \u_coder/n153 , \u_coder/n152 ,
         \u_coder/n148 , \u_coder/n147 , \u_coder/n146 , \u_coder/n145 ,
         \u_coder/n144 , \u_coder/n141 , \u_coder/n140 , \u_coder/n139 ,
         \u_coder/n138 , \u_coder/n137 , \u_coder/n135 , \u_coder/n134 ,
         \u_coder/n131 , \u_coder/n130 , \u_coder/n129 , \u_coder/n128 ,
         \u_coder/n127 , \u_coder/n126 , \u_coder/n125 , \u_coder/n124 ,
         \u_coder/n123 , \u_coder/n122 , \u_coder/n121 , \u_coder/n120 ,
         \u_coder/n119 , \u_coder/n118 , \u_coder/n117 , \u_coder/n90 ,
         \u_coder/n89 , \u_coder/n88 , \u_coder/n86 , \u_coder/n85 ,
         \u_coder/n76 , \u_coder/n72 , \u_coder/n69 , \u_coder/n33 ,
         \u_coder/N1149 , \u_coder/N1143 , \u_coder/N1031 , \u_coder/N1030 ,
         \u_coder/N1029 , \u_coder/N1028 , \u_coder/N1027 , \u_coder/N1026 ,
         \u_coder/N1025 , \u_coder/N1024 , \u_coder/N1023 , \u_coder/N1022 ,
         \u_coder/N1021 , \u_coder/N1020 , \u_coder/N1019 , \u_coder/N1018 ,
         \u_coder/N1017 , \u_coder/N1016 , \u_coder/N1015 , \u_coder/N1014 ,
         \u_coder/N974 , \u_coder/N726 , \u_coder/N725 , \u_coder/N724 ,
         \u_coder/N723 , \u_coder/N722 , \u_coder/N721 , \u_coder/N720 ,
         \u_coder/N719 , \u_coder/N718 , \u_coder/N717 , \u_coder/N716 ,
         \u_coder/N715 , \u_coder/N714 , \u_coder/N713 , \u_coder/N712 ,
         \u_coder/N711 , \u_coder/N710 , \u_coder/N709 , \u_coder/N708 ,
         \u_coder/N668 , \u_coder/N522 , \u_coder/N521 , \u_coder/N520 ,
         \u_coder/N519 , \u_coder/N518 , \u_coder/N517 , \u_coder/N516 ,
         \u_coder/N515 , \u_coder/N514 , \u_coder/N513 , \u_coder/N512 ,
         \u_coder/N511 , \u_coder/N510 , \u_coder/N509 , \u_coder/N508 ,
         \u_coder/N507 , \u_coder/N506 , \u_coder/N505 , \u_coder/N504 ,
         \u_coder/N503 , \u_coder/N501 , \u_coder/N499 , \u_coder/my_clk_10M ,
         \u_coder/old_i_data , \u_coder/is9 , \u_coder/isPositiveQ ,
         \u_coder/isPositiveI , \u_coder/sin_was_positiveQ ,
         \u_coder/sin_was_positiveI , \u_coder/IorQ , \u_coder/stateQ[0] ,
         \u_coder/stateI[0] , \u_coder/N476 , \u_coder/N475 , \u_coder/N474 ,
         \u_coder/N473 , \u_coder/N472 , \u_coder/N471 , \u_coder/N470 ,
         \u_coder/N469 , \u_coder/N468 , \u_coder/N467 , \u_coder/N466 ,
         \u_coder/N465 , \u_coder/N464 , \u_coder/N463 , \u_coder/N462 ,
         \u_coder/N461 , \u_coder/N460 , \u_coder/N459 , \u_coder/clk_10M ,
         \u_decoder/sample_ready , \u_cordic/n37 , \u_cordic/n36 ,
         \u_cordic/n35 , \u_cordic/n34 , \u_cordic/n33 , \u_cordic/n32 ,
         \u_cordic/n31 , \u_cordic/n30 , \u_cordic/n29 , \u_cordic/n28 ,
         \u_cordic/n27 , \u_cordic/n26 , \u_cordic/n25 , \u_cordic/n24 ,
         \u_cordic/n23 , \u_cordic/n22 , \u_cordic/n21 , \u_cordic/n20 ,
         \u_cordic/n19 , \u_cordic/n18 , \u_cordic/n17 , \u_cordic/n16 ,
         \u_cordic/n13 , \u_cordic/n12 , \u_cordic/n11 , \u_cordic/N17 ,
         \u_cordic/N16 , \u_cordic/N15 , \u_cordic/dir , \u_cdr/n58 ,
         \u_cdr/n57 , \u_cdr/n56 , \u_cdr/n55 , \u_cdr/n54 , \u_cdr/n53 ,
         \u_cdr/n52 , \u_cdr/n51 , \u_cdr/n50 , \u_cdr/n49 , \u_cdr/n48 ,
         \u_cdr/n47 , \u_cdr/n46 , \u_cdr/n45 , \u_cdr/n44 , \u_cdr/n43 ,
         \u_cdr/n42 , \u_cdr/n41 , \u_cdr/n40 , \u_cdr/n39 , \u_cdr/n38 ,
         \u_cdr/n37 , \u_cdr/n36 , \u_cdr/n35 , \u_cdr/n34 , \u_cdr/n33 ,
         \u_cdr/n32 , \u_cdr/n31 , \u_cdr/n30 , \u_cdr/n29 , \u_cdr/n28 ,
         \u_cdr/n27 , \u_cdr/n26 , \u_cdr/n25 , \u_cdr/n24 , \u_cdr/n23 ,
         \u_cdr/n22 , \u_cdr/n19 , \u_cdr/n18 , \u_cdr/n17 , \u_cdr/n16 ,
         \u_cdr/n15 , \u_cdr/n14 , \u_cdr/n3 , \u_cdr/N100 , \u_cdr/w_sE ,
         \u_cdr/w_sT , \u_cdr/dir , \u_cdr/flag , \u_outFIFO/n731 ,
         \u_outFIFO/n730 , \u_outFIFO/n729 , \u_outFIFO/n728 ,
         \u_outFIFO/n727 , \u_outFIFO/n726 , \u_outFIFO/n725 ,
         \u_outFIFO/n724 , \u_outFIFO/n723 , \u_outFIFO/n722 ,
         \u_outFIFO/n721 , \u_outFIFO/n720 , \u_outFIFO/n719 ,
         \u_outFIFO/n718 , \u_outFIFO/n717 , \u_outFIFO/n716 ,
         \u_outFIFO/n715 , \u_outFIFO/n714 , \u_outFIFO/n713 ,
         \u_outFIFO/n712 , \u_outFIFO/n711 , \u_outFIFO/n710 ,
         \u_outFIFO/n709 , \u_outFIFO/n708 , \u_outFIFO/n707 ,
         \u_outFIFO/n706 , \u_outFIFO/n705 , \u_outFIFO/n704 ,
         \u_outFIFO/n703 , \u_outFIFO/n702 , \u_outFIFO/n701 ,
         \u_outFIFO/n700 , \u_outFIFO/n699 , \u_outFIFO/n698 ,
         \u_outFIFO/n697 , \u_outFIFO/n696 , \u_outFIFO/n695 ,
         \u_outFIFO/n694 , \u_outFIFO/n693 , \u_outFIFO/n692 ,
         \u_outFIFO/n690 , \u_outFIFO/n689 , \u_outFIFO/n688 ,
         \u_outFIFO/n687 , \u_outFIFO/n686 , \u_outFIFO/n685 ,
         \u_outFIFO/n684 , \u_outFIFO/n683 , \u_outFIFO/n682 ,
         \u_outFIFO/n681 , \u_outFIFO/n680 , \u_outFIFO/n679 ,
         \u_outFIFO/n678 , \u_outFIFO/n677 , \u_outFIFO/n676 ,
         \u_outFIFO/n675 , \u_outFIFO/n674 , \u_outFIFO/n673 ,
         \u_outFIFO/n672 , \u_outFIFO/n671 , \u_outFIFO/n670 ,
         \u_outFIFO/n669 , \u_outFIFO/n668 , \u_outFIFO/n667 ,
         \u_outFIFO/n666 , \u_outFIFO/n665 , \u_outFIFO/n664 ,
         \u_outFIFO/n663 , \u_outFIFO/n662 , \u_outFIFO/n661 ,
         \u_outFIFO/n660 , \u_outFIFO/n659 , \u_outFIFO/n658 ,
         \u_outFIFO/n657 , \u_outFIFO/n656 , \u_outFIFO/n655 ,
         \u_outFIFO/n654 , \u_outFIFO/n653 , \u_outFIFO/n652 ,
         \u_outFIFO/n651 , \u_outFIFO/n650 , \u_outFIFO/n649 ,
         \u_outFIFO/n648 , \u_outFIFO/n647 , \u_outFIFO/n646 ,
         \u_outFIFO/n645 , \u_outFIFO/n644 , \u_outFIFO/n643 ,
         \u_outFIFO/n642 , \u_outFIFO/n641 , \u_outFIFO/n640 ,
         \u_outFIFO/n639 , \u_outFIFO/n638 , \u_outFIFO/n637 ,
         \u_outFIFO/n636 , \u_outFIFO/n635 , \u_outFIFO/n634 ,
         \u_outFIFO/n633 , \u_outFIFO/n632 , \u_outFIFO/n631 ,
         \u_outFIFO/n630 , \u_outFIFO/n629 , \u_outFIFO/n628 ,
         \u_outFIFO/n627 , \u_outFIFO/n626 , \u_outFIFO/n625 ,
         \u_outFIFO/n624 , \u_outFIFO/n623 , \u_outFIFO/n622 ,
         \u_outFIFO/n621 , \u_outFIFO/n620 , \u_outFIFO/n619 ,
         \u_outFIFO/n618 , \u_outFIFO/n617 , \u_outFIFO/n616 ,
         \u_outFIFO/n615 , \u_outFIFO/n614 , \u_outFIFO/n613 ,
         \u_outFIFO/n612 , \u_outFIFO/n611 , \u_outFIFO/n610 ,
         \u_outFIFO/n609 , \u_outFIFO/n608 , \u_outFIFO/n607 ,
         \u_outFIFO/n606 , \u_outFIFO/n605 , \u_outFIFO/n604 ,
         \u_outFIFO/n603 , \u_outFIFO/n602 , \u_outFIFO/n601 ,
         \u_outFIFO/n600 , \u_outFIFO/n599 , \u_outFIFO/n598 ,
         \u_outFIFO/n597 , \u_outFIFO/n596 , \u_outFIFO/n595 ,
         \u_outFIFO/n594 , \u_outFIFO/n593 , \u_outFIFO/n592 ,
         \u_outFIFO/n591 , \u_outFIFO/n590 , \u_outFIFO/n589 ,
         \u_outFIFO/n588 , \u_outFIFO/n587 , \u_outFIFO/n586 ,
         \u_outFIFO/n585 , \u_outFIFO/n584 , \u_outFIFO/n583 ,
         \u_outFIFO/n582 , \u_outFIFO/n581 , \u_outFIFO/n580 ,
         \u_outFIFO/n579 , \u_outFIFO/n578 , \u_outFIFO/n577 ,
         \u_outFIFO/n576 , \u_outFIFO/n575 , \u_outFIFO/n574 ,
         \u_outFIFO/n573 , \u_outFIFO/n572 , \u_outFIFO/n571 ,
         \u_outFIFO/n570 , \u_outFIFO/n569 , \u_outFIFO/n568 ,
         \u_outFIFO/n567 , \u_outFIFO/n566 , \u_outFIFO/n565 ,
         \u_outFIFO/n564 , \u_outFIFO/n563 , \u_outFIFO/n562 ,
         \u_outFIFO/n561 , \u_outFIFO/n560 , \u_outFIFO/n559 ,
         \u_outFIFO/n558 , \u_outFIFO/n557 , \u_outFIFO/n556 ,
         \u_outFIFO/n555 , \u_outFIFO/n554 , \u_outFIFO/n553 ,
         \u_outFIFO/n552 , \u_outFIFO/n551 , \u_outFIFO/n549 ,
         \u_outFIFO/n548 , \u_outFIFO/n547 , \u_outFIFO/n546 ,
         \u_outFIFO/n545 , \u_outFIFO/n544 , \u_outFIFO/n543 ,
         \u_outFIFO/n542 , \u_outFIFO/n541 , \u_outFIFO/n540 ,
         \u_outFIFO/n539 , \u_outFIFO/n538 , \u_outFIFO/n537 ,
         \u_outFIFO/n536 , \u_outFIFO/n535 , \u_outFIFO/n534 ,
         \u_outFIFO/n533 , \u_outFIFO/n532 , \u_outFIFO/n531 ,
         \u_outFIFO/n530 , \u_outFIFO/n529 , \u_outFIFO/n528 ,
         \u_outFIFO/n527 , \u_outFIFO/n526 , \u_outFIFO/n525 ,
         \u_outFIFO/n524 , \u_outFIFO/n523 , \u_outFIFO/n522 ,
         \u_outFIFO/n521 , \u_outFIFO/n520 , \u_outFIFO/n519 ,
         \u_outFIFO/n518 , \u_outFIFO/n517 , \u_outFIFO/n516 ,
         \u_outFIFO/n515 , \u_outFIFO/n514 , \u_outFIFO/n513 ,
         \u_outFIFO/n512 , \u_outFIFO/n511 , \u_outFIFO/n510 ,
         \u_outFIFO/n509 , \u_outFIFO/n508 , \u_outFIFO/n507 ,
         \u_outFIFO/n506 , \u_outFIFO/n505 , \u_outFIFO/n504 ,
         \u_outFIFO/n503 , \u_outFIFO/n502 , \u_outFIFO/n501 ,
         \u_outFIFO/n500 , \u_outFIFO/n499 , \u_outFIFO/n498 ,
         \u_outFIFO/n497 , \u_outFIFO/n496 , \u_outFIFO/n495 ,
         \u_outFIFO/n494 , \u_outFIFO/n493 , \u_outFIFO/n492 ,
         \u_outFIFO/n491 , \u_outFIFO/n490 , \u_outFIFO/n489 ,
         \u_outFIFO/n488 , \u_outFIFO/n487 , \u_outFIFO/n486 ,
         \u_outFIFO/n485 , \u_outFIFO/n484 , \u_outFIFO/n483 ,
         \u_outFIFO/n482 , \u_outFIFO/n481 , \u_outFIFO/n480 ,
         \u_outFIFO/n479 , \u_outFIFO/n478 , \u_outFIFO/n477 ,
         \u_outFIFO/n476 , \u_outFIFO/n475 , \u_outFIFO/n474 ,
         \u_outFIFO/n473 , \u_outFIFO/n472 , \u_outFIFO/n471 ,
         \u_outFIFO/n470 , \u_outFIFO/n469 , \u_outFIFO/n468 ,
         \u_outFIFO/n467 , \u_outFIFO/n466 , \u_outFIFO/n465 ,
         \u_outFIFO/n464 , \u_outFIFO/n463 , \u_outFIFO/n462 ,
         \u_outFIFO/n461 , \u_outFIFO/n460 , \u_outFIFO/n459 ,
         \u_outFIFO/n458 , \u_outFIFO/n457 , \u_outFIFO/n456 ,
         \u_outFIFO/n455 , \u_outFIFO/n454 , \u_outFIFO/n453 ,
         \u_outFIFO/n452 , \u_outFIFO/n451 , \u_outFIFO/n450 ,
         \u_outFIFO/n449 , \u_outFIFO/n448 , \u_outFIFO/n447 ,
         \u_outFIFO/n446 , \u_outFIFO/n445 , \u_outFIFO/n444 ,
         \u_outFIFO/n443 , \u_outFIFO/n442 , \u_outFIFO/n441 ,
         \u_outFIFO/n440 , \u_outFIFO/n439 , \u_outFIFO/n438 ,
         \u_outFIFO/n437 , \u_outFIFO/n436 , \u_outFIFO/n435 ,
         \u_outFIFO/n434 , \u_outFIFO/n433 , \u_outFIFO/n432 ,
         \u_outFIFO/n431 , \u_outFIFO/n430 , \u_outFIFO/n429 ,
         \u_outFIFO/n428 , \u_outFIFO/n427 , \u_outFIFO/n426 ,
         \u_outFIFO/n425 , \u_outFIFO/n424 , \u_outFIFO/n423 ,
         \u_outFIFO/n422 , \u_outFIFO/n421 , \u_outFIFO/n420 ,
         \u_outFIFO/n419 , \u_outFIFO/n418 , \u_outFIFO/n417 ,
         \u_outFIFO/n416 , \u_outFIFO/n415 , \u_outFIFO/n414 ,
         \u_outFIFO/n413 , \u_outFIFO/n412 , \u_outFIFO/n411 ,
         \u_outFIFO/n410 , \u_outFIFO/n409 , \u_outFIFO/n408 ,
         \u_outFIFO/n407 , \u_outFIFO/n406 , \u_outFIFO/n405 ,
         \u_outFIFO/n404 , \u_outFIFO/n403 , \u_outFIFO/n402 ,
         \u_outFIFO/n401 , \u_outFIFO/n400 , \u_outFIFO/n399 ,
         \u_outFIFO/n398 , \u_outFIFO/n397 , \u_outFIFO/n396 ,
         \u_outFIFO/n395 , \u_outFIFO/n394 , \u_outFIFO/n393 ,
         \u_outFIFO/n392 , \u_outFIFO/n391 , \u_outFIFO/n390 ,
         \u_outFIFO/n389 , \u_outFIFO/n388 , \u_outFIFO/n387 ,
         \u_outFIFO/n386 , \u_outFIFO/n385 , \u_outFIFO/n384 ,
         \u_outFIFO/n383 , \u_outFIFO/n382 , \u_outFIFO/n381 ,
         \u_outFIFO/n380 , \u_outFIFO/n379 , \u_outFIFO/n378 ,
         \u_outFIFO/n377 , \u_outFIFO/n376 , \u_outFIFO/n375 ,
         \u_outFIFO/n374 , \u_outFIFO/n373 , \u_outFIFO/n372 ,
         \u_outFIFO/n371 , \u_outFIFO/n370 , \u_outFIFO/n369 ,
         \u_outFIFO/n368 , \u_outFIFO/n367 , \u_outFIFO/n366 ,
         \u_outFIFO/n365 , \u_outFIFO/n364 , \u_outFIFO/n363 ,
         \u_outFIFO/n362 , \u_outFIFO/n361 , \u_outFIFO/n360 ,
         \u_outFIFO/n359 , \u_outFIFO/n358 , \u_outFIFO/n357 ,
         \u_outFIFO/n356 , \u_outFIFO/n355 , \u_outFIFO/n354 ,
         \u_outFIFO/n353 , \u_outFIFO/n352 , \u_outFIFO/n351 ,
         \u_outFIFO/n350 , \u_outFIFO/n349 , \u_outFIFO/n348 ,
         \u_outFIFO/n347 , \u_outFIFO/n346 , \u_outFIFO/n345 ,
         \u_outFIFO/n344 , \u_outFIFO/n343 , \u_outFIFO/n342 ,
         \u_outFIFO/n341 , \u_outFIFO/n340 , \u_outFIFO/n339 ,
         \u_outFIFO/n338 , \u_outFIFO/n337 , \u_outFIFO/n336 ,
         \u_outFIFO/n335 , \u_outFIFO/n334 , \u_outFIFO/n333 ,
         \u_outFIFO/n332 , \u_outFIFO/n331 , \u_outFIFO/n330 ,
         \u_outFIFO/n329 , \u_outFIFO/n328 , \u_outFIFO/n327 ,
         \u_outFIFO/n326 , \u_outFIFO/n325 , \u_outFIFO/n324 ,
         \u_outFIFO/n323 , \u_outFIFO/n322 , \u_outFIFO/n321 ,
         \u_outFIFO/n320 , \u_outFIFO/n319 , \u_outFIFO/n318 ,
         \u_outFIFO/n317 , \u_outFIFO/n316 , \u_outFIFO/n315 ,
         \u_outFIFO/n314 , \u_outFIFO/n313 , \u_outFIFO/n312 ,
         \u_outFIFO/n311 , \u_outFIFO/n310 , \u_outFIFO/n309 ,
         \u_outFIFO/n308 , \u_outFIFO/n307 , \u_outFIFO/n306 ,
         \u_outFIFO/n305 , \u_outFIFO/n304 , \u_outFIFO/n303 ,
         \u_outFIFO/n302 , \u_outFIFO/n301 , \u_outFIFO/n300 ,
         \u_outFIFO/n299 , \u_outFIFO/n298 , \u_outFIFO/n297 ,
         \u_outFIFO/n296 , \u_outFIFO/n295 , \u_outFIFO/n294 ,
         \u_outFIFO/n293 , \u_outFIFO/n292 , \u_outFIFO/n291 ,
         \u_outFIFO/n290 , \u_outFIFO/n289 , \u_outFIFO/n288 ,
         \u_outFIFO/n287 , \u_outFIFO/n286 , \u_outFIFO/n285 ,
         \u_outFIFO/n284 , \u_outFIFO/n283 , \u_outFIFO/n282 ,
         \u_outFIFO/n281 , \u_outFIFO/n280 , \u_outFIFO/n279 ,
         \u_outFIFO/n278 , \u_outFIFO/n277 , \u_outFIFO/n276 ,
         \u_outFIFO/n275 , \u_outFIFO/n274 , \u_outFIFO/n273 ,
         \u_outFIFO/n272 , \u_outFIFO/n271 , \u_outFIFO/n270 ,
         \u_outFIFO/n269 , \u_outFIFO/n268 , \u_outFIFO/n267 ,
         \u_outFIFO/n266 , \u_outFIFO/n265 , \u_outFIFO/n264 ,
         \u_outFIFO/n263 , \u_outFIFO/n262 , \u_outFIFO/n261 ,
         \u_outFIFO/n260 , \u_outFIFO/n259 , \u_outFIFO/n258 ,
         \u_outFIFO/n257 , \u_outFIFO/n256 , \u_outFIFO/n255 ,
         \u_outFIFO/n254 , \u_outFIFO/n253 , \u_outFIFO/n252 ,
         \u_outFIFO/n251 , \u_outFIFO/n250 , \u_outFIFO/n249 ,
         \u_outFIFO/n248 , \u_outFIFO/n247 , \u_outFIFO/n246 ,
         \u_outFIFO/n245 , \u_outFIFO/n244 , \u_outFIFO/n243 ,
         \u_outFIFO/n242 , \u_outFIFO/n241 , \u_outFIFO/n240 ,
         \u_outFIFO/n239 , \u_outFIFO/n238 , \u_outFIFO/n237 ,
         \u_outFIFO/n236 , \u_outFIFO/n235 , \u_outFIFO/n234 ,
         \u_outFIFO/n233 , \u_outFIFO/n232 , \u_outFIFO/n231 ,
         \u_outFIFO/n230 , \u_outFIFO/n229 , \u_outFIFO/n228 ,
         \u_outFIFO/n227 , \u_outFIFO/n226 , \u_outFIFO/n225 ,
         \u_outFIFO/n224 , \u_outFIFO/n223 , \u_outFIFO/n222 ,
         \u_outFIFO/n221 , \u_outFIFO/n220 , \u_outFIFO/n219 ,
         \u_outFIFO/n218 , \u_outFIFO/n217 , \u_outFIFO/n216 ,
         \u_outFIFO/n215 , \u_outFIFO/n214 , \u_outFIFO/n213 ,
         \u_outFIFO/n212 , \u_outFIFO/n211 , \u_outFIFO/n210 ,
         \u_outFIFO/n209 , \u_outFIFO/n208 , \u_outFIFO/n207 ,
         \u_outFIFO/n206 , \u_outFIFO/n205 , \u_outFIFO/n197 ,
         \u_outFIFO/n196 , \u_outFIFO/n195 , \u_outFIFO/n194 ,
         \u_outFIFO/n193 , \u_outFIFO/n192 , \u_outFIFO/n191 ,
         \u_outFIFO/n185 , \u_outFIFO/n184 , \u_outFIFO/n183 ,
         \u_outFIFO/n182 , \u_outFIFO/n181 , \u_outFIFO/n180 ,
         \u_outFIFO/n178 , \u_outFIFO/n177 , \u_outFIFO/n176 ,
         \u_outFIFO/n174 , \u_outFIFO/n173 , \u_outFIFO/N474 ,
         \u_outFIFO/N473 , \u_outFIFO/N199 , \u_outFIFO/N198 ,
         \u_outFIFO/N197 , \u_outFIFO/N196 , \u_outFIFO/N185 ,
         \u_outFIFO/N184 , \u_outFIFO/N183 , \u_outFIFO/N182 ,
         \u_outFIFO/FIFO[31][3] , \u_outFIFO/FIFO[31][2] ,
         \u_outFIFO/FIFO[31][1] , \u_outFIFO/FIFO[31][0] ,
         \u_outFIFO/FIFO[30][3] , \u_outFIFO/FIFO[30][2] ,
         \u_outFIFO/FIFO[30][1] , \u_outFIFO/FIFO[30][0] ,
         \u_outFIFO/FIFO[29][3] , \u_outFIFO/FIFO[29][2] ,
         \u_outFIFO/FIFO[29][1] , \u_outFIFO/FIFO[29][0] ,
         \u_outFIFO/FIFO[28][3] , \u_outFIFO/FIFO[28][2] ,
         \u_outFIFO/FIFO[28][1] , \u_outFIFO/FIFO[28][0] ,
         \u_outFIFO/FIFO[27][3] , \u_outFIFO/FIFO[27][2] ,
         \u_outFIFO/FIFO[27][1] , \u_outFIFO/FIFO[27][0] ,
         \u_outFIFO/FIFO[26][3] , \u_outFIFO/FIFO[26][2] ,
         \u_outFIFO/FIFO[26][1] , \u_outFIFO/FIFO[26][0] ,
         \u_outFIFO/FIFO[25][3] , \u_outFIFO/FIFO[25][2] ,
         \u_outFIFO/FIFO[25][1] , \u_outFIFO/FIFO[25][0] ,
         \u_outFIFO/FIFO[24][3] , \u_outFIFO/FIFO[24][2] ,
         \u_outFIFO/FIFO[24][1] , \u_outFIFO/FIFO[24][0] ,
         \u_outFIFO/FIFO[23][3] , \u_outFIFO/FIFO[23][2] ,
         \u_outFIFO/FIFO[23][1] , \u_outFIFO/FIFO[23][0] ,
         \u_outFIFO/FIFO[22][3] , \u_outFIFO/FIFO[22][2] ,
         \u_outFIFO/FIFO[22][1] , \u_outFIFO/FIFO[22][0] ,
         \u_outFIFO/FIFO[21][3] , \u_outFIFO/FIFO[21][2] ,
         \u_outFIFO/FIFO[21][1] , \u_outFIFO/FIFO[21][0] ,
         \u_outFIFO/FIFO[20][3] , \u_outFIFO/FIFO[20][2] ,
         \u_outFIFO/FIFO[20][1] , \u_outFIFO/FIFO[20][0] ,
         \u_outFIFO/FIFO[19][3] , \u_outFIFO/FIFO[19][2] ,
         \u_outFIFO/FIFO[19][1] , \u_outFIFO/FIFO[19][0] ,
         \u_outFIFO/FIFO[18][3] , \u_outFIFO/FIFO[18][2] ,
         \u_outFIFO/FIFO[18][1] , \u_outFIFO/FIFO[18][0] ,
         \u_outFIFO/FIFO[17][3] , \u_outFIFO/FIFO[17][2] ,
         \u_outFIFO/FIFO[17][1] , \u_outFIFO/FIFO[17][0] ,
         \u_outFIFO/FIFO[16][3] , \u_outFIFO/FIFO[16][2] ,
         \u_outFIFO/FIFO[16][1] , \u_outFIFO/FIFO[16][0] ,
         \u_outFIFO/FIFO[15][3] , \u_outFIFO/FIFO[15][2] ,
         \u_outFIFO/FIFO[15][1] , \u_outFIFO/FIFO[15][0] ,
         \u_outFIFO/FIFO[14][3] , \u_outFIFO/FIFO[14][2] ,
         \u_outFIFO/FIFO[14][1] , \u_outFIFO/FIFO[14][0] ,
         \u_outFIFO/FIFO[13][3] , \u_outFIFO/FIFO[13][2] ,
         \u_outFIFO/FIFO[13][1] , \u_outFIFO/FIFO[13][0] ,
         \u_outFIFO/FIFO[12][3] , \u_outFIFO/FIFO[12][2] ,
         \u_outFIFO/FIFO[12][1] , \u_outFIFO/FIFO[12][0] ,
         \u_outFIFO/FIFO[11][3] , \u_outFIFO/FIFO[11][2] ,
         \u_outFIFO/FIFO[11][1] , \u_outFIFO/FIFO[11][0] ,
         \u_outFIFO/FIFO[10][3] , \u_outFIFO/FIFO[10][2] ,
         \u_outFIFO/FIFO[10][1] , \u_outFIFO/FIFO[10][0] ,
         \u_outFIFO/FIFO[9][3] , \u_outFIFO/FIFO[9][2] ,
         \u_outFIFO/FIFO[9][1] , \u_outFIFO/FIFO[9][0] ,
         \u_outFIFO/FIFO[8][3] , \u_outFIFO/FIFO[8][2] ,
         \u_outFIFO/FIFO[8][1] , \u_outFIFO/FIFO[8][0] ,
         \u_outFIFO/FIFO[7][3] , \u_outFIFO/FIFO[7][2] ,
         \u_outFIFO/FIFO[7][1] , \u_outFIFO/FIFO[7][0] ,
         \u_outFIFO/FIFO[6][3] , \u_outFIFO/FIFO[6][2] ,
         \u_outFIFO/FIFO[6][1] , \u_outFIFO/FIFO[6][0] ,
         \u_outFIFO/FIFO[5][3] , \u_outFIFO/FIFO[5][2] ,
         \u_outFIFO/FIFO[5][1] , \u_outFIFO/FIFO[5][0] ,
         \u_outFIFO/FIFO[4][3] , \u_outFIFO/FIFO[4][2] ,
         \u_outFIFO/FIFO[4][1] , \u_outFIFO/FIFO[4][0] ,
         \u_outFIFO/FIFO[3][3] , \u_outFIFO/FIFO[3][2] ,
         \u_outFIFO/FIFO[3][1] , \u_outFIFO/FIFO[3][0] ,
         \u_outFIFO/FIFO[2][3] , \u_outFIFO/FIFO[2][2] ,
         \u_outFIFO/FIFO[2][1] , \u_outFIFO/FIFO[2][0] ,
         \u_outFIFO/FIFO[1][3] , \u_outFIFO/FIFO[1][2] ,
         \u_outFIFO/FIFO[1][1] , \u_outFIFO/FIFO[1][0] ,
         \u_outFIFO/FIFO[0][3] , \u_outFIFO/FIFO[0][2] ,
         \u_outFIFO/FIFO[0][1] , \u_outFIFO/FIFO[0][0] , \u_outFIFO/N178 ,
         \u_outFIFO/N136 , \u_outFIFO/N135 , \u_outFIFO/N134 ,
         \u_outFIFO/N133 , \u_outFIFO/N132 , \u_outFIFO/N131 ,
         \u_outFIFO/N129 , \u_outFIFO/N128 , \u_outFIFO/N127 ,
         \u_outFIFO/N126 , \u_outFIFO/N122 , \u_outFIFO/N121 ,
         \u_outFIFO/N120 , \u_outFIFO/N118 , \u_outFIFO/N117 ,
         \u_outFIFO/N116 , \u_outFIFO/N115 , \u_outFIFO/N114 ,
         \u_outFIFO/sigEnableCounter , \u_outFIFO/N44 , \u_outFIFO/N43 ,
         \u_outFIFO/N42 , \u_outFIFO/N41 , \u_outFIFO/sig_fsm_start_W ,
         \u_outFIFO/sig_fsm_start_R , \u_outFIFO/outReadCount[0] ,
         \u_outFIFO/outReadCount[1] , \u_outFIFO/outReadCount[2] ,
         \u_outFIFO/outReadCount[3] , \u_outFIFO/outReadCount[4] ,
         \u_outFIFO/outWriteCount[0] , \u_outFIFO/outWriteCount[1] ,
         \u_outFIFO/outWriteCount[2] , \u_outFIFO/outWriteCount[3] ,
         \u_outFIFO/outWriteCount[4] , \u_outFIFO/outWriteCount[5] ,
         \u_outFIFO/N39 , \u_outFIFO/N38 , \u_outFIFO/N37 , \u_outFIFO/N36 ,
         \u_demux1/n5 , \u_demux1/n4 , \u_mux3/n3 , \u_mux8/n4 , \u_mux8/n3 ,
         \u_inFIFO/os1/sigQout2 , \u_inFIFO/os1/sigQout1 ,
         \u_decoder/iq_demod/n71 , \u_decoder/iq_demod/n70 ,
         \u_decoder/iq_demod/n69 , \u_decoder/iq_demod/n68 ,
         \u_decoder/iq_demod/n67 , \u_decoder/iq_demod/n66 ,
         \u_decoder/iq_demod/n65 , \u_decoder/iq_demod/n64 ,
         \u_decoder/iq_demod/n63 , \u_decoder/iq_demod/n62 ,
         \u_decoder/iq_demod/n61 , \u_decoder/iq_demod/n60 ,
         \u_decoder/iq_demod/n59 , \u_decoder/iq_demod/n58 ,
         \u_decoder/iq_demod/n57 , \u_decoder/iq_demod/n56 ,
         \u_decoder/iq_demod/n55 , \u_decoder/iq_demod/n54 ,
         \u_decoder/iq_demod/n53 , \u_decoder/iq_demod/n52 ,
         \u_decoder/iq_demod/n51 , \u_decoder/iq_demod/n50 ,
         \u_decoder/iq_demod/n49 , \u_decoder/iq_demod/n48 ,
         \u_decoder/iq_demod/n47 , \u_decoder/iq_demod/n46 ,
         \u_decoder/iq_demod/n45 , \u_decoder/iq_demod/n44 ,
         \u_decoder/iq_demod/n43 , \u_decoder/iq_demod/n42 ,
         \u_decoder/iq_demod/n41 , \u_decoder/iq_demod/n30 ,
         \u_decoder/iq_demod/I_if_buff[3] , \u_decoder/iq_demod/Q_if_buff[3] ,
         \u_decoder/iq_demod/N13 , \u_decoder/fir_filter/n1451 ,
         \u_decoder/fir_filter/n1450 , \u_decoder/fir_filter/n1449 ,
         \u_decoder/fir_filter/n1448 , \u_decoder/fir_filter/n1447 ,
         \u_decoder/fir_filter/n1446 , \u_decoder/fir_filter/n1445 ,
         \u_decoder/fir_filter/n1444 , \u_decoder/fir_filter/n1443 ,
         \u_decoder/fir_filter/n1442 , \u_decoder/fir_filter/n1441 ,
         \u_decoder/fir_filter/n1440 , \u_decoder/fir_filter/n1439 ,
         \u_decoder/fir_filter/n1438 , \u_decoder/fir_filter/n1437 ,
         \u_decoder/fir_filter/n1436 , \u_decoder/fir_filter/n1434 ,
         \u_decoder/fir_filter/n1433 , \u_decoder/fir_filter/n1432 ,
         \u_decoder/fir_filter/n1431 , \u_decoder/fir_filter/n1430 ,
         \u_decoder/fir_filter/n1429 , \u_decoder/fir_filter/n1428 ,
         \u_decoder/fir_filter/n1427 , \u_decoder/fir_filter/n1426 ,
         \u_decoder/fir_filter/n1425 , \u_decoder/fir_filter/n1424 ,
         \u_decoder/fir_filter/n1423 , \u_decoder/fir_filter/n1422 ,
         \u_decoder/fir_filter/n1421 , \u_decoder/fir_filter/n1420 ,
         \u_decoder/fir_filter/n1418 , \u_decoder/fir_filter/n1417 ,
         \u_decoder/fir_filter/n1416 , \u_decoder/fir_filter/n1415 ,
         \u_decoder/fir_filter/n1414 , \u_decoder/fir_filter/n1413 ,
         \u_decoder/fir_filter/n1412 , \u_decoder/fir_filter/n1411 ,
         \u_decoder/fir_filter/n1410 , \u_decoder/fir_filter/n1409 ,
         \u_decoder/fir_filter/n1408 , \u_decoder/fir_filter/n1407 ,
         \u_decoder/fir_filter/n1406 , \u_decoder/fir_filter/n1405 ,
         \u_decoder/fir_filter/n1402 , \u_decoder/fir_filter/n1401 ,
         \u_decoder/fir_filter/n1400 , \u_decoder/fir_filter/n1399 ,
         \u_decoder/fir_filter/n1398 , \u_decoder/fir_filter/n1397 ,
         \u_decoder/fir_filter/n1396 , \u_decoder/fir_filter/n1395 ,
         \u_decoder/fir_filter/n1394 , \u_decoder/fir_filter/n1393 ,
         \u_decoder/fir_filter/n1392 , \u_decoder/fir_filter/n1391 ,
         \u_decoder/fir_filter/n1390 , \u_decoder/fir_filter/n1389 ,
         \u_decoder/fir_filter/n1388 , \u_decoder/fir_filter/n1386 ,
         \u_decoder/fir_filter/n1385 , \u_decoder/fir_filter/n1384 ,
         \u_decoder/fir_filter/n1383 , \u_decoder/fir_filter/n1382 ,
         \u_decoder/fir_filter/n1381 , \u_decoder/fir_filter/n1380 ,
         \u_decoder/fir_filter/n1379 , \u_decoder/fir_filter/n1378 ,
         \u_decoder/fir_filter/n1377 , \u_decoder/fir_filter/n1376 ,
         \u_decoder/fir_filter/n1375 , \u_decoder/fir_filter/n1374 ,
         \u_decoder/fir_filter/n1373 , \u_decoder/fir_filter/n1372 ,
         \u_decoder/fir_filter/n1370 , \u_decoder/fir_filter/n1369 ,
         \u_decoder/fir_filter/n1368 , \u_decoder/fir_filter/n1367 ,
         \u_decoder/fir_filter/n1366 , \u_decoder/fir_filter/n1365 ,
         \u_decoder/fir_filter/n1364 , \u_decoder/fir_filter/n1363 ,
         \u_decoder/fir_filter/n1362 , \u_decoder/fir_filter/n1361 ,
         \u_decoder/fir_filter/n1360 , \u_decoder/fir_filter/n1359 ,
         \u_decoder/fir_filter/n1358 , \u_decoder/fir_filter/n1357 ,
         \u_decoder/fir_filter/n1354 , \u_decoder/fir_filter/n1353 ,
         \u_decoder/fir_filter/n1352 , \u_decoder/fir_filter/n1351 ,
         \u_decoder/fir_filter/n1350 , \u_decoder/fir_filter/n1349 ,
         \u_decoder/fir_filter/n1348 , \u_decoder/fir_filter/n1347 ,
         \u_decoder/fir_filter/n1346 , \u_decoder/fir_filter/n1345 ,
         \u_decoder/fir_filter/n1344 , \u_decoder/fir_filter/n1343 ,
         \u_decoder/fir_filter/n1342 , \u_decoder/fir_filter/n1341 ,
         \u_decoder/fir_filter/n1340 , \u_decoder/fir_filter/n1338 ,
         \u_decoder/fir_filter/n1337 , \u_decoder/fir_filter/n1336 ,
         \u_decoder/fir_filter/n1335 , \u_decoder/fir_filter/n1334 ,
         \u_decoder/fir_filter/n1333 , \u_decoder/fir_filter/n1332 ,
         \u_decoder/fir_filter/n1331 , \u_decoder/fir_filter/n1330 ,
         \u_decoder/fir_filter/n1329 , \u_decoder/fir_filter/n1328 ,
         \u_decoder/fir_filter/n1327 , \u_decoder/fir_filter/n1326 ,
         \u_decoder/fir_filter/n1325 , \u_decoder/fir_filter/n1324 ,
         \u_decoder/fir_filter/n1317 , \u_decoder/fir_filter/n1316 ,
         \u_decoder/fir_filter/n1315 , \u_decoder/fir_filter/n1314 ,
         \u_decoder/fir_filter/n1313 , \u_decoder/fir_filter/n1312 ,
         \u_decoder/fir_filter/n1311 , \u_decoder/fir_filter/n1310 ,
         \u_decoder/fir_filter/n1309 , \u_decoder/fir_filter/n1308 ,
         \u_decoder/fir_filter/n1307 , \u_decoder/fir_filter/n1306 ,
         \u_decoder/fir_filter/n1305 , \u_decoder/fir_filter/n1304 ,
         \u_decoder/fir_filter/n1303 , \u_decoder/fir_filter/n1302 ,
         \u_decoder/fir_filter/n1301 , \u_decoder/fir_filter/n1300 ,
         \u_decoder/fir_filter/n1299 , \u_decoder/fir_filter/n1298 ,
         \u_decoder/fir_filter/n1297 , \u_decoder/fir_filter/n1296 ,
         \u_decoder/fir_filter/n1295 , \u_decoder/fir_filter/n1294 ,
         \u_decoder/fir_filter/n1293 , \u_decoder/fir_filter/n1292 ,
         \u_decoder/fir_filter/n1291 , \u_decoder/fir_filter/n1290 ,
         \u_decoder/fir_filter/n1289 , \u_decoder/fir_filter/n1288 ,
         \u_decoder/fir_filter/n1286 , \u_decoder/fir_filter/n1285 ,
         \u_decoder/fir_filter/n1284 , \u_decoder/fir_filter/n1283 ,
         \u_decoder/fir_filter/n1282 , \u_decoder/fir_filter/n1281 ,
         \u_decoder/fir_filter/n1280 , \u_decoder/fir_filter/n1279 ,
         \u_decoder/fir_filter/n1278 , \u_decoder/fir_filter/n1277 ,
         \u_decoder/fir_filter/n1276 , \u_decoder/fir_filter/n1275 ,
         \u_decoder/fir_filter/n1274 , \u_decoder/fir_filter/n1273 ,
         \u_decoder/fir_filter/n1272 , \u_decoder/fir_filter/n1270 ,
         \u_decoder/fir_filter/n1269 , \u_decoder/fir_filter/n1268 ,
         \u_decoder/fir_filter/n1267 , \u_decoder/fir_filter/n1266 ,
         \u_decoder/fir_filter/n1265 , \u_decoder/fir_filter/n1264 ,
         \u_decoder/fir_filter/n1263 , \u_decoder/fir_filter/n1262 ,
         \u_decoder/fir_filter/n1261 , \u_decoder/fir_filter/n1260 ,
         \u_decoder/fir_filter/n1259 , \u_decoder/fir_filter/n1258 ,
         \u_decoder/fir_filter/n1257 , \u_decoder/fir_filter/n1254 ,
         \u_decoder/fir_filter/n1253 , \u_decoder/fir_filter/n1252 ,
         \u_decoder/fir_filter/n1251 , \u_decoder/fir_filter/n1250 ,
         \u_decoder/fir_filter/n1249 , \u_decoder/fir_filter/n1248 ,
         \u_decoder/fir_filter/n1247 , \u_decoder/fir_filter/n1246 ,
         \u_decoder/fir_filter/n1245 , \u_decoder/fir_filter/n1244 ,
         \u_decoder/fir_filter/n1243 , \u_decoder/fir_filter/n1242 ,
         \u_decoder/fir_filter/n1241 , \u_decoder/fir_filter/n1240 ,
         \u_decoder/fir_filter/n1238 , \u_decoder/fir_filter/n1237 ,
         \u_decoder/fir_filter/n1236 , \u_decoder/fir_filter/n1235 ,
         \u_decoder/fir_filter/n1234 , \u_decoder/fir_filter/n1233 ,
         \u_decoder/fir_filter/n1232 , \u_decoder/fir_filter/n1231 ,
         \u_decoder/fir_filter/n1230 , \u_decoder/fir_filter/n1229 ,
         \u_decoder/fir_filter/n1228 , \u_decoder/fir_filter/n1227 ,
         \u_decoder/fir_filter/n1226 , \u_decoder/fir_filter/n1225 ,
         \u_decoder/fir_filter/n1224 , \u_decoder/fir_filter/n1222 ,
         \u_decoder/fir_filter/n1221 , \u_decoder/fir_filter/n1220 ,
         \u_decoder/fir_filter/n1219 , \u_decoder/fir_filter/n1218 ,
         \u_decoder/fir_filter/n1217 , \u_decoder/fir_filter/n1216 ,
         \u_decoder/fir_filter/n1215 , \u_decoder/fir_filter/n1214 ,
         \u_decoder/fir_filter/n1213 , \u_decoder/fir_filter/n1212 ,
         \u_decoder/fir_filter/n1211 , \u_decoder/fir_filter/n1210 ,
         \u_decoder/fir_filter/n1209 , \u_decoder/fir_filter/n1206 ,
         \u_decoder/fir_filter/n1205 , \u_decoder/fir_filter/n1204 ,
         \u_decoder/fir_filter/n1203 , \u_decoder/fir_filter/n1202 ,
         \u_decoder/fir_filter/n1201 , \u_decoder/fir_filter/n1200 ,
         \u_decoder/fir_filter/n1199 , \u_decoder/fir_filter/n1198 ,
         \u_decoder/fir_filter/n1197 , \u_decoder/fir_filter/n1196 ,
         \u_decoder/fir_filter/n1195 , \u_decoder/fir_filter/n1194 ,
         \u_decoder/fir_filter/n1193 , \u_decoder/fir_filter/n1192 ,
         \u_decoder/fir_filter/n1190 , \u_decoder/fir_filter/n1189 ,
         \u_decoder/fir_filter/n1188 , \u_decoder/fir_filter/n1187 ,
         \u_decoder/fir_filter/n1186 , \u_decoder/fir_filter/n1185 ,
         \u_decoder/fir_filter/n1184 , \u_decoder/fir_filter/n1183 ,
         \u_decoder/fir_filter/n1182 , \u_decoder/fir_filter/n1181 ,
         \u_decoder/fir_filter/n1180 , \u_decoder/fir_filter/n1179 ,
         \u_decoder/fir_filter/n1178 , \u_decoder/fir_filter/n1177 ,
         \u_decoder/fir_filter/n1176 , \u_decoder/fir_filter/n1169 ,
         \u_decoder/fir_filter/n1168 , \u_decoder/fir_filter/n1167 ,
         \u_decoder/fir_filter/n1166 , \u_decoder/fir_filter/n1165 ,
         \u_decoder/fir_filter/n1164 , \u_decoder/fir_filter/n1163 ,
         \u_decoder/fir_filter/n1162 , \u_decoder/fir_filter/n1161 ,
         \u_decoder/fir_filter/n1160 , \u_decoder/fir_filter/n1159 ,
         \u_decoder/fir_filter/n1158 , \u_decoder/fir_filter/n1157 ,
         \u_decoder/fir_filter/n1156 , \u_decoder/fir_filter/n1155 ,
         \u_decoder/fir_filter/n1154 , \u_decoder/fir_filter/n1153 ,
         \u_decoder/fir_filter/n1152 , \u_decoder/fir_filter/n1151 ,
         \u_decoder/fir_filter/n1150 , \u_decoder/fir_filter/n1149 ,
         \u_decoder/fir_filter/n1148 , \u_decoder/fir_filter/n1147 ,
         \u_decoder/fir_filter/n1146 , \u_decoder/fir_filter/n1145 ,
         \u_decoder/fir_filter/n1144 , \u_decoder/fir_filter/n1143 ,
         \u_decoder/fir_filter/n1142 , \u_decoder/fir_filter/n1141 ,
         \u_decoder/fir_filter/n1140 , \u_decoder/fir_filter/n1139 ,
         \u_decoder/fir_filter/n1138 , \u_decoder/fir_filter/n1137 ,
         \u_decoder/fir_filter/n1136 , \u_decoder/fir_filter/n1135 ,
         \u_decoder/fir_filter/n1134 , \u_decoder/fir_filter/n1132 ,
         \u_decoder/fir_filter/n1131 , \u_decoder/fir_filter/n1130 ,
         \u_decoder/fir_filter/n1129 , \u_decoder/fir_filter/n1128 ,
         \u_decoder/fir_filter/n1127 , \u_decoder/fir_filter/n1126 ,
         \u_decoder/fir_filter/n1125 , \u_decoder/fir_filter/n1124 ,
         \u_decoder/fir_filter/n1123 , \u_decoder/fir_filter/n1122 ,
         \u_decoder/fir_filter/n1121 , \u_decoder/fir_filter/n1120 ,
         \u_decoder/fir_filter/n1119 , \u_decoder/fir_filter/n1118 ,
         \u_decoder/fir_filter/n1116 , \u_decoder/fir_filter/n1115 ,
         \u_decoder/fir_filter/n1114 , \u_decoder/fir_filter/n1113 ,
         \u_decoder/fir_filter/n1112 , \u_decoder/fir_filter/n1111 ,
         \u_decoder/fir_filter/n1110 , \u_decoder/fir_filter/n1109 ,
         \u_decoder/fir_filter/n1108 , \u_decoder/fir_filter/n1107 ,
         \u_decoder/fir_filter/n1106 , \u_decoder/fir_filter/n1105 ,
         \u_decoder/fir_filter/n1104 , \u_decoder/fir_filter/n1103 ,
         \u_decoder/fir_filter/n1102 , \u_decoder/fir_filter/n1100 ,
         \u_decoder/fir_filter/n1099 , \u_decoder/fir_filter/n1098 ,
         \u_decoder/fir_filter/n1097 , \u_decoder/fir_filter/n1096 ,
         \u_decoder/fir_filter/n1095 , \u_decoder/fir_filter/n1094 ,
         \u_decoder/fir_filter/n1093 , \u_decoder/fir_filter/n1092 ,
         \u_decoder/fir_filter/n1091 , \u_decoder/fir_filter/n1090 ,
         \u_decoder/fir_filter/n1089 , \u_decoder/fir_filter/n1088 ,
         \u_decoder/fir_filter/n1087 , \u_decoder/fir_filter/n1086 ,
         \u_decoder/fir_filter/n1084 , \u_decoder/fir_filter/n1083 ,
         \u_decoder/fir_filter/n1082 , \u_decoder/fir_filter/n1081 ,
         \u_decoder/fir_filter/n1080 , \u_decoder/fir_filter/n1079 ,
         \u_decoder/fir_filter/n1078 , \u_decoder/fir_filter/n1077 ,
         \u_decoder/fir_filter/n1076 , \u_decoder/fir_filter/n1075 ,
         \u_decoder/fir_filter/n1074 , \u_decoder/fir_filter/n1073 ,
         \u_decoder/fir_filter/n1072 , \u_decoder/fir_filter/n1071 ,
         \u_decoder/fir_filter/n1070 , \u_decoder/fir_filter/n1068 ,
         \u_decoder/fir_filter/n1067 , \u_decoder/fir_filter/n1066 ,
         \u_decoder/fir_filter/n1065 , \u_decoder/fir_filter/n1064 ,
         \u_decoder/fir_filter/n1063 , \u_decoder/fir_filter/n1062 ,
         \u_decoder/fir_filter/n1061 , \u_decoder/fir_filter/n1060 ,
         \u_decoder/fir_filter/n1059 , \u_decoder/fir_filter/n1058 ,
         \u_decoder/fir_filter/n1057 , \u_decoder/fir_filter/n1056 ,
         \u_decoder/fir_filter/n1055 , \u_decoder/fir_filter/n1054 ,
         \u_decoder/fir_filter/n1052 , \u_decoder/fir_filter/n1051 ,
         \u_decoder/fir_filter/n1050 , \u_decoder/fir_filter/n1049 ,
         \u_decoder/fir_filter/n1048 , \u_decoder/fir_filter/n1047 ,
         \u_decoder/fir_filter/n1046 , \u_decoder/fir_filter/n1045 ,
         \u_decoder/fir_filter/n1044 , \u_decoder/fir_filter/n1043 ,
         \u_decoder/fir_filter/n1042 , \u_decoder/fir_filter/n1041 ,
         \u_decoder/fir_filter/n1040 , \u_decoder/fir_filter/n1039 ,
         \u_decoder/fir_filter/n1038 , \u_decoder/fir_filter/n1037 ,
         \u_decoder/fir_filter/n1035 , \u_decoder/fir_filter/n1034 ,
         \u_decoder/fir_filter/n1033 , \u_decoder/fir_filter/n1032 ,
         \u_decoder/fir_filter/n1031 , \u_decoder/fir_filter/n1030 ,
         \u_decoder/fir_filter/n1029 , \u_decoder/fir_filter/n1028 ,
         \u_decoder/fir_filter/n1027 , \u_decoder/fir_filter/n1026 ,
         \u_decoder/fir_filter/n1025 , \u_decoder/fir_filter/n1024 ,
         \u_decoder/fir_filter/n1023 , \u_decoder/fir_filter/n1022 ,
         \u_decoder/fir_filter/n1021 , \u_decoder/fir_filter/n1020 ,
         \u_decoder/fir_filter/n1019 , \u_decoder/fir_filter/n1011 ,
         \u_decoder/fir_filter/n1010 , \u_decoder/fir_filter/n1009 ,
         \u_decoder/fir_filter/n1008 , \u_decoder/fir_filter/n1007 ,
         \u_decoder/fir_filter/n1006 , \u_decoder/fir_filter/n1005 ,
         \u_decoder/fir_filter/n1004 , \u_decoder/fir_filter/n1003 ,
         \u_decoder/fir_filter/n1002 , \u_decoder/fir_filter/n1001 ,
         \u_decoder/fir_filter/n1000 , \u_decoder/fir_filter/n999 ,
         \u_decoder/fir_filter/n998 , \u_decoder/fir_filter/n997 ,
         \u_decoder/fir_filter/n996 , \u_decoder/fir_filter/n995 ,
         \u_decoder/fir_filter/n994 , \u_decoder/fir_filter/n993 ,
         \u_decoder/fir_filter/n992 , \u_decoder/fir_filter/n991 ,
         \u_decoder/fir_filter/n990 , \u_decoder/fir_filter/n989 ,
         \u_decoder/fir_filter/n988 , \u_decoder/fir_filter/n987 ,
         \u_decoder/fir_filter/n986 , \u_decoder/fir_filter/n985 ,
         \u_decoder/fir_filter/n984 , \u_decoder/fir_filter/n983 ,
         \u_decoder/fir_filter/n982 , \u_decoder/fir_filter/n975 ,
         \u_decoder/fir_filter/n974 , \u_decoder/fir_filter/n973 ,
         \u_decoder/fir_filter/n972 , \u_decoder/fir_filter/n971 ,
         \u_decoder/fir_filter/n970 , \u_decoder/fir_filter/n969 ,
         \u_decoder/fir_filter/n968 , \u_decoder/fir_filter/n967 ,
         \u_decoder/fir_filter/n966 , \u_decoder/fir_filter/n965 ,
         \u_decoder/fir_filter/n964 , \u_decoder/fir_filter/n963 ,
         \u_decoder/fir_filter/n962 , \u_decoder/fir_filter/n961 ,
         \u_decoder/fir_filter/n954 , \u_decoder/fir_filter/n953 ,
         \u_decoder/fir_filter/n952 , \u_decoder/fir_filter/n951 ,
         \u_decoder/fir_filter/n950 , \u_decoder/fir_filter/n949 ,
         \u_decoder/fir_filter/n948 , \u_decoder/fir_filter/n947 ,
         \u_decoder/fir_filter/n946 , \u_decoder/fir_filter/n945 ,
         \u_decoder/fir_filter/n944 , \u_decoder/fir_filter/n943 ,
         \u_decoder/fir_filter/n942 , \u_decoder/fir_filter/n941 ,
         \u_decoder/fir_filter/n940 , \u_decoder/fir_filter/n933 ,
         \u_decoder/fir_filter/n932 , \u_decoder/fir_filter/n931 ,
         \u_decoder/fir_filter/n930 , \u_decoder/fir_filter/n929 ,
         \u_decoder/fir_filter/n928 , \u_decoder/fir_filter/n927 ,
         \u_decoder/fir_filter/n926 , \u_decoder/fir_filter/n925 ,
         \u_decoder/fir_filter/n924 , \u_decoder/fir_filter/n923 ,
         \u_decoder/fir_filter/n922 , \u_decoder/fir_filter/n921 ,
         \u_decoder/fir_filter/n920 , \u_decoder/fir_filter/n919 ,
         \u_decoder/fir_filter/n912 , \u_decoder/fir_filter/n911 ,
         \u_decoder/fir_filter/n910 , \u_decoder/fir_filter/n909 ,
         \u_decoder/fir_filter/n908 , \u_decoder/fir_filter/n907 ,
         \u_decoder/fir_filter/n906 , \u_decoder/fir_filter/n905 ,
         \u_decoder/fir_filter/n904 , \u_decoder/fir_filter/n903 ,
         \u_decoder/fir_filter/n902 , \u_decoder/fir_filter/n901 ,
         \u_decoder/fir_filter/n900 , \u_decoder/fir_filter/n899 ,
         \u_decoder/fir_filter/n898 , \u_decoder/fir_filter/n891 ,
         \u_decoder/fir_filter/n890 , \u_decoder/fir_filter/n889 ,
         \u_decoder/fir_filter/n888 , \u_decoder/fir_filter/n887 ,
         \u_decoder/fir_filter/n886 , \u_decoder/fir_filter/n885 ,
         \u_decoder/fir_filter/n884 , \u_decoder/fir_filter/n883 ,
         \u_decoder/fir_filter/n882 , \u_decoder/fir_filter/n881 ,
         \u_decoder/fir_filter/n880 , \u_decoder/fir_filter/n879 ,
         \u_decoder/fir_filter/n878 , \u_decoder/fir_filter/n877 ,
         \u_decoder/fir_filter/n870 , \u_decoder/fir_filter/n869 ,
         \u_decoder/fir_filter/n868 , \u_decoder/fir_filter/n867 ,
         \u_decoder/fir_filter/n866 , \u_decoder/fir_filter/n865 ,
         \u_decoder/fir_filter/n864 , \u_decoder/fir_filter/n863 ,
         \u_decoder/fir_filter/n862 , \u_decoder/fir_filter/n861 ,
         \u_decoder/fir_filter/n860 , \u_decoder/fir_filter/n859 ,
         \u_decoder/fir_filter/n858 , \u_decoder/fir_filter/n857 ,
         \u_decoder/fir_filter/n856 , \u_decoder/fir_filter/n855 ,
         \u_decoder/fir_filter/n854 , \u_decoder/fir_filter/n853 ,
         \u_decoder/fir_filter/n852 , \u_decoder/fir_filter/n851 ,
         \u_decoder/fir_filter/n850 , \u_decoder/fir_filter/n849 ,
         \u_decoder/fir_filter/n848 , \u_decoder/fir_filter/n847 ,
         \u_decoder/fir_filter/n846 , \u_decoder/fir_filter/n845 ,
         \u_decoder/fir_filter/n844 , \u_decoder/fir_filter/n843 ,
         \u_decoder/fir_filter/n842 , \u_decoder/fir_filter/n841 ,
         \u_decoder/fir_filter/n840 , \u_decoder/fir_filter/n839 ,
         \u_decoder/fir_filter/n838 , \u_decoder/fir_filter/n837 ,
         \u_decoder/fir_filter/n835 , \u_decoder/fir_filter/n834 ,
         \u_decoder/fir_filter/n833 , \u_decoder/fir_filter/n832 ,
         \u_decoder/fir_filter/n831 , \u_decoder/fir_filter/n830 ,
         \u_decoder/fir_filter/n829 , \u_decoder/fir_filter/n828 ,
         \u_decoder/fir_filter/n827 , \u_decoder/fir_filter/n826 ,
         \u_decoder/fir_filter/n825 , \u_decoder/fir_filter/n824 ,
         \u_decoder/fir_filter/n823 , \u_decoder/fir_filter/n822 ,
         \u_decoder/fir_filter/n821 , \u_decoder/fir_filter/n819 ,
         \u_decoder/fir_filter/n818 , \u_decoder/fir_filter/n817 ,
         \u_decoder/fir_filter/n816 , \u_decoder/fir_filter/n815 ,
         \u_decoder/fir_filter/n814 , \u_decoder/fir_filter/n813 ,
         \u_decoder/fir_filter/n812 , \u_decoder/fir_filter/n811 ,
         \u_decoder/fir_filter/n810 , \u_decoder/fir_filter/n809 ,
         \u_decoder/fir_filter/n808 , \u_decoder/fir_filter/n807 ,
         \u_decoder/fir_filter/n806 , \u_decoder/fir_filter/n805 ,
         \u_decoder/fir_filter/n803 , \u_decoder/fir_filter/n802 ,
         \u_decoder/fir_filter/n801 , \u_decoder/fir_filter/n800 ,
         \u_decoder/fir_filter/n799 , \u_decoder/fir_filter/n798 ,
         \u_decoder/fir_filter/n797 , \u_decoder/fir_filter/n796 ,
         \u_decoder/fir_filter/n795 , \u_decoder/fir_filter/n794 ,
         \u_decoder/fir_filter/n793 , \u_decoder/fir_filter/n792 ,
         \u_decoder/fir_filter/n791 , \u_decoder/fir_filter/n790 ,
         \u_decoder/fir_filter/n789 , \u_decoder/fir_filter/n787 ,
         \u_decoder/fir_filter/n786 , \u_decoder/fir_filter/n785 ,
         \u_decoder/fir_filter/n784 , \u_decoder/fir_filter/n783 ,
         \u_decoder/fir_filter/n782 , \u_decoder/fir_filter/n781 ,
         \u_decoder/fir_filter/n780 , \u_decoder/fir_filter/n779 ,
         \u_decoder/fir_filter/n778 , \u_decoder/fir_filter/n777 ,
         \u_decoder/fir_filter/n776 , \u_decoder/fir_filter/n775 ,
         \u_decoder/fir_filter/n774 , \u_decoder/fir_filter/n773 ,
         \u_decoder/fir_filter/n771 , \u_decoder/fir_filter/n770 ,
         \u_decoder/fir_filter/n769 , \u_decoder/fir_filter/n768 ,
         \u_decoder/fir_filter/n767 , \u_decoder/fir_filter/n766 ,
         \u_decoder/fir_filter/n765 , \u_decoder/fir_filter/n764 ,
         \u_decoder/fir_filter/n763 , \u_decoder/fir_filter/n762 ,
         \u_decoder/fir_filter/n761 , \u_decoder/fir_filter/n760 ,
         \u_decoder/fir_filter/n759 , \u_decoder/fir_filter/n758 ,
         \u_decoder/fir_filter/n757 , \u_decoder/fir_filter/n755 ,
         \u_decoder/fir_filter/n754 , \u_decoder/fir_filter/n753 ,
         \u_decoder/fir_filter/n752 , \u_decoder/fir_filter/n751 ,
         \u_decoder/fir_filter/n750 , \u_decoder/fir_filter/n749 ,
         \u_decoder/fir_filter/n748 , \u_decoder/fir_filter/n747 ,
         \u_decoder/fir_filter/n746 , \u_decoder/fir_filter/n745 ,
         \u_decoder/fir_filter/n744 , \u_decoder/fir_filter/n743 ,
         \u_decoder/fir_filter/n742 , \u_decoder/fir_filter/n741 ,
         \u_decoder/fir_filter/n740 , \u_decoder/fir_filter/n738 ,
         \u_decoder/fir_filter/n737 , \u_decoder/fir_filter/n736 ,
         \u_decoder/fir_filter/n735 , \u_decoder/fir_filter/n734 ,
         \u_decoder/fir_filter/n733 , \u_decoder/fir_filter/n732 ,
         \u_decoder/fir_filter/n731 , \u_decoder/fir_filter/n730 ,
         \u_decoder/fir_filter/n729 , \u_decoder/fir_filter/n728 ,
         \u_decoder/fir_filter/n727 , \u_decoder/fir_filter/n726 ,
         \u_decoder/fir_filter/n725 , \u_decoder/fir_filter/n724 ,
         \u_decoder/fir_filter/n723 , \u_decoder/fir_filter/n722 ,
         \u_decoder/fir_filter/n721 , \u_decoder/fir_filter/n713 ,
         \u_decoder/fir_filter/n712 , \u_decoder/fir_filter/n711 ,
         \u_decoder/fir_filter/n710 , \u_decoder/fir_filter/n709 ,
         \u_decoder/fir_filter/n708 , \u_decoder/fir_filter/n707 ,
         \u_decoder/fir_filter/n706 , \u_decoder/fir_filter/n705 ,
         \u_decoder/fir_filter/n704 , \u_decoder/fir_filter/n703 ,
         \u_decoder/fir_filter/n702 , \u_decoder/fir_filter/n701 ,
         \u_decoder/fir_filter/n700 , \u_decoder/fir_filter/n699 ,
         \u_decoder/fir_filter/n698 , \u_decoder/fir_filter/n697 ,
         \u_decoder/fir_filter/n696 , \u_decoder/fir_filter/n695 ,
         \u_decoder/fir_filter/n694 , \u_decoder/fir_filter/n693 ,
         \u_decoder/fir_filter/n692 , \u_decoder/fir_filter/n691 ,
         \u_decoder/fir_filter/n690 , \u_decoder/fir_filter/n689 ,
         \u_decoder/fir_filter/n688 , \u_decoder/fir_filter/n687 ,
         \u_decoder/fir_filter/n686 , \u_decoder/fir_filter/n685 ,
         \u_decoder/fir_filter/n684 , \u_decoder/fir_filter/n677 ,
         \u_decoder/fir_filter/n676 , \u_decoder/fir_filter/n675 ,
         \u_decoder/fir_filter/n674 , \u_decoder/fir_filter/n673 ,
         \u_decoder/fir_filter/n672 , \u_decoder/fir_filter/n671 ,
         \u_decoder/fir_filter/n670 , \u_decoder/fir_filter/n669 ,
         \u_decoder/fir_filter/n668 , \u_decoder/fir_filter/n667 ,
         \u_decoder/fir_filter/n666 , \u_decoder/fir_filter/n665 ,
         \u_decoder/fir_filter/n664 , \u_decoder/fir_filter/n663 ,
         \u_decoder/fir_filter/n656 , \u_decoder/fir_filter/n655 ,
         \u_decoder/fir_filter/n654 , \u_decoder/fir_filter/n653 ,
         \u_decoder/fir_filter/n652 , \u_decoder/fir_filter/n651 ,
         \u_decoder/fir_filter/n650 , \u_decoder/fir_filter/n649 ,
         \u_decoder/fir_filter/n648 , \u_decoder/fir_filter/n647 ,
         \u_decoder/fir_filter/n646 , \u_decoder/fir_filter/n645 ,
         \u_decoder/fir_filter/n644 , \u_decoder/fir_filter/n643 ,
         \u_decoder/fir_filter/n642 , \u_decoder/fir_filter/n635 ,
         \u_decoder/fir_filter/n634 , \u_decoder/fir_filter/n633 ,
         \u_decoder/fir_filter/n632 , \u_decoder/fir_filter/n631 ,
         \u_decoder/fir_filter/n630 , \u_decoder/fir_filter/n629 ,
         \u_decoder/fir_filter/n628 , \u_decoder/fir_filter/n627 ,
         \u_decoder/fir_filter/n626 , \u_decoder/fir_filter/n625 ,
         \u_decoder/fir_filter/n624 , \u_decoder/fir_filter/n623 ,
         \u_decoder/fir_filter/n622 , \u_decoder/fir_filter/n621 ,
         \u_decoder/fir_filter/n614 , \u_decoder/fir_filter/n613 ,
         \u_decoder/fir_filter/n612 , \u_decoder/fir_filter/n611 ,
         \u_decoder/fir_filter/n610 , \u_decoder/fir_filter/n609 ,
         \u_decoder/fir_filter/n608 , \u_decoder/fir_filter/n607 ,
         \u_decoder/fir_filter/n606 , \u_decoder/fir_filter/n605 ,
         \u_decoder/fir_filter/n604 , \u_decoder/fir_filter/n603 ,
         \u_decoder/fir_filter/n602 , \u_decoder/fir_filter/n601 ,
         \u_decoder/fir_filter/n600 , \u_decoder/fir_filter/n593 ,
         \u_decoder/fir_filter/n592 , \u_decoder/fir_filter/n591 ,
         \u_decoder/fir_filter/n590 , \u_decoder/fir_filter/n589 ,
         \u_decoder/fir_filter/n588 , \u_decoder/fir_filter/n587 ,
         \u_decoder/fir_filter/n586 , \u_decoder/fir_filter/n585 ,
         \u_decoder/fir_filter/n584 , \u_decoder/fir_filter/n583 ,
         \u_decoder/fir_filter/n582 , \u_decoder/fir_filter/n581 ,
         \u_decoder/fir_filter/n580 , \u_decoder/fir_filter/n579 ,
         \u_decoder/fir_filter/n572 , \u_decoder/fir_filter/n571 ,
         \u_decoder/fir_filter/n570 , \u_decoder/fir_filter/n569 ,
         \u_decoder/fir_filter/n568 , \u_decoder/fir_filter/n567 ,
         \u_decoder/fir_filter/n566 , \u_decoder/fir_filter/n565 ,
         \u_decoder/fir_filter/n564 , \u_decoder/fir_filter/n563 ,
         \u_decoder/fir_filter/n562 , \u_decoder/fir_filter/n561 ,
         \u_decoder/fir_filter/n560 , \u_decoder/fir_filter/n559 ,
         \u_decoder/fir_filter/n558 , \u_decoder/fir_filter/n557 ,
         \u_decoder/fir_filter/n556 , \u_decoder/fir_filter/n555 ,
         \u_decoder/fir_filter/n554 , \u_decoder/fir_filter/n553 ,
         \u_decoder/fir_filter/n442 , \u_decoder/fir_filter/n441 ,
         \u_decoder/fir_filter/n440 , \u_decoder/fir_filter/n439 ,
         \u_decoder/fir_filter/n438 , \u_decoder/fir_filter/n437 ,
         \u_decoder/fir_filter/n436 , \u_decoder/fir_filter/n435 ,
         \u_decoder/fir_filter/n434 , \u_decoder/fir_filter/n433 ,
         \u_decoder/fir_filter/n432 , \u_decoder/fir_filter/n431 ,
         \u_decoder/fir_filter/n430 , \u_decoder/fir_filter/n429 ,
         \u_decoder/fir_filter/n428 , \u_decoder/fir_filter/n426 ,
         \u_decoder/fir_filter/n425 , \u_decoder/fir_filter/n424 ,
         \u_decoder/fir_filter/n423 , \u_decoder/fir_filter/n422 ,
         \u_decoder/fir_filter/n421 , \u_decoder/fir_filter/n420 ,
         \u_decoder/fir_filter/n419 , \u_decoder/fir_filter/n418 ,
         \u_decoder/fir_filter/n417 , \u_decoder/fir_filter/n416 ,
         \u_decoder/fir_filter/n415 , \u_decoder/fir_filter/n414 ,
         \u_decoder/fir_filter/n413 , \u_decoder/fir_filter/n412 ,
         \u_decoder/fir_filter/n410 , \u_decoder/fir_filter/Q_data_mult_2[8] ,
         \u_decoder/fir_filter/Q_data_mult_2_15 ,
         \u_decoder/fir_filter/Q_data_mult_1[4] ,
         \u_decoder/fir_filter/Q_data_mult_1_15 ,
         \u_decoder/fir_filter/Q_data_mult_0_15 ,
         \u_decoder/fir_filter/I_data_mult_2[8] ,
         \u_decoder/fir_filter/I_data_mult_2_15 ,
         \u_decoder/fir_filter/I_data_mult_1[4] ,
         \u_decoder/fir_filter/I_data_mult_1_15 ,
         \u_decoder/fir_filter/I_data_mult_0_15 , \u_decoder/fir_filter/N12 ,
         \u_decoder/fir_filter/N11 , \u_cordic/mycordic/n586 ,
         \u_cordic/mycordic/n585 , \u_cordic/mycordic/n584 ,
         \u_cordic/mycordic/n583 , \u_cordic/mycordic/n582 ,
         \u_cordic/mycordic/n581 , \u_cordic/mycordic/n580 ,
         \u_cordic/mycordic/n579 , \u_cordic/mycordic/n578 ,
         \u_cordic/mycordic/n577 , \u_cordic/mycordic/n576 ,
         \u_cordic/mycordic/n575 , \u_cordic/mycordic/n574 ,
         \u_cordic/mycordic/n573 , \u_cordic/mycordic/n572 ,
         \u_cordic/mycordic/n571 , \u_cordic/mycordic/n570 ,
         \u_cordic/mycordic/n569 , \u_cordic/mycordic/n568 ,
         \u_cordic/mycordic/n567 , \u_cordic/mycordic/n566 ,
         \u_cordic/mycordic/n565 , \u_cordic/mycordic/n564 ,
         \u_cordic/mycordic/n563 , \u_cordic/mycordic/n562 ,
         \u_cordic/mycordic/n561 , \u_cordic/mycordic/n560 ,
         \u_cordic/mycordic/n559 , \u_cordic/mycordic/n558 ,
         \u_cordic/mycordic/n557 , \u_cordic/mycordic/n556 ,
         \u_cordic/mycordic/n555 , \u_cordic/mycordic/n554 ,
         \u_cordic/mycordic/n553 , \u_cordic/mycordic/n552 ,
         \u_cordic/mycordic/n551 , \u_cordic/mycordic/n550 ,
         \u_cordic/mycordic/n549 , \u_cordic/mycordic/n548 ,
         \u_cordic/mycordic/n547 , \u_cordic/mycordic/n546 ,
         \u_cordic/mycordic/n545 , \u_cordic/mycordic/n544 ,
         \u_cordic/mycordic/n543 , \u_cordic/mycordic/n542 ,
         \u_cordic/mycordic/n541 , \u_cordic/mycordic/n540 ,
         \u_cordic/mycordic/n539 , \u_cordic/mycordic/n538 ,
         \u_cordic/mycordic/n537 , \u_cordic/mycordic/n536 ,
         \u_cordic/mycordic/n520 , \u_cordic/mycordic/n519 ,
         \u_cordic/mycordic/n518 , \u_cordic/mycordic/n517 ,
         \u_cordic/mycordic/n516 , \u_cordic/mycordic/n515 ,
         \u_cordic/mycordic/n514 , \u_cordic/mycordic/n513 ,
         \u_cordic/mycordic/n512 , \u_cordic/mycordic/n511 ,
         \u_cordic/mycordic/n510 , \u_cordic/mycordic/n509 ,
         \u_cordic/mycordic/n508 , \u_cordic/mycordic/n507 ,
         \u_cordic/mycordic/n506 , \u_cordic/mycordic/n505 ,
         \u_cordic/mycordic/n504 , \u_cordic/mycordic/n503 ,
         \u_cordic/mycordic/n502 , \u_cordic/mycordic/n501 ,
         \u_cordic/mycordic/n500 , \u_cordic/mycordic/n499 ,
         \u_cordic/mycordic/n498 , \u_cordic/mycordic/n497 ,
         \u_cordic/mycordic/n496 , \u_cordic/mycordic/n495 ,
         \u_cordic/mycordic/n494 , \u_cordic/mycordic/n493 ,
         \u_cordic/mycordic/n492 , \u_cordic/mycordic/n491 ,
         \u_cordic/mycordic/n490 , \u_cordic/mycordic/n489 ,
         \u_cordic/mycordic/n488 , \u_cordic/mycordic/n487 ,
         \u_cordic/mycordic/n486 , \u_cordic/mycordic/n485 ,
         \u_cordic/mycordic/n484 , \u_cordic/mycordic/n483 ,
         \u_cordic/mycordic/n482 , \u_cordic/mycordic/n481 ,
         \u_cordic/mycordic/n480 , \u_cordic/mycordic/n479 ,
         \u_cordic/mycordic/n478 , \u_cordic/mycordic/n477 ,
         \u_cordic/mycordic/n476 , \u_cordic/mycordic/n475 ,
         \u_cordic/mycordic/n474 , \u_cordic/mycordic/n473 ,
         \u_cordic/mycordic/n472 , \u_cordic/mycordic/n471 ,
         \u_cordic/mycordic/n470 , \u_cordic/mycordic/n469 ,
         \u_cordic/mycordic/n468 , \u_cordic/mycordic/n467 ,
         \u_cordic/mycordic/n466 , \u_cordic/mycordic/n465 ,
         \u_cordic/mycordic/n464 , \u_cordic/mycordic/n463 ,
         \u_cordic/mycordic/n462 , \u_cordic/mycordic/n461 ,
         \u_cordic/mycordic/n460 , \u_cordic/mycordic/n459 ,
         \u_cordic/mycordic/n458 , \u_cordic/mycordic/n457 ,
         \u_cordic/mycordic/n456 , \u_cordic/mycordic/n455 ,
         \u_cordic/mycordic/n454 , \u_cordic/mycordic/n453 ,
         \u_cordic/mycordic/n452 , \u_cordic/mycordic/n451 ,
         \u_cordic/mycordic/n450 , \u_cordic/mycordic/n449 ,
         \u_cordic/mycordic/n448 , \u_cordic/mycordic/n447 ,
         \u_cordic/mycordic/n446 , \u_cordic/mycordic/n445 ,
         \u_cordic/mycordic/n444 , \u_cordic/mycordic/n443 ,
         \u_cordic/mycordic/n442 , \u_cordic/mycordic/n441 ,
         \u_cordic/mycordic/n440 , \u_cordic/mycordic/n439 ,
         \u_cordic/mycordic/n438 , \u_cordic/mycordic/n437 ,
         \u_cordic/mycordic/n436 , \u_cordic/mycordic/n435 ,
         \u_cordic/mycordic/n433 , \u_cordic/mycordic/n432 ,
         \u_cordic/mycordic/n431 , \u_cordic/mycordic/n430 ,
         \u_cordic/mycordic/n429 , \u_cordic/mycordic/n428 ,
         \u_cordic/mycordic/n427 , \u_cordic/mycordic/n426 ,
         \u_cordic/mycordic/n425 , \u_cordic/mycordic/n424 ,
         \u_cordic/mycordic/n423 , \u_cordic/mycordic/n422 ,
         \u_cordic/mycordic/n421 , \u_cordic/mycordic/n420 ,
         \u_cordic/mycordic/n419 , \u_cordic/mycordic/n418 ,
         \u_cordic/mycordic/n417 , \u_cordic/mycordic/n416 ,
         \u_cordic/mycordic/n415 , \u_cordic/mycordic/n414 ,
         \u_cordic/mycordic/n413 , \u_cordic/mycordic/n412 ,
         \u_cordic/mycordic/n411 , \u_cordic/mycordic/n410 ,
         \u_cordic/mycordic/n409 , \u_cordic/mycordic/n408 ,
         \u_cordic/mycordic/n407 , \u_cordic/mycordic/n406 ,
         \u_cordic/mycordic/n405 , \u_cordic/mycordic/n404 ,
         \u_cordic/mycordic/n403 , \u_cordic/mycordic/n402 ,
         \u_cordic/mycordic/n401 , \u_cordic/mycordic/n400 ,
         \u_cordic/mycordic/n399 , \u_cordic/mycordic/n395 ,
         \u_cordic/mycordic/n394 , \u_cordic/mycordic/n393 ,
         \u_cordic/mycordic/n392 , \u_cordic/mycordic/n391 ,
         \u_cordic/mycordic/n387 , \u_cordic/mycordic/n386 ,
         \u_cordic/mycordic/n385 , \u_cordic/mycordic/n384 ,
         \u_cordic/mycordic/n383 , \u_cordic/mycordic/n382 ,
         \u_cordic/mycordic/n381 , \u_cordic/mycordic/n380 ,
         \u_cordic/mycordic/n379 , \u_cordic/mycordic/n378 ,
         \u_cordic/mycordic/n377 , \u_cordic/mycordic/n376 ,
         \u_cordic/mycordic/n375 , \u_cordic/mycordic/n374 ,
         \u_cordic/mycordic/n373 , \u_cordic/mycordic/n372 ,
         \u_cordic/mycordic/n371 , \u_cordic/mycordic/n370 ,
         \u_cordic/mycordic/n369 , \u_cordic/mycordic/n368 ,
         \u_cordic/mycordic/n367 , \u_cordic/mycordic/n366 ,
         \u_cordic/mycordic/n365 , \u_cordic/mycordic/n364 ,
         \u_cordic/mycordic/n363 , \u_cordic/mycordic/n362 ,
         \u_cordic/mycordic/n358 , \u_cordic/mycordic/n357 ,
         \u_cordic/mycordic/n356 , \u_cordic/mycordic/n355 ,
         \u_cordic/mycordic/n354 , \u_cordic/mycordic/n353 ,
         \u_cordic/mycordic/n349 , \u_cordic/mycordic/n348 ,
         \u_cordic/mycordic/n347 , \u_cordic/mycordic/n346 ,
         \u_cordic/mycordic/n345 , \u_cordic/mycordic/n344 ,
         \u_cordic/mycordic/n343 , \u_cordic/mycordic/n342 ,
         \u_cordic/mycordic/n341 , \u_cordic/mycordic/n340 ,
         \u_cordic/mycordic/n339 , \u_cordic/mycordic/n338 ,
         \u_cordic/mycordic/n337 , \u_cordic/mycordic/n336 ,
         \u_cordic/mycordic/n335 , \u_cordic/mycordic/n334 ,
         \u_cordic/mycordic/n333 , \u_cordic/mycordic/n332 ,
         \u_cordic/mycordic/n331 , \u_cordic/mycordic/n110 ,
         \u_cordic/mycordic/n108 , \u_cordic/mycordic/N630 ,
         \u_cordic/mycordic/N629 , \u_cordic/mycordic/N628 ,
         \u_cordic/mycordic/N627 , \u_cordic/mycordic/N626 ,
         \u_cordic/mycordic/N625 , \u_cordic/mycordic/N624 ,
         \u_cordic/mycordic/N623 , \u_cordic/mycordic/N622 ,
         \u_cordic/mycordic/N621 , \u_cordic/mycordic/N620 ,
         \u_cordic/mycordic/N619 , \u_cordic/mycordic/N615 ,
         \u_cordic/mycordic/N565 , \u_cordic/mycordic/N564 ,
         \u_cordic/mycordic/N563 , \u_cordic/mycordic/N562 ,
         \u_cordic/mycordic/N561 , \u_cordic/mycordic/N560 ,
         \u_cordic/mycordic/N559 , \u_cordic/mycordic/N558 ,
         \u_cordic/mycordic/N557 , \u_cordic/mycordic/N556 ,
         \u_cordic/mycordic/N555 , \u_cordic/mycordic/N554 ,
         \u_cordic/mycordic/N553 , \u_cordic/mycordic/N552 ,
         \u_cordic/mycordic/N550 , \u_cordic/mycordic/N549 ,
         \u_cordic/mycordic/N548 , \u_cordic/mycordic/N547 ,
         \u_cordic/mycordic/N546 , \u_cordic/mycordic/N545 ,
         \u_cordic/mycordic/N544 , \u_cordic/mycordic/N543 ,
         \u_cordic/mycordic/N542 , \u_cordic/mycordic/N541 ,
         \u_cordic/mycordic/N540 , \u_cordic/mycordic/N539 ,
         \u_cordic/mycordic/N538 , \u_cordic/mycordic/N537 ,
         \u_cordic/mycordic/N536 , \u_cordic/mycordic/N533 ,
         \u_cordic/mycordic/N532 , \u_cordic/mycordic/N531 ,
         \u_cordic/mycordic/N530 , \u_cordic/mycordic/N529 ,
         \u_cordic/mycordic/N528 , \u_cordic/mycordic/N527 ,
         \u_cordic/mycordic/N526 , \u_cordic/mycordic/N525 ,
         \u_cordic/mycordic/N524 , \u_cordic/mycordic/N523 ,
         \u_cordic/mycordic/N522 , \u_cordic/mycordic/N521 ,
         \u_cordic/mycordic/N520 , \u_cordic/mycordic/N519 ,
         \u_cordic/mycordic/N517 , \u_cordic/mycordic/N516 ,
         \u_cordic/mycordic/N515 , \u_cordic/mycordic/N514 ,
         \u_cordic/mycordic/N513 , \u_cordic/mycordic/N512 ,
         \u_cordic/mycordic/N511 , \u_cordic/mycordic/N510 ,
         \u_cordic/mycordic/N509 , \u_cordic/mycordic/N508 ,
         \u_cordic/mycordic/N507 , \u_cordic/mycordic/N506 ,
         \u_cordic/mycordic/N505 , \u_cordic/mycordic/N504 ,
         \u_cordic/mycordic/N503 , \u_cordic/mycordic/N502 ,
         \u_cordic/mycordic/N500 , \u_cordic/mycordic/N499 ,
         \u_cordic/mycordic/N498 , \u_cordic/mycordic/N497 ,
         \u_cordic/mycordic/N496 , \u_cordic/mycordic/N495 ,
         \u_cordic/mycordic/N494 , \u_cordic/mycordic/N493 ,
         \u_cordic/mycordic/N492 , \u_cordic/mycordic/N491 ,
         \u_cordic/mycordic/N490 , \u_cordic/mycordic/N489 ,
         \u_cordic/mycordic/N488 , \u_cordic/mycordic/N487 ,
         \u_cordic/mycordic/N486 , \u_cordic/mycordic/N485 ,
         \u_cordic/mycordic/N483 , \u_cordic/mycordic/N482 ,
         \u_cordic/mycordic/N481 , \u_cordic/mycordic/N480 ,
         \u_cordic/mycordic/N479 , \u_cordic/mycordic/N478 ,
         \u_cordic/mycordic/N477 , \u_cordic/mycordic/N476 ,
         \u_cordic/mycordic/N475 , \u_cordic/mycordic/N474 ,
         \u_cordic/mycordic/N473 , \u_cordic/mycordic/N472 ,
         \u_cordic/mycordic/N471 , \u_cordic/mycordic/N470 ,
         \u_cordic/mycordic/N469 , \u_cordic/mycordic/N468 ,
         \u_cordic/mycordic/N467 , \u_cordic/mycordic/N466 ,
         \u_cordic/mycordic/N465 , \u_cordic/mycordic/N464 ,
         \u_cordic/mycordic/N463 , \u_cordic/mycordic/N462 ,
         \u_cordic/mycordic/N461 , \u_cordic/mycordic/N460 ,
         \u_cordic/mycordic/N459 , \u_cordic/mycordic/N458 ,
         \u_cordic/mycordic/N457 , \u_cordic/mycordic/N455 ,
         \u_cordic/mycordic/N454 , \u_cordic/mycordic/N453 ,
         \u_cordic/mycordic/N452 , \u_cordic/mycordic/N451 ,
         \u_cordic/mycordic/N450 , \u_cordic/mycordic/N449 ,
         \u_cordic/mycordic/N448 , \u_cordic/mycordic/N447 ,
         \u_cordic/mycordic/N446 , \u_cordic/mycordic/N445 ,
         \u_cordic/mycordic/N444 , \u_cordic/mycordic/N443 ,
         \u_cordic/mycordic/N442 , \u_cordic/mycordic/N441 ,
         \u_cordic/mycordic/N440 , \u_cordic/mycordic/N439 ,
         \u_cordic/mycordic/N438 , \u_cordic/mycordic/N437 ,
         \u_cordic/mycordic/N436 , \u_cordic/mycordic/N435 ,
         \u_cordic/mycordic/N434 , \u_cordic/mycordic/N433 ,
         \u_cordic/mycordic/N432 , \u_cordic/mycordic/N431 ,
         \u_cordic/mycordic/N430 , \u_cordic/mycordic/N428 ,
         \u_cordic/mycordic/N427 , \u_cordic/mycordic/N426 ,
         \u_cordic/mycordic/N425 , \u_cordic/mycordic/N424 ,
         \u_cordic/mycordic/N423 , \u_cordic/mycordic/N422 ,
         \u_cordic/mycordic/N421 , \u_cordic/mycordic/N420 ,
         \u_cordic/mycordic/N419 , \u_cordic/mycordic/N418 ,
         \u_cordic/mycordic/N417 , \u_cordic/mycordic/N416 ,
         \u_cordic/mycordic/N415 , \u_cordic/mycordic/N414 ,
         \u_cordic/mycordic/N413 , \u_cordic/mycordic/N412 ,
         \u_cordic/mycordic/N411 , \u_cordic/mycordic/N410 ,
         \u_cordic/mycordic/N409 , \u_cordic/mycordic/N408 ,
         \u_cordic/mycordic/N407 , \u_cordic/mycordic/N406 ,
         \u_cordic/mycordic/N405 , \u_cordic/mycordic/N404 ,
         \u_cordic/mycordic/N403 , \u_cordic/mycordic/N402 ,
         \u_cordic/mycordic/N401 , \u_cordic/mycordic/N400 ,
         \u_cordic/mycordic/N399 , \u_cordic/mycordic/N398 ,
         \u_cordic/mycordic/N395 , \u_cordic/mycordic/N394 ,
         \u_cordic/mycordic/N393 , \u_cordic/mycordic/N392 ,
         \u_cordic/mycordic/N391 , \u_cordic/mycordic/N390 ,
         \u_cordic/mycordic/N389 , \u_cordic/mycordic/N388 ,
         \u_cordic/mycordic/N387 , \u_cordic/mycordic/N386 ,
         \u_cordic/mycordic/N385 , \u_cordic/mycordic/N384 ,
         \u_cordic/mycordic/N383 , \u_cordic/mycordic/N382 ,
         \u_cordic/mycordic/N381 , \u_cordic/mycordic/N380 ,
         \u_cordic/mycordic/N379 , \u_cordic/mycordic/N378 ,
         \u_cordic/mycordic/N377 , \u_cordic/mycordic/N376 ,
         \u_cordic/mycordic/N375 , \u_cordic/mycordic/N374 ,
         \u_cordic/mycordic/N373 , \u_cordic/mycordic/N372 ,
         \u_cordic/mycordic/N371 , \u_cordic/mycordic/N370 ,
         \u_cordic/mycordic/N369 , \u_cordic/mycordic/N368 ,
         \u_cordic/mycordic/N367 , \u_cordic/mycordic/N366 ,
         \u_cordic/mycordic/N365 , \u_cordic/mycordic/N363 ,
         \u_cordic/mycordic/N362 , \u_cordic/mycordic/N361 ,
         \u_cordic/mycordic/N360 , \u_cordic/mycordic/N359 ,
         \u_cordic/mycordic/N358 , \u_cordic/mycordic/N357 ,
         \u_cordic/mycordic/N356 , \u_cordic/mycordic/N355 ,
         \u_cordic/mycordic/N354 , \u_cordic/mycordic/N353 ,
         \u_cordic/mycordic/N352 , \u_cordic/mycordic/N351 ,
         \u_cordic/mycordic/N350 , \u_cordic/mycordic/N349 ,
         \u_cordic/mycordic/N348 , \u_cordic/mycordic/N347 ,
         \u_cordic/mycordic/N346 , \u_cordic/mycordic/N345 ,
         \u_cordic/mycordic/N344 , \u_cordic/mycordic/N343 ,
         \u_cordic/mycordic/N342 , \u_cordic/mycordic/N341 ,
         \u_cordic/mycordic/N340 , \u_cordic/mycordic/N339 ,
         \u_cordic/mycordic/N338 , \u_cordic/mycordic/N337 ,
         \u_cordic/mycordic/N336 , \u_cordic/mycordic/N335 ,
         \u_cordic/mycordic/N334 , \u_cordic/mycordic/N333 ,
         \u_cordic/mycordic/N331 , \u_cordic/mycordic/N330 ,
         \u_cordic/mycordic/N329 , \u_cordic/mycordic/N328 ,
         \u_cordic/mycordic/N327 , \u_cordic/mycordic/N326 ,
         \u_cordic/mycordic/N325 , \u_cordic/mycordic/N324 ,
         \u_cordic/mycordic/N323 , \u_cordic/mycordic/N322 ,
         \u_cordic/mycordic/N321 , \u_cordic/mycordic/N320 ,
         \u_cordic/mycordic/N319 , \u_cordic/mycordic/N318 ,
         \u_cordic/mycordic/N317 , \u_cordic/mycordic/N316 ,
         \u_cordic/mycordic/N291 , \u_cordic/mycordic/N290 ,
         \u_cordic/mycordic/N289 , \u_cordic/mycordic/N288 ,
         \u_cordic/mycordic/N287 , \u_cordic/mycordic/N267 ,
         \u_cordic/mycordic/N266 , \u_cordic/mycordic/N265 ,
         \u_cordic/mycordic/N264 , \u_cordic/mycordic/N263 ,
         \u_cordic/mycordic/N259 , \u_cordic/mycordic/N258 ,
         \u_cordic/mycordic/N257 , \u_cordic/mycordic/N256 ,
         \u_cordic/mycordic/N255 , \u_cordic/mycordic/N247 ,
         \u_cordic/mycordic/N246 , \u_cordic/mycordic/N245 ,
         \u_cordic/mycordic/N244 , \u_cordic/mycordic/N238 ,
         \u_cordic/mycordic/N237 , \u_cordic/mycordic/N236 ,
         \u_cordic/mycordic/N212 , \u_cordic/mycordic/N211 ,
         \u_cordic/mycordic/N44 , \u_cordic/mycordic/next_ANGLE_table[6][15] ,
         \u_cordic/mycordic/next_ANGLE_table[6][14] ,
         \u_cordic/mycordic/next_ANGLE_table[6][13] ,
         \u_cordic/mycordic/next_ANGLE_table[6][12] ,
         \u_cordic/mycordic/next_ANGLE_table[6][11] ,
         \u_cordic/mycordic/next_ANGLE_table[6][10] ,
         \u_cordic/mycordic/next_ANGLE_table[6][9] ,
         \u_cordic/mycordic/next_ANGLE_table[6][8] ,
         \u_cordic/mycordic/next_ANGLE_table[6][7] ,
         \u_cordic/mycordic/next_ANGLE_table[6][6] ,
         \u_cordic/mycordic/next_ANGLE_table[6][5] ,
         \u_cordic/mycordic/next_ANGLE_table[6][4] ,
         \u_cordic/mycordic/next_ANGLE_table[6][3] ,
         \u_cordic/mycordic/next_ANGLE_table[6][2] ,
         \u_cordic/mycordic/next_ANGLE_table[6][1] ,
         \u_cordic/mycordic/next_ANGLE_table[6][0] ,
         \u_cordic/mycordic/present_C_table[1][0] ,
         \u_cordic/mycordic/present_C_table[1][1] ,
         \u_cordic/mycordic/present_C_table[1][2] ,
         \u_cordic/mycordic/present_C_table[2][0] ,
         \u_cordic/mycordic/present_C_table[2][1] ,
         \u_cordic/mycordic/present_C_table[2][2] ,
         \u_cordic/mycordic/present_C_table[3][0] ,
         \u_cordic/mycordic/present_C_table[3][1] ,
         \u_cordic/mycordic/present_C_table[3][2] ,
         \u_cordic/mycordic/present_C_table[4][0] ,
         \u_cordic/mycordic/present_C_table[4][1] ,
         \u_cordic/mycordic/present_C_table[4][2] ,
         \u_cordic/mycordic/present_C_table[5][0] ,
         \u_cordic/mycordic/present_C_table[5][1] ,
         \u_cordic/mycordic/present_C_table[5][2] ,
         \u_cordic/mycordic/present_C_table[6][0] ,
         \u_cordic/mycordic/present_C_table[6][1] ,
         \u_cordic/mycordic/present_C_table[6][2] ,
         \u_cordic/mycordic/present_C_table[7][0] ,
         \u_cordic/mycordic/present_C_table[7][1] ,
         \u_cordic/mycordic/present_ANGLE_table[6][15] ,
         \u_cordic/mycordic/present_ANGLE_table[6][14] ,
         \u_cordic/mycordic/present_ANGLE_table[6][13] ,
         \u_cordic/mycordic/present_ANGLE_table[6][12] ,
         \u_cordic/mycordic/present_ANGLE_table[6][11] ,
         \u_cordic/mycordic/present_ANGLE_table[6][10] ,
         \u_cordic/mycordic/present_ANGLE_table[6][9] ,
         \u_cordic/mycordic/present_ANGLE_table[6][8] ,
         \u_cordic/mycordic/present_ANGLE_table[6][7] ,
         \u_cordic/mycordic/present_ANGLE_table[6][6] ,
         \u_cordic/mycordic/present_ANGLE_table[6][5] ,
         \u_cordic/mycordic/present_ANGLE_table[6][4] ,
         \u_cordic/mycordic/present_ANGLE_table[6][3] ,
         \u_cordic/mycordic/present_ANGLE_table[6][2] ,
         \u_cordic/mycordic/present_ANGLE_table[6][1] ,
         \u_cordic/mycordic/present_ANGLE_table[5][15] ,
         \u_cordic/mycordic/present_ANGLE_table[5][14] ,
         \u_cordic/mycordic/present_ANGLE_table[5][13] ,
         \u_cordic/mycordic/present_ANGLE_table[5][12] ,
         \u_cordic/mycordic/present_ANGLE_table[5][11] ,
         \u_cordic/mycordic/present_ANGLE_table[5][10] ,
         \u_cordic/mycordic/present_ANGLE_table[5][9] ,
         \u_cordic/mycordic/present_ANGLE_table[5][8] ,
         \u_cordic/mycordic/present_ANGLE_table[5][7] ,
         \u_cordic/mycordic/present_ANGLE_table[5][6] ,
         \u_cordic/mycordic/present_ANGLE_table[5][5] ,
         \u_cordic/mycordic/present_ANGLE_table[5][4] ,
         \u_cordic/mycordic/present_ANGLE_table[5][3] ,
         \u_cordic/mycordic/present_ANGLE_table[5][2] ,
         \u_cordic/mycordic/present_ANGLE_table[5][1] ,
         \u_cordic/mycordic/present_ANGLE_table[4][15] ,
         \u_cordic/mycordic/present_ANGLE_table[4][14] ,
         \u_cordic/mycordic/present_ANGLE_table[4][13] ,
         \u_cordic/mycordic/present_ANGLE_table[4][12] ,
         \u_cordic/mycordic/present_ANGLE_table[4][11] ,
         \u_cordic/mycordic/present_ANGLE_table[4][10] ,
         \u_cordic/mycordic/present_ANGLE_table[4][9] ,
         \u_cordic/mycordic/present_ANGLE_table[4][8] ,
         \u_cordic/mycordic/present_ANGLE_table[4][7] ,
         \u_cordic/mycordic/present_ANGLE_table[4][6] ,
         \u_cordic/mycordic/present_ANGLE_table[4][5] ,
         \u_cordic/mycordic/present_ANGLE_table[4][4] ,
         \u_cordic/mycordic/present_ANGLE_table[4][3] ,
         \u_cordic/mycordic/present_ANGLE_table[4][2] ,
         \u_cordic/mycordic/present_ANGLE_table[4][1] ,
         \u_cordic/mycordic/present_ANGLE_table[4][0] ,
         \u_cordic/mycordic/present_ANGLE_table[3][15] ,
         \u_cordic/mycordic/present_ANGLE_table[3][14] ,
         \u_cordic/mycordic/present_ANGLE_table[3][13] ,
         \u_cordic/mycordic/present_ANGLE_table[3][12] ,
         \u_cordic/mycordic/present_ANGLE_table[3][11] ,
         \u_cordic/mycordic/present_ANGLE_table[3][10] ,
         \u_cordic/mycordic/present_ANGLE_table[3][9] ,
         \u_cordic/mycordic/present_ANGLE_table[3][8] ,
         \u_cordic/mycordic/present_ANGLE_table[3][7] ,
         \u_cordic/mycordic/present_ANGLE_table[3][6] ,
         \u_cordic/mycordic/present_ANGLE_table[3][5] ,
         \u_cordic/mycordic/present_ANGLE_table[3][4] ,
         \u_cordic/mycordic/present_ANGLE_table[3][3] ,
         \u_cordic/mycordic/present_ANGLE_table[3][2] ,
         \u_cordic/mycordic/present_ANGLE_table[3][1] ,
         \u_cordic/mycordic/present_ANGLE_table[3][0] ,
         \u_cordic/mycordic/present_ANGLE_table[2][15] ,
         \u_cordic/mycordic/present_ANGLE_table[2][14] ,
         \u_cordic/mycordic/present_ANGLE_table[2][13] ,
         \u_cordic/mycordic/present_ANGLE_table[2][12] ,
         \u_cordic/mycordic/present_ANGLE_table[2][11] ,
         \u_cordic/mycordic/present_ANGLE_table[2][10] ,
         \u_cordic/mycordic/present_ANGLE_table[2][9] ,
         \u_cordic/mycordic/present_ANGLE_table[2][8] ,
         \u_cordic/mycordic/present_ANGLE_table[2][7] ,
         \u_cordic/mycordic/present_ANGLE_table[2][6] ,
         \u_cordic/mycordic/present_ANGLE_table[2][5] ,
         \u_cordic/mycordic/present_ANGLE_table[2][4] ,
         \u_cordic/mycordic/present_ANGLE_table[2][3] ,
         \u_cordic/mycordic/present_ANGLE_table[2][2] ,
         \u_cordic/mycordic/present_ANGLE_table[2][1] ,
         \u_cordic/mycordic/present_ANGLE_table[1][15] ,
         \u_cordic/mycordic/present_ANGLE_table[1][14] ,
         \u_cordic/mycordic/present_ANGLE_table[1][13] ,
         \u_cordic/mycordic/present_ANGLE_table[1][12] ,
         \u_cordic/mycordic/present_ANGLE_table[1][11] ,
         \u_cordic/mycordic/present_ANGLE_table[1][10] ,
         \u_cordic/mycordic/present_ANGLE_table[1][9] ,
         \u_cordic/mycordic/present_ANGLE_table[1][8] ,
         \u_cordic/mycordic/present_ANGLE_table[1][7] ,
         \u_cordic/mycordic/present_ANGLE_table[1][6] ,
         \u_cordic/mycordic/present_ANGLE_table[1][5] ,
         \u_cordic/mycordic/present_ANGLE_table[1][4] ,
         \u_cordic/mycordic/present_ANGLE_table[1][3] ,
         \u_cordic/mycordic/present_ANGLE_table[1][2] ,
         \u_cordic/mycordic/present_ANGLE_table[1][1] ,
         \u_cordic/mycordic/present_ANGLE_table[1][0] ,
         \u_cordic/mycordic/present_Q_table[0][3] ,
         \u_cordic/mycordic/present_Q_table[0][4] ,
         \u_cordic/mycordic/present_Q_table[0][5] ,
         \u_cordic/mycordic/present_Q_table[0][6] ,
         \u_cordic/mycordic/present_Q_table[0][7] ,
         \u_cordic/mycordic/present_Q_table[1][3] ,
         \u_cordic/mycordic/present_Q_table[1][4] ,
         \u_cordic/mycordic/present_Q_table[1][5] ,
         \u_cordic/mycordic/present_Q_table[1][6] ,
         \u_cordic/mycordic/present_Q_table[1][7] ,
         \u_cordic/mycordic/present_Q_table[2][0] ,
         \u_cordic/mycordic/present_Q_table[2][1] ,
         \u_cordic/mycordic/present_Q_table[2][2] ,
         \u_cordic/mycordic/present_Q_table[2][3] ,
         \u_cordic/mycordic/present_Q_table[2][4] ,
         \u_cordic/mycordic/present_Q_table[2][5] ,
         \u_cordic/mycordic/present_Q_table[2][6] ,
         \u_cordic/mycordic/present_Q_table[2][7] ,
         \u_cordic/mycordic/present_Q_table[3][0] ,
         \u_cordic/mycordic/present_Q_table[3][1] ,
         \u_cordic/mycordic/present_Q_table[3][2] ,
         \u_cordic/mycordic/present_Q_table[3][3] ,
         \u_cordic/mycordic/present_Q_table[3][4] ,
         \u_cordic/mycordic/present_Q_table[3][5] ,
         \u_cordic/mycordic/present_Q_table[3][6] ,
         \u_cordic/mycordic/present_Q_table[3][7] ,
         \u_cordic/mycordic/present_Q_table[4][0] ,
         \u_cordic/mycordic/present_Q_table[4][1] ,
         \u_cordic/mycordic/present_Q_table[4][2] ,
         \u_cordic/mycordic/present_Q_table[4][3] ,
         \u_cordic/mycordic/present_Q_table[4][4] ,
         \u_cordic/mycordic/present_Q_table[4][5] ,
         \u_cordic/mycordic/present_Q_table[4][6] ,
         \u_cordic/mycordic/present_Q_table[4][7] ,
         \u_cordic/mycordic/present_Q_table[5][0] ,
         \u_cordic/mycordic/present_Q_table[5][1] ,
         \u_cordic/mycordic/present_Q_table[5][2] ,
         \u_cordic/mycordic/present_Q_table[5][3] ,
         \u_cordic/mycordic/present_Q_table[5][4] ,
         \u_cordic/mycordic/present_Q_table[5][5] ,
         \u_cordic/mycordic/present_Q_table[5][6] ,
         \u_cordic/mycordic/present_Q_table[5][7] ,
         \u_cordic/mycordic/present_Q_table[6][7] ,
         \u_cordic/mycordic/present_I_table[0][3] ,
         \u_cordic/mycordic/present_I_table[0][4] ,
         \u_cordic/mycordic/present_I_table[0][5] ,
         \u_cordic/mycordic/present_I_table[0][6] ,
         \u_cordic/mycordic/present_I_table[0][7] ,
         \u_cordic/mycordic/present_I_table[1][3] ,
         \u_cordic/mycordic/present_I_table[1][4] ,
         \u_cordic/mycordic/present_I_table[1][5] ,
         \u_cordic/mycordic/present_I_table[1][6] ,
         \u_cordic/mycordic/present_I_table[1][7] ,
         \u_cordic/mycordic/present_I_table[2][0] ,
         \u_cordic/mycordic/present_I_table[2][1] ,
         \u_cordic/mycordic/present_I_table[2][2] ,
         \u_cordic/mycordic/present_I_table[2][3] ,
         \u_cordic/mycordic/present_I_table[2][4] ,
         \u_cordic/mycordic/present_I_table[2][5] ,
         \u_cordic/mycordic/present_I_table[2][6] ,
         \u_cordic/mycordic/present_I_table[2][7] ,
         \u_cordic/mycordic/present_I_table[3][0] ,
         \u_cordic/mycordic/present_I_table[3][1] ,
         \u_cordic/mycordic/present_I_table[3][2] ,
         \u_cordic/mycordic/present_I_table[3][3] ,
         \u_cordic/mycordic/present_I_table[3][4] ,
         \u_cordic/mycordic/present_I_table[3][5] ,
         \u_cordic/mycordic/present_I_table[3][6] ,
         \u_cordic/mycordic/present_I_table[3][7] ,
         \u_cordic/mycordic/present_I_table[4][0] ,
         \u_cordic/mycordic/present_I_table[4][1] ,
         \u_cordic/mycordic/present_I_table[4][2] ,
         \u_cordic/mycordic/present_I_table[4][3] ,
         \u_cordic/mycordic/present_I_table[4][4] ,
         \u_cordic/mycordic/present_I_table[4][5] ,
         \u_cordic/mycordic/present_I_table[4][6] ,
         \u_cordic/mycordic/present_I_table[4][7] ,
         \u_cordic/mycordic/present_I_table[5][4] ,
         \u_cordic/mycordic/present_I_table[5][5] ,
         \u_cordic/mycordic/present_I_table[5][6] ,
         \u_cordic/mycordic/present_I_table[5][7] ,
         \u_cordic/my_rotation/n117 , \u_cordic/my_rotation/n116 ,
         \u_cordic/my_rotation/n115 , \u_cordic/my_rotation/n114 ,
         \u_cordic/my_rotation/n113 , \u_cordic/my_rotation/n112 ,
         \u_cordic/my_rotation/n111 , \u_cordic/my_rotation/n110 ,
         \u_cordic/my_rotation/n109 , \u_cordic/my_rotation/n108 ,
         \u_cordic/my_rotation/n107 , \u_cordic/my_rotation/n106 ,
         \u_cordic/my_rotation/n105 , \u_cordic/my_rotation/n104 ,
         \u_cordic/my_rotation/n103 , \u_cordic/my_rotation/n102 ,
         \u_cordic/my_rotation/n101 , \u_cordic/my_rotation/n100 ,
         \u_cordic/my_rotation/n99 , \u_cordic/my_rotation/n98 ,
         \u_cordic/my_rotation/n97 , \u_cordic/my_rotation/n96 ,
         \u_cordic/my_rotation/n95 , \u_cordic/my_rotation/n94 ,
         \u_cordic/my_rotation/n93 , \u_cordic/my_rotation/n92 ,
         \u_cordic/my_rotation/n91 , \u_cordic/my_rotation/n90 ,
         \u_cordic/my_rotation/n89 , \u_cordic/my_rotation/n88 ,
         \u_cordic/my_rotation/n87 , \u_cordic/my_rotation/n86 ,
         \u_cordic/my_rotation/n85 , \u_cordic/my_rotation/n84 ,
         \u_cordic/my_rotation/n83 , \u_cordic/my_rotation/n82 ,
         \u_cordic/my_rotation/n81 , \u_cordic/my_rotation/n80 ,
         \u_cordic/my_rotation/n79 , \u_cordic/my_rotation/n78 ,
         \u_cordic/my_rotation/n77 , \u_cordic/my_rotation/n76 ,
         \u_cordic/my_rotation/n75 , \u_cordic/my_rotation/n74 ,
         \u_cordic/my_rotation/n73 , \u_cordic/my_rotation/n72 ,
         \u_cordic/my_rotation/n71 , \u_cordic/my_rotation/n70 ,
         \u_cordic/my_rotation/n69 , \u_cordic/my_rotation/n68 ,
         \u_cordic/my_rotation/n67 , \u_cordic/my_rotation/n66 ,
         \u_cordic/my_rotation/n65 , \u_cordic/my_rotation/n64 ,
         \u_cordic/my_rotation/n63 , \u_cordic/my_rotation/N56 ,
         \u_cordic/my_rotation/N55 , \u_cordic/my_rotation/N54 ,
         \u_cordic/my_rotation/N53 , \u_cordic/my_rotation/N52 ,
         \u_cordic/my_rotation/N51 , \u_cordic/my_rotation/N50 ,
         \u_cordic/my_rotation/N49 , \u_cordic/my_rotation/N48 ,
         \u_cordic/my_rotation/N47 , \u_cordic/my_rotation/N46 ,
         \u_cordic/my_rotation/N45 , \u_cordic/my_rotation/N41 ,
         \u_cordic/my_rotation/N39 ,
         \u_cordic/my_rotation/present_angle[0][15] ,
         \u_cordic/my_rotation/present_angle[0][14] ,
         \u_cordic/my_rotation/present_angle[0][13] ,
         \u_cordic/my_rotation/present_angle[0][12] ,
         \u_cordic/my_rotation/present_angle[0][11] ,
         \u_cordic/my_rotation/present_angle[0][10] ,
         \u_cordic/my_rotation/present_angle[0][9] ,
         \u_cordic/my_rotation/present_angle[0][8] ,
         \u_cordic/my_rotation/present_angle[0][7] ,
         \u_cordic/my_rotation/present_angle[0][6] ,
         \u_cordic/my_rotation/present_angle[0][5] ,
         \u_cordic/my_rotation/present_angle[0][4] ,
         \u_cordic/my_rotation/present_angle[0][3] ,
         \u_cordic/my_rotation/present_angle[0][2] ,
         \u_cordic/my_rotation/present_angle[0][1] ,
         \u_cordic/my_rotation/present_angle[0][0] , \u_cdr/div1/n39 ,
         \u_cdr/div1/n38 , \u_cdr/div1/n37 , \u_cdr/div1/n36 ,
         \u_cdr/div1/n35 , \u_cdr/div1/n34 , \u_cdr/div1/n31 ,
         \u_cdr/div1/n30 , \u_cdr/div1/n26 , \u_cdr/div1/n10 , \u_cdr/div1/n9 ,
         \u_cdr/div1/n8 , \u_cdr/div1/n7 , \u_cdr/div1/N34 ,
         \u_cdr/div1/w_en_freq_synch , \u_cdr/phd1/n21 , \u_cdr/phd1/n20 ,
         \u_cdr/phd1/n19 , \u_cdr/phd1/n18 , \u_cdr/phd1/n17 ,
         \u_cdr/phd1/n16 , \u_cdr/phd1/n15 , \u_cdr/phd1/n14 ,
         \u_cdr/phd1/n13 , \u_cdr/phd1/n12 , \u_cdr/phd1/n11 ,
         \u_cdr/phd1/n10 , \u_cdr/phd1/n9 , \u_cdr/phd1/w_s4 ,
         \u_cdr/phd1/w_s3 , \u_cdr/phd1/w_s2 , \u_cdr/phd1/w_s1 ,
         \u_cdr/phd1/w_en_f , \u_cdr/phd1/w_en_m , \u_cdr/phd1/w_en_d ,
         \u_cdr/dec1/n33 , \u_cdr/dec1/n32 , \u_cdr/dec1/n31 ,
         \u_cdr/dec1/n30 , \u_cdr/dec1/n29 , \u_cdr/dec1/n26 ,
         \u_cdr/dec1/n25 , \u_cdr/dec1/n24 , \u_cdr/dec1/n20 ,
         \u_cdr/dec1/w_en_dec , \u_cdr/dec1/N73 , \u_cdr/dec1/N65 ,
         \u_cdr/dec1/N64 , \u_cdr/dec1/N63 , \u_cdr/dec1/N62 ,
         \u_cdr/dec1/N61 , \u_cdr/dec1/w_s_r , \u_inFIFO/os1/dff1/n2 ,
         \u_decoder/iq_demod/cossin_dig/n56 ,
         \u_decoder/iq_demod/cossin_dig/n55 ,
         \u_decoder/iq_demod/cossin_dig/n54 ,
         \u_decoder/iq_demod/cossin_dig/n53 ,
         \u_decoder/iq_demod/cossin_dig/n52 ,
         \u_decoder/iq_demod/cossin_dig/n51 ,
         \u_decoder/iq_demod/cossin_dig/n50 ,
         \u_decoder/iq_demod/cossin_dig/n49 ,
         \u_decoder/iq_demod/cossin_dig/n48 ,
         \u_decoder/iq_demod/cossin_dig/n47 ,
         \u_decoder/iq_demod/cossin_dig/n46 ,
         \u_decoder/iq_demod/cossin_dig/n45 ,
         \u_decoder/iq_demod/cossin_dig/n44 ,
         \u_decoder/iq_demod/cossin_dig/n43 ,
         \u_decoder/iq_demod/cossin_dig/n42 ,
         \u_decoder/iq_demod/cossin_dig/n41 ,
         \u_decoder/iq_demod/cossin_dig/n40 ,
         \u_decoder/iq_demod/cossin_dig/n39 ,
         \u_decoder/iq_demod/cossin_dig/n38 ,
         \u_decoder/iq_demod/cossin_dig/n37 ,
         \u_decoder/iq_demod/cossin_dig/n36 ,
         \u_decoder/iq_demod/cossin_dig/n35 ,
         \u_decoder/iq_demod/cossin_dig/n34 ,
         \u_decoder/iq_demod/cossin_dig/n33 ,
         \u_decoder/iq_demod/cossin_dig/n32 ,
         \u_decoder/iq_demod/cossin_dig/n31 ,
         \u_decoder/iq_demod/cossin_dig/n30 ,
         \u_decoder/iq_demod/cossin_dig/n29 ,
         \u_decoder/iq_demod/cossin_dig/n28 ,
         \u_decoder/iq_demod/cossin_dig/n27 ,
         \u_decoder/iq_demod/cossin_dig/n26 ,
         \u_decoder/iq_demod/cossin_dig/n25 ,
         \u_decoder/iq_demod/cossin_dig/n23 ,
         \u_decoder/iq_demod/cossin_dig/n21 ,
         \u_decoder/iq_demod/cossin_dig/n19 ,
         \u_decoder/iq_demod/cossin_dig/n10 ,
         \u_decoder/iq_demod/cossin_dig/N60 ,
         \u_decoder/iq_demod/cossin_dig/N55 ,
         \u_decoder/iq_demod/cossin_dig/N52 ,
         \u_decoder/iq_demod/cossin_dig/N42 ,
         \u_decoder/iq_demod/cossin_dig/N41 ,
         \u_decoder/iq_demod/cossin_dig/N22 ,
         \u_decoder/iq_demod/cossin_dig/N21 ,
         \u_decoder/iq_demod/cossin_dig/N20 ,
         \u_decoder/iq_demod/cossin_dig/state[0] , \u_cdr/div1/cnt_div/n50 ,
         \u_cdr/div1/cnt_div/n48 , \u_cdr/div1/cnt_div/n47 ,
         \u_cdr/div1/cnt_div/n46 , \u_cdr/div1/cnt_div/n45 ,
         \u_cdr/div1/cnt_div/n44 , \u_cdr/div1/cnt_div/n43 ,
         \u_cdr/div1/cnt_div/n42 , \u_cdr/div1/cnt_div/n41 ,
         \u_cdr/div1/cnt_div/n40 , \u_cdr/div1/cnt_div/N84 ,
         \u_cdr/div1/cnt_div/N83 , \u_cdr/div1/cnt_div/N82 ,
         \u_cdr/div1/cnt_div/N81 , \u_cdr/div1/cnt_div/N80 ,
         \u_cdr/div1/cnt_div/N76 , \u_cdr/div1/cnt_div/N67 ,
         \u_cdr/phd1/f1/n2 , \u_outFIFO/os2/sigQout2 ,
         \u_outFIFO/os2/sigQout1 , \u_outFIFO/os1/sigQout2 ,
         \u_outFIFO/os1/sigQout1 , \u_inFIFO/os2/sigQout2 ,
         \u_inFIFO/os2/sigQout1 , \u_cdr/dec1/cnt_dec/N84 ,
         \u_cdr/dec1/cnt_dec/N83 , \u_cdr/dec1/cnt_dec/N82 ,
         \u_cdr/dec1/cnt_dec/N81 , \u_cdr/dec1/cnt_dec/N80 ,
         \u_cdr/dec1/cnt_dec/N76 , \u_cdr/dec1/cnt_dec/N43 ,
         \u_cdr/phd1/cnt_phd/N92 , \u_cdr/phd1/cnt_phd/N84 ,
         \u_cdr/phd1/cnt_phd/N83 , \u_cdr/phd1/cnt_phd/N82 ,
         \u_cdr/phd1/cnt_phd/N81 , \u_cdr/phd1/cnt_phd/N80 ,
         \u_cdr/phd1/cnt_phd/N76 , \u_cdr/phd1/cnt_phd/N59 ,
         \u_cdr/phd1/cnt_phd/N51 , \u_cdr/phd1/cnt_phd/N42 ,
         \u_cdr/phd1/cnt_phd/N41 , \u_cdr/phd1/cnt_phd/N14 ,
         \u_cdr/phd1/cnt_phd/N13 , \u_cdr/phd1/cnt_phd/N12 ,
         \u_cordic/mycordic/add_191/carry[2] ,
         \u_cordic/mycordic/add_191/carry[3] ,
         \u_cordic/mycordic/add_191/carry[4] ,
         \u_cordic/mycordic/add_191/carry[5] ,
         \u_cordic/mycordic/add_191/carry[6] ,
         \u_cordic/mycordic/add_191/carry[7] ,
         \u_cordic/mycordic/add_191/carry[8] ,
         \u_cordic/mycordic/add_191/carry[9] ,
         \u_cordic/mycordic/add_191/carry[10] ,
         \u_cordic/mycordic/add_191/carry[11] ,
         \u_cordic/mycordic/add_191/carry[12] ,
         \u_cordic/mycordic/add_191/carry[13] ,
         \u_cordic/mycordic/add_191/carry[14] ,
         \u_cordic/mycordic/add_191/carry[15] ,
         \u_cordic/mycordic/sub_196/carry[2] ,
         \u_cordic/mycordic/sub_196/carry[3] ,
         \u_cordic/mycordic/sub_196/carry[4] ,
         \u_cordic/mycordic/sub_196/carry[5] ,
         \u_cordic/mycordic/sub_196/carry[6] ,
         \u_cordic/mycordic/sub_196/carry[7] ,
         \u_cordic/mycordic/sub_196/carry[8] ,
         \u_cordic/mycordic/sub_196/carry[9] ,
         \u_cordic/mycordic/sub_196/carry[10] ,
         \u_cordic/mycordic/sub_196/carry[11] ,
         \u_cordic/mycordic/sub_196/carry[12] ,
         \u_cordic/mycordic/sub_196/carry[13] ,
         \u_cordic/mycordic/sub_196/carry[14] ,
         \u_cordic/mycordic/sub_196/carry[15] ,
         \u_cordic/mycordic/add_213/carry[2] ,
         \u_cordic/mycordic/add_213/carry[3] ,
         \u_cordic/mycordic/add_213/carry[4] ,
         \u_cordic/mycordic/add_213/carry[5] ,
         \u_cordic/mycordic/add_213/carry[6] ,
         \u_cordic/mycordic/add_213/carry[7] ,
         \u_cordic/mycordic/add_213/carry[8] ,
         \u_cordic/mycordic/add_213/carry[9] ,
         \u_cordic/mycordic/add_213/carry[10] ,
         \u_cordic/mycordic/add_213/carry[11] ,
         \u_cordic/mycordic/add_213/carry[12] ,
         \u_cordic/mycordic/add_213/carry[13] ,
         \u_cordic/mycordic/add_213/carry[14] ,
         \u_cordic/mycordic/add_213/carry[15] ,
         \u_cordic/mycordic/sub_218/carry[2] ,
         \u_cordic/mycordic/sub_218/carry[3] ,
         \u_cordic/mycordic/sub_218/carry[4] ,
         \u_cordic/mycordic/sub_218/carry[5] ,
         \u_cordic/mycordic/sub_218/carry[6] ,
         \u_cordic/mycordic/sub_218/carry[7] ,
         \u_cordic/mycordic/sub_218/carry[8] ,
         \u_cordic/mycordic/sub_218/carry[9] ,
         \u_cordic/mycordic/sub_218/carry[10] ,
         \u_cordic/mycordic/sub_218/carry[11] ,
         \u_cordic/mycordic/sub_218/carry[12] ,
         \u_cordic/mycordic/sub_218/carry[13] ,
         \u_cordic/mycordic/sub_218/carry[14] ,
         \u_cordic/mycordic/sub_218/carry[15] ,
         \u_cordic/mycordic/sub_223/carry[7] ,
         \u_cordic/mycordic/add_224/carry[2] ,
         \u_cordic/mycordic/add_224/carry[3] ,
         \u_cordic/mycordic/add_224/carry[4] ,
         \u_cordic/mycordic/add_224/carry[5] ,
         \u_cordic/mycordic/add_224/carry[6] ,
         \u_cordic/mycordic/add_224/carry[7] ,
         \u_cordic/mycordic/add_224/carry[8] ,
         \u_cordic/mycordic/add_224/carry[9] ,
         \u_cordic/mycordic/add_224/carry[10] ,
         \u_cordic/mycordic/add_224/carry[11] ,
         \u_cordic/mycordic/add_224/carry[12] ,
         \u_cordic/mycordic/add_224/carry[13] ,
         \u_cordic/mycordic/add_224/carry[14] ,
         \u_cordic/mycordic/add_224/carry[15] ,
         \u_cordic/mycordic/add_228/carry[7] ,
         \u_cordic/mycordic/sub_229/carry[2] ,
         \u_cordic/mycordic/sub_229/carry[3] ,
         \u_cordic/mycordic/sub_229/carry[4] ,
         \u_cordic/mycordic/sub_229/carry[5] ,
         \u_cordic/mycordic/sub_229/carry[6] ,
         \u_cordic/mycordic/sub_229/carry[7] ,
         \u_cordic/mycordic/sub_229/carry[8] ,
         \u_cordic/mycordic/sub_229/carry[9] ,
         \u_cordic/mycordic/sub_229/carry[10] ,
         \u_cordic/mycordic/sub_229/carry[11] ,
         \u_cordic/mycordic/sub_229/carry[12] ,
         \u_cordic/mycordic/sub_229/carry[13] ,
         \u_cordic/mycordic/sub_229/carry[14] ,
         \u_cordic/mycordic/sub_229/carry[15] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_276/A2[7] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_276/A2[8] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_276/A2[9] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_276/A2[10] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_276/A2[11] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_276/A1[7] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_276/A1[8] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_276/A1[9] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_276/A1[10] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_276/SUMB[1][5] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_276/SUMB[2][3] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_276/SUMB[2][5] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_276/SUMB[3][3] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_276/SUMB[3][5] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_276/SUMB[4][3] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_276/SUMB[4][5] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_276/SUMB[5][3] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_276/SUMB[5][5] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_276/SUMB[6][3] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_276/SUMB[6][5] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_276/SUMB[7][0] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_276/SUMB[7][1] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_276/SUMB[7][2] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_276/SUMB[7][3] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_276/SUMB[7][4] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_276/SUMB[7][5] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[1][5] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[2][3] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[2][5] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[3][0] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[3][3] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[3][5] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[4][0] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[4][3] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[4][5] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[5][0] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[5][3] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[5][5] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[6][0] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[6][3] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[6][5] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[7][0] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[7][1] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[7][2] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[7][3] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[7][4] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[7][5] ,
         \u_decoder/fir_filter/dp_cluster_0/r167/A2[7] ,
         \u_decoder/fir_filter/dp_cluster_0/r167/A2[8] ,
         \u_decoder/fir_filter/dp_cluster_0/r167/A2[9] ,
         \u_decoder/fir_filter/dp_cluster_0/r167/A2[10] ,
         \u_decoder/fir_filter/dp_cluster_0/r167/A2[11] ,
         \u_decoder/fir_filter/dp_cluster_0/r167/A1[7] ,
         \u_decoder/fir_filter/dp_cluster_0/r167/A1[8] ,
         \u_decoder/fir_filter/dp_cluster_0/r167/A1[9] ,
         \u_decoder/fir_filter/dp_cluster_0/r167/A1[10] ,
         \u_decoder/fir_filter/dp_cluster_0/r167/SUMB[2][1] ,
         \u_decoder/fir_filter/dp_cluster_0/r167/SUMB[3][1] ,
         \u_decoder/fir_filter/dp_cluster_0/r167/SUMB[3][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r167/SUMB[4][1] ,
         \u_decoder/fir_filter/dp_cluster_0/r167/SUMB[4][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r167/SUMB[5][1] ,
         \u_decoder/fir_filter/dp_cluster_0/r167/SUMB[5][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r167/SUMB[6][1] ,
         \u_decoder/fir_filter/dp_cluster_0/r167/SUMB[6][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r167/SUMB[7][0] ,
         \u_decoder/fir_filter/dp_cluster_0/r167/SUMB[7][1] ,
         \u_decoder/fir_filter/dp_cluster_0/r167/SUMB[7][2] ,
         \u_decoder/fir_filter/dp_cluster_0/r167/SUMB[7][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r167/SUMB[7][4] ,
         \u_decoder/fir_filter/dp_cluster_0/r167/SUMB[7][5] ,
         \u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[1][0] ,
         \u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[2][0] ,
         \u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[2][1] ,
         \u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[3][0] ,
         \u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[3][1] ,
         \u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[3][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[4][0] ,
         \u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[4][1] ,
         \u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[4][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[5][0] ,
         \u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[5][1] ,
         \u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[5][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[6][0] ,
         \u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[6][1] ,
         \u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[6][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[7][0] ,
         \u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[7][1] ,
         \u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[7][2] ,
         \u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[7][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[7][4] ,
         \u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[7][5] ,
         \u_decoder/fir_filter/dp_cluster_0/r166/A2[6] ,
         \u_decoder/fir_filter/dp_cluster_0/r166/A2[7] ,
         \u_decoder/fir_filter/dp_cluster_0/r166/A2[8] ,
         \u_decoder/fir_filter/dp_cluster_0/r166/A2[9] ,
         \u_decoder/fir_filter/dp_cluster_0/r166/A1[6] ,
         \u_decoder/fir_filter/dp_cluster_0/r166/A1[7] ,
         \u_decoder/fir_filter/dp_cluster_0/r166/A1[8] ,
         \u_decoder/fir_filter/dp_cluster_0/r166/SUMB[1][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r166/SUMB[2][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r166/SUMB[3][1] ,
         \u_decoder/fir_filter/dp_cluster_0/r166/SUMB[3][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r166/SUMB[4][1] ,
         \u_decoder/fir_filter/dp_cluster_0/r166/SUMB[4][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r166/SUMB[5][1] ,
         \u_decoder/fir_filter/dp_cluster_0/r166/SUMB[5][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r166/SUMB[6][1] ,
         \u_decoder/fir_filter/dp_cluster_0/r166/SUMB[6][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r166/SUMB[7][0] ,
         \u_decoder/fir_filter/dp_cluster_0/r166/SUMB[7][1] ,
         \u_decoder/fir_filter/dp_cluster_0/r166/SUMB[7][2] ,
         \u_decoder/fir_filter/dp_cluster_0/r166/SUMB[7][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r166/CARRYB[1][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r166/CARRYB[2][1] ,
         \u_decoder/fir_filter/dp_cluster_0/r166/CARRYB[2][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r166/CARRYB[3][1] ,
         \u_decoder/fir_filter/dp_cluster_0/r166/CARRYB[3][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r166/CARRYB[4][1] ,
         \u_decoder/fir_filter/dp_cluster_0/r166/CARRYB[4][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r166/CARRYB[5][1] ,
         \u_decoder/fir_filter/dp_cluster_0/r166/CARRYB[5][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r166/CARRYB[6][1] ,
         \u_decoder/fir_filter/dp_cluster_0/r166/CARRYB[6][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r166/CARRYB[7][0] ,
         \u_decoder/fir_filter/dp_cluster_0/r166/CARRYB[7][1] ,
         \u_decoder/fir_filter/dp_cluster_0/r166/CARRYB[7][2] ,
         \u_decoder/fir_filter/dp_cluster_0/r166/CARRYB[7][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r165/A2[6] ,
         \u_decoder/fir_filter/dp_cluster_0/r165/A2[7] ,
         \u_decoder/fir_filter/dp_cluster_0/r165/A2[8] ,
         \u_decoder/fir_filter/dp_cluster_0/r165/A2[9] ,
         \u_decoder/fir_filter/dp_cluster_0/r165/A2[10] ,
         \u_decoder/fir_filter/dp_cluster_0/r165/A1[4] ,
         \u_decoder/fir_filter/dp_cluster_0/r165/A1[5] ,
         \u_decoder/fir_filter/dp_cluster_0/r165/A1[6] ,
         \u_decoder/fir_filter/dp_cluster_0/r165/A1[7] ,
         \u_decoder/fir_filter/dp_cluster_0/r165/A1[8] ,
         \u_decoder/fir_filter/dp_cluster_0/r165/A1[9] ,
         \u_decoder/fir_filter/dp_cluster_0/r165/PROD1[5] ,
         \u_decoder/fir_filter/dp_cluster_0/r165/SUMB[2][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r165/SUMB[3][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r165/SUMB[4][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r165/SUMB[5][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r165/SUMB[6][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r165/SUMB[7][0] ,
         \u_decoder/fir_filter/dp_cluster_0/r165/SUMB[7][1] ,
         \u_decoder/fir_filter/dp_cluster_0/r165/SUMB[7][2] ,
         \u_decoder/fir_filter/dp_cluster_0/r165/SUMB[7][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r165/SUMB[7][4] ,
         \u_decoder/fir_filter/dp_cluster_0/r165/CARRYB[2][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r165/CARRYB[3][0] ,
         \u_decoder/fir_filter/dp_cluster_0/r165/CARRYB[3][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r165/CARRYB[4][0] ,
         \u_decoder/fir_filter/dp_cluster_0/r165/CARRYB[4][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r165/CARRYB[5][0] ,
         \u_decoder/fir_filter/dp_cluster_0/r165/CARRYB[5][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r165/CARRYB[6][0] ,
         \u_decoder/fir_filter/dp_cluster_0/r165/CARRYB[6][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r165/CARRYB[7][0] ,
         \u_decoder/fir_filter/dp_cluster_0/r165/CARRYB[7][1] ,
         \u_decoder/fir_filter/dp_cluster_0/r165/CARRYB[7][2] ,
         \u_decoder/fir_filter/dp_cluster_0/r165/CARRYB[7][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r165/CARRYB[7][4] ,
         \u_decoder/fir_filter/dp_cluster_0/r164/A2[6] ,
         \u_decoder/fir_filter/dp_cluster_0/r164/A2[7] ,
         \u_decoder/fir_filter/dp_cluster_0/r164/A2[8] ,
         \u_decoder/fir_filter/dp_cluster_0/r164/A2[9] ,
         \u_decoder/fir_filter/dp_cluster_0/r164/A1[3] ,
         \u_decoder/fir_filter/dp_cluster_0/r164/A1[4] ,
         \u_decoder/fir_filter/dp_cluster_0/r164/A1[5] ,
         \u_decoder/fir_filter/dp_cluster_0/r164/A1[6] ,
         \u_decoder/fir_filter/dp_cluster_0/r164/A1[7] ,
         \u_decoder/fir_filter/dp_cluster_0/r164/A1[8] ,
         \u_decoder/fir_filter/dp_cluster_0/r164/PROD1[4] ,
         \u_decoder/fir_filter/dp_cluster_0/r164/SUMB[2][2] ,
         \u_decoder/fir_filter/dp_cluster_0/r164/SUMB[3][2] ,
         \u_decoder/fir_filter/dp_cluster_0/r164/SUMB[4][2] ,
         \u_decoder/fir_filter/dp_cluster_0/r164/SUMB[5][2] ,
         \u_decoder/fir_filter/dp_cluster_0/r164/SUMB[6][2] ,
         \u_decoder/fir_filter/dp_cluster_0/r164/SUMB[7][0] ,
         \u_decoder/fir_filter/dp_cluster_0/r164/SUMB[7][1] ,
         \u_decoder/fir_filter/dp_cluster_0/r164/SUMB[7][2] ,
         \u_decoder/fir_filter/dp_cluster_0/r164/SUMB[7][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r164/CARRYB[2][0] ,
         \u_decoder/fir_filter/dp_cluster_0/r164/CARRYB[2][2] ,
         \u_decoder/fir_filter/dp_cluster_0/r164/CARRYB[3][0] ,
         \u_decoder/fir_filter/dp_cluster_0/r164/CARRYB[3][2] ,
         \u_decoder/fir_filter/dp_cluster_0/r164/CARRYB[4][0] ,
         \u_decoder/fir_filter/dp_cluster_0/r164/CARRYB[4][2] ,
         \u_decoder/fir_filter/dp_cluster_0/r164/CARRYB[5][0] ,
         \u_decoder/fir_filter/dp_cluster_0/r164/CARRYB[5][2] ,
         \u_decoder/fir_filter/dp_cluster_0/r164/CARRYB[6][0] ,
         \u_decoder/fir_filter/dp_cluster_0/r164/CARRYB[6][2] ,
         \u_decoder/fir_filter/dp_cluster_0/r164/CARRYB[7][0] ,
         \u_decoder/fir_filter/dp_cluster_0/r164/CARRYB[7][1] ,
         \u_decoder/fir_filter/dp_cluster_0/r164/CARRYB[7][2] ,
         \u_decoder/fir_filter/dp_cluster_0/r164/CARRYB[7][3] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_308/A2[7] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_308/A2[8] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_308/A2[9] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_308/A2[10] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_308/A2[11] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_308/A1[7] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_308/A1[8] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_308/A1[9] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_308/A1[10] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_308/SUMB[1][5] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_308/SUMB[2][3] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_308/SUMB[2][5] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_308/SUMB[3][3] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_308/SUMB[3][5] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_308/SUMB[4][3] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_308/SUMB[4][5] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_308/SUMB[5][3] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_308/SUMB[5][5] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_308/SUMB[6][3] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_308/SUMB[6][5] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_308/SUMB[7][0] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_308/SUMB[7][1] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_308/SUMB[7][2] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_308/SUMB[7][3] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_308/SUMB[7][4] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_308/SUMB[7][5] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[1][5] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[2][3] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[2][5] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[3][0] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[3][3] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[3][5] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[4][0] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[4][3] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[4][5] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[5][0] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[5][3] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[5][5] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[6][0] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[6][3] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[6][5] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[7][0] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[7][1] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[7][2] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[7][3] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[7][4] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[7][5] ,
         \u_decoder/fir_filter/dp_cluster_0/r180/A2[7] ,
         \u_decoder/fir_filter/dp_cluster_0/r180/A2[8] ,
         \u_decoder/fir_filter/dp_cluster_0/r180/A2[9] ,
         \u_decoder/fir_filter/dp_cluster_0/r180/A2[10] ,
         \u_decoder/fir_filter/dp_cluster_0/r180/A2[11] ,
         \u_decoder/fir_filter/dp_cluster_0/r180/A1[7] ,
         \u_decoder/fir_filter/dp_cluster_0/r180/A1[8] ,
         \u_decoder/fir_filter/dp_cluster_0/r180/A1[9] ,
         \u_decoder/fir_filter/dp_cluster_0/r180/A1[10] ,
         \u_decoder/fir_filter/dp_cluster_0/r180/SUMB[2][1] ,
         \u_decoder/fir_filter/dp_cluster_0/r180/SUMB[3][1] ,
         \u_decoder/fir_filter/dp_cluster_0/r180/SUMB[3][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r180/SUMB[4][1] ,
         \u_decoder/fir_filter/dp_cluster_0/r180/SUMB[4][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r180/SUMB[5][1] ,
         \u_decoder/fir_filter/dp_cluster_0/r180/SUMB[5][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r180/SUMB[6][1] ,
         \u_decoder/fir_filter/dp_cluster_0/r180/SUMB[6][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r180/SUMB[7][0] ,
         \u_decoder/fir_filter/dp_cluster_0/r180/SUMB[7][1] ,
         \u_decoder/fir_filter/dp_cluster_0/r180/SUMB[7][2] ,
         \u_decoder/fir_filter/dp_cluster_0/r180/SUMB[7][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r180/SUMB[7][4] ,
         \u_decoder/fir_filter/dp_cluster_0/r180/SUMB[7][5] ,
         \u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[1][0] ,
         \u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[2][0] ,
         \u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[2][1] ,
         \u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[3][0] ,
         \u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[3][1] ,
         \u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[3][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[4][0] ,
         \u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[4][1] ,
         \u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[4][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[5][0] ,
         \u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[5][1] ,
         \u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[5][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[6][0] ,
         \u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[6][1] ,
         \u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[6][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[7][0] ,
         \u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[7][1] ,
         \u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[7][2] ,
         \u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[7][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[7][4] ,
         \u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[7][5] ,
         \u_decoder/fir_filter/dp_cluster_0/r179/A2[6] ,
         \u_decoder/fir_filter/dp_cluster_0/r179/A2[7] ,
         \u_decoder/fir_filter/dp_cluster_0/r179/A2[8] ,
         \u_decoder/fir_filter/dp_cluster_0/r179/A2[9] ,
         \u_decoder/fir_filter/dp_cluster_0/r179/A1[6] ,
         \u_decoder/fir_filter/dp_cluster_0/r179/A1[7] ,
         \u_decoder/fir_filter/dp_cluster_0/r179/A1[8] ,
         \u_decoder/fir_filter/dp_cluster_0/r179/SUMB[1][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r179/SUMB[2][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r179/SUMB[3][1] ,
         \u_decoder/fir_filter/dp_cluster_0/r179/SUMB[3][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r179/SUMB[4][1] ,
         \u_decoder/fir_filter/dp_cluster_0/r179/SUMB[4][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r179/SUMB[5][1] ,
         \u_decoder/fir_filter/dp_cluster_0/r179/SUMB[5][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r179/SUMB[6][1] ,
         \u_decoder/fir_filter/dp_cluster_0/r179/SUMB[6][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r179/SUMB[7][0] ,
         \u_decoder/fir_filter/dp_cluster_0/r179/SUMB[7][1] ,
         \u_decoder/fir_filter/dp_cluster_0/r179/SUMB[7][2] ,
         \u_decoder/fir_filter/dp_cluster_0/r179/SUMB[7][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r179/CARRYB[1][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r179/CARRYB[2][1] ,
         \u_decoder/fir_filter/dp_cluster_0/r179/CARRYB[2][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r179/CARRYB[3][1] ,
         \u_decoder/fir_filter/dp_cluster_0/r179/CARRYB[3][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r179/CARRYB[4][1] ,
         \u_decoder/fir_filter/dp_cluster_0/r179/CARRYB[4][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r179/CARRYB[5][1] ,
         \u_decoder/fir_filter/dp_cluster_0/r179/CARRYB[5][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r179/CARRYB[6][1] ,
         \u_decoder/fir_filter/dp_cluster_0/r179/CARRYB[6][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r179/CARRYB[7][0] ,
         \u_decoder/fir_filter/dp_cluster_0/r179/CARRYB[7][1] ,
         \u_decoder/fir_filter/dp_cluster_0/r179/CARRYB[7][2] ,
         \u_decoder/fir_filter/dp_cluster_0/r179/CARRYB[7][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r178/A2[6] ,
         \u_decoder/fir_filter/dp_cluster_0/r178/A2[7] ,
         \u_decoder/fir_filter/dp_cluster_0/r178/A2[8] ,
         \u_decoder/fir_filter/dp_cluster_0/r178/A2[9] ,
         \u_decoder/fir_filter/dp_cluster_0/r178/A2[10] ,
         \u_decoder/fir_filter/dp_cluster_0/r178/A1[4] ,
         \u_decoder/fir_filter/dp_cluster_0/r178/A1[5] ,
         \u_decoder/fir_filter/dp_cluster_0/r178/A1[6] ,
         \u_decoder/fir_filter/dp_cluster_0/r178/A1[7] ,
         \u_decoder/fir_filter/dp_cluster_0/r178/A1[8] ,
         \u_decoder/fir_filter/dp_cluster_0/r178/A1[9] ,
         \u_decoder/fir_filter/dp_cluster_0/r178/PROD1[5] ,
         \u_decoder/fir_filter/dp_cluster_0/r178/SUMB[2][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r178/SUMB[3][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r178/SUMB[4][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r178/SUMB[5][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r178/SUMB[6][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r178/SUMB[7][0] ,
         \u_decoder/fir_filter/dp_cluster_0/r178/SUMB[7][1] ,
         \u_decoder/fir_filter/dp_cluster_0/r178/SUMB[7][2] ,
         \u_decoder/fir_filter/dp_cluster_0/r178/SUMB[7][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r178/SUMB[7][4] ,
         \u_decoder/fir_filter/dp_cluster_0/r178/CARRYB[2][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r178/CARRYB[3][0] ,
         \u_decoder/fir_filter/dp_cluster_0/r178/CARRYB[3][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r178/CARRYB[4][0] ,
         \u_decoder/fir_filter/dp_cluster_0/r178/CARRYB[4][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r178/CARRYB[5][0] ,
         \u_decoder/fir_filter/dp_cluster_0/r178/CARRYB[5][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r178/CARRYB[6][0] ,
         \u_decoder/fir_filter/dp_cluster_0/r178/CARRYB[6][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r178/CARRYB[7][0] ,
         \u_decoder/fir_filter/dp_cluster_0/r178/CARRYB[7][1] ,
         \u_decoder/fir_filter/dp_cluster_0/r178/CARRYB[7][2] ,
         \u_decoder/fir_filter/dp_cluster_0/r178/CARRYB[7][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r178/CARRYB[7][4] ,
         \u_decoder/fir_filter/dp_cluster_0/r177/A2[6] ,
         \u_decoder/fir_filter/dp_cluster_0/r177/A2[7] ,
         \u_decoder/fir_filter/dp_cluster_0/r177/A2[8] ,
         \u_decoder/fir_filter/dp_cluster_0/r177/A2[9] ,
         \u_decoder/fir_filter/dp_cluster_0/r177/A1[3] ,
         \u_decoder/fir_filter/dp_cluster_0/r177/A1[4] ,
         \u_decoder/fir_filter/dp_cluster_0/r177/A1[5] ,
         \u_decoder/fir_filter/dp_cluster_0/r177/A1[6] ,
         \u_decoder/fir_filter/dp_cluster_0/r177/A1[7] ,
         \u_decoder/fir_filter/dp_cluster_0/r177/A1[8] ,
         \u_decoder/fir_filter/dp_cluster_0/r177/PROD1[4] ,
         \u_decoder/fir_filter/dp_cluster_0/r177/SUMB[2][2] ,
         \u_decoder/fir_filter/dp_cluster_0/r177/SUMB[3][2] ,
         \u_decoder/fir_filter/dp_cluster_0/r177/SUMB[4][2] ,
         \u_decoder/fir_filter/dp_cluster_0/r177/SUMB[5][2] ,
         \u_decoder/fir_filter/dp_cluster_0/r177/SUMB[6][2] ,
         \u_decoder/fir_filter/dp_cluster_0/r177/SUMB[7][0] ,
         \u_decoder/fir_filter/dp_cluster_0/r177/SUMB[7][1] ,
         \u_decoder/fir_filter/dp_cluster_0/r177/SUMB[7][2] ,
         \u_decoder/fir_filter/dp_cluster_0/r177/SUMB[7][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r177/CARRYB[2][0] ,
         \u_decoder/fir_filter/dp_cluster_0/r177/CARRYB[2][2] ,
         \u_decoder/fir_filter/dp_cluster_0/r177/CARRYB[3][0] ,
         \u_decoder/fir_filter/dp_cluster_0/r177/CARRYB[3][2] ,
         \u_decoder/fir_filter/dp_cluster_0/r177/CARRYB[4][0] ,
         \u_decoder/fir_filter/dp_cluster_0/r177/CARRYB[4][2] ,
         \u_decoder/fir_filter/dp_cluster_0/r177/CARRYB[5][0] ,
         \u_decoder/fir_filter/dp_cluster_0/r177/CARRYB[5][2] ,
         \u_decoder/fir_filter/dp_cluster_0/r177/CARRYB[6][0] ,
         \u_decoder/fir_filter/dp_cluster_0/r177/CARRYB[6][2] ,
         \u_decoder/fir_filter/dp_cluster_0/r177/CARRYB[7][0] ,
         \u_decoder/fir_filter/dp_cluster_0/r177/CARRYB[7][1] ,
         \u_decoder/fir_filter/dp_cluster_0/r177/CARRYB[7][2] ,
         \u_decoder/fir_filter/dp_cluster_0/r177/CARRYB[7][3] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_151/A2[2] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_151/A2[3] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_151/A2[4] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_151/A2[5] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_151/A1[2] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_151/A1[3] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_151/A1[4] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_151/SUMB[1][1] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_151/SUMB[1][2] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_151/SUMB[2][1] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_151/SUMB[2][2] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_151/SUMB[3][0] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_151/SUMB[3][1] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_151/SUMB[3][2] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_151/SUMB[3][3] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_151/CARRYB[1][0] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_151/CARRYB[1][1] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_151/CARRYB[1][2] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_151/CARRYB[2][0] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_151/CARRYB[2][1] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_151/CARRYB[2][2] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_151/CARRYB[3][0] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_151/CARRYB[3][1] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_151/CARRYB[3][2] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_151/CARRYB[3][3] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_151/ab[0][1] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_151/ab[0][2] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_151/ab[0][3] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_151/ab[1][0] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_151/ab[1][1] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_151/ab[1][2] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_151/ab[1][3] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_151/ab[2][0] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_151/ab[2][1] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_151/ab[2][2] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_151/ab[2][3] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_151/ab[3][0] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_151/ab[3][1] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_151/ab[3][2] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_151/ab[3][3] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_148/A2[2] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_148/A2[3] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_148/A2[4] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_148/A2[5] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_148/A1[2] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_148/A1[3] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_148/A1[4] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_148/SUMB[1][1] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_148/SUMB[1][2] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_148/SUMB[2][1] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_148/SUMB[2][2] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_148/SUMB[3][0] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_148/SUMB[3][1] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_148/SUMB[3][2] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_148/SUMB[3][3] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_148/CARRYB[1][0] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_148/CARRYB[1][1] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_148/CARRYB[1][2] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_148/CARRYB[2][0] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_148/CARRYB[2][1] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_148/CARRYB[2][2] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_148/CARRYB[3][0] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_148/CARRYB[3][1] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_148/CARRYB[3][2] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_148/CARRYB[3][3] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_148/ab[0][1] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_148/ab[0][2] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_148/ab[0][3] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_148/ab[1][0] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_148/ab[1][1] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_148/ab[1][2] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_148/ab[1][3] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_148/ab[2][0] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_148/ab[2][1] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_148/ab[2][2] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_148/ab[2][3] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_148/ab[3][0] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_148/ab[3][1] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_148/ab[3][2] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_148/ab[3][3] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_150/A2[2] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_150/A2[3] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_150/A2[4] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_150/A2[5] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_150/A1[2] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_150/A1[3] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_150/A1[4] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_150/SUMB[1][1] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_150/SUMB[1][2] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_150/SUMB[2][1] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_150/SUMB[2][2] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_150/SUMB[3][0] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_150/SUMB[3][1] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_150/SUMB[3][2] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_150/SUMB[3][3] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_150/CARRYB[1][0] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_150/CARRYB[1][1] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_150/CARRYB[1][2] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_150/CARRYB[2][0] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_150/CARRYB[2][1] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_150/CARRYB[2][2] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_150/CARRYB[3][0] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_150/CARRYB[3][1] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_150/CARRYB[3][2] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_150/CARRYB[3][3] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_150/ab[0][1] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_150/ab[0][2] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_150/ab[0][3] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_150/ab[1][0] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_150/ab[1][1] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_150/ab[1][2] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_150/ab[1][3] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_150/ab[2][0] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_150/ab[2][1] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_150/ab[2][2] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_150/ab[2][3] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_150/ab[3][0] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_150/ab[3][1] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_150/ab[3][2] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_150/ab[3][3] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_149/A2[2] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_149/A2[3] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_149/A2[4] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_149/A2[5] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_149/A1[2] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_149/A1[3] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_149/A1[4] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_149/SUMB[1][1] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_149/SUMB[1][2] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_149/SUMB[2][1] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_149/SUMB[2][2] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_149/SUMB[3][0] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_149/SUMB[3][1] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_149/SUMB[3][2] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_149/SUMB[3][3] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_149/CARRYB[1][0] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_149/CARRYB[1][1] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_149/CARRYB[1][2] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_149/CARRYB[2][0] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_149/CARRYB[2][1] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_149/CARRYB[2][2] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_149/CARRYB[3][0] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_149/CARRYB[3][1] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_149/CARRYB[3][2] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_149/CARRYB[3][3] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_149/ab[0][1] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_149/ab[0][2] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_149/ab[0][3] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_149/ab[1][0] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_149/ab[1][1] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_149/ab[1][2] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_149/ab[1][3] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_149/ab[2][0] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_149/ab[2][1] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_149/ab[2][2] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_149/ab[2][3] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_149/ab[3][0] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_149/ab[3][1] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_149/ab[3][2] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_149/ab[3][3] ,
         \u_cdr/dp_cluster_0/mult_add_59_aco/PROD_not[0] ,
         \u_cdr/dp_cluster_0/mult_add_59_aco/PROD_not[1] ,
         \u_cdr/dp_cluster_0/mult_add_59_aco/PROD_not[2] ,
         \u_cdr/dp_cluster_0/mult_add_59_aco/PROD_not[3] , n1, n2, n3, n4, n5,
         n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
         n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
         n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
         n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
         n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
         n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
         n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
         n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
         n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
         n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
         n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
         n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
         n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
         n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
         n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
         n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
         n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
         n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
         n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
         n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
         n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
         n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
         n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
         n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
         n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
         n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404,
         n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414,
         n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424,
         n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434,
         n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444,
         n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454,
         n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464,
         n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474,
         n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484,
         n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494,
         n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504,
         n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514,
         n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524,
         n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534,
         n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544,
         n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554,
         n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564,
         n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574,
         n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584,
         n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594,
         n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604,
         n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614,
         n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624,
         n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634,
         n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644,
         n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654,
         n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664,
         n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674,
         n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684,
         n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694,
         n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704,
         n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714,
         n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724,
         n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734,
         n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744,
         n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754,
         n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764,
         n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774,
         n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784,
         n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794,
         n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804,
         n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814,
         n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824,
         n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834,
         n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844,
         n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854,
         n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864,
         n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874,
         n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884,
         n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894,
         n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904,
         n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914,
         n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924,
         n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934,
         n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944,
         n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954,
         n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964,
         n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974,
         n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984,
         n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994,
         n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004,
         n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014,
         n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024,
         n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034,
         n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044,
         n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054,
         n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064,
         n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074,
         n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084,
         n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094,
         n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104,
         n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114,
         n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124,
         n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134,
         n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144,
         n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154,
         n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164,
         n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174,
         n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184,
         n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194,
         n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204,
         n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214,
         n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224,
         n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234,
         n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244,
         n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254,
         n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264,
         n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274,
         n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284,
         n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294,
         n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304,
         n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314,
         n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324,
         n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334,
         n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344,
         n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354,
         n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364,
         n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374,
         n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384,
         n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394,
         n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404,
         n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414,
         n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424,
         n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434,
         n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444,
         n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454,
         n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464,
         n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474,
         n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484,
         n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494,
         n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504,
         n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514,
         n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524,
         n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534,
         n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544,
         n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554,
         n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564,
         n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574,
         n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584,
         n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594,
         n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604,
         n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614,
         n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624,
         n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634,
         n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644,
         n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654,
         n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664,
         n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674,
         n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684,
         n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693;
  wire   [3:0] sig_coder_outSinI;
  wire   [3:0] sig_coder_outSinQ;
  wire   [3:0] sig_coder_outSinIMasked;
  wire   [3:0] sig_coder_outSinQMasked;
  wire   [3:0] sig_decod_outI;
  wire   [3:0] sig_decod_outQ;
  wire   [3:0] sig_outFIFO_outData;
  wire   [7:0] sig_DEMUX_outDEMUX1;
  wire   [7:0] sig_DEMUX_outDEMUX2;
  wire   [7:0] sig_DEMUX_outDEMUX17;
  wire   [7:0] sig_DEMUX_outDEMUX18;
  wire   [3:0] sig_MUX_outMUX6;
  wire   [3:0] sig_MUX_outMUX7;
  wire   [4:0] \u_inFIFO/j_FIFO ;
  wire   [3:0] \u_inFIFO/currentState ;
  wire   [19:0] \u_coder/j ;
  wire   [19:0] \u_coder/i ;
  wire   [19:0] \u_coder/c ;
  wire   [7:0] \u_decoder/Q_prefilter ;
  wire   [7:0] \u_decoder/I_prefilter ;
  wire   [2:0] \u_cordic/present_state ;
  wire   [3:0] \u_cordic/Q ;
  wire   [3:0] \u_cordic/I ;
  wire   [15:0] \u_cordic/cordic_to_rotation ;
  wire   [5:0] \u_cdr/w_nb_P ;
  wire   [2:0] \u_cdr/cnt ;
  wire   [1:0] \u_cdr/cnt_d ;
  wire   [3:0] \u_cdr/cnt_in ;
  wire   [1:0] \u_outFIFO/k_FIFO ;
  wire   [4:0] \u_outFIFO/i_FIFO ;
  wire   [3:0] \u_outFIFO/currentState ;
  wire   [7:0] \u_decoder/iq_demod/dp_cluster_1/mult_I_sin_out ;
  wire   [7:0] \u_decoder/iq_demod/dp_cluster_1/mult_Q_cos_out ;
  wire   [7:0] \u_decoder/iq_demod/dp_cluster_0/mult_I_cos_out ;
  wire   [7:0] \u_decoder/iq_demod/dp_cluster_0/mult_Q_sin_out ;
  wire   [3:0] \u_decoder/iq_demod/Q_if_signed ;
  wire   [3:0] \u_decoder/iq_demod/I_if_signed ;
  wire   [7:0] \u_decoder/iq_demod/add_Q_out ;
  wire   [7:0] \u_decoder/iq_demod/add_I_out ;
  wire   [1:0] \u_decoder/iq_demod/state ;
  wire   [3:0] \u_decoder/iq_demod/sin_out ;
  wire   [3:0] \u_decoder/iq_demod/cos_out ;
  wire   [20:0] \u_decoder/fir_filter/Q_data_mult_8_buff ;
  wire   [15:0] \u_decoder/fir_filter/Q_data_mult_7_buff ;
  wire   [15:0] \u_decoder/fir_filter/Q_data_mult_6_buff ;
  wire   [15:0] \u_decoder/fir_filter/Q_data_mult_5_buff ;
  wire   [15:0] \u_decoder/fir_filter/Q_data_mult_4 ;
  wire   [15:0] \u_decoder/fir_filter/Q_data_mult_4_buff ;
  wire   [15:0] \u_decoder/fir_filter/Q_data_mult_3 ;
  wire   [15:0] \u_decoder/fir_filter/Q_data_mult_3_buff ;
  wire   [15:0] \u_decoder/fir_filter/Q_data_mult_2_buff ;
  wire   [15:0] \u_decoder/fir_filter/Q_data_mult_1_buff ;
  wire   [11:0] \u_decoder/fir_filter/Q_data_mult_0 ;
  wire   [14:0] \u_decoder/fir_filter/Q_data_mult_0_buff ;
  wire   [20:0] \u_decoder/fir_filter/Q_data_add_7 ;
  wire   [20:0] \u_decoder/fir_filter/Q_data_add_7_buff ;
  wire   [20:0] \u_decoder/fir_filter/Q_data_add_6 ;
  wire   [20:0] \u_decoder/fir_filter/Q_data_add_6_buff ;
  wire   [20:0] \u_decoder/fir_filter/Q_data_add_5 ;
  wire   [20:0] \u_decoder/fir_filter/Q_data_add_5_buff ;
  wire   [20:0] \u_decoder/fir_filter/Q_data_add_4 ;
  wire   [20:0] \u_decoder/fir_filter/Q_data_add_4_buff ;
  wire   [20:0] \u_decoder/fir_filter/Q_data_add_3 ;
  wire   [20:0] \u_decoder/fir_filter/Q_data_add_3_buff ;
  wire   [20:0] \u_decoder/fir_filter/Q_data_add_2 ;
  wire   [20:0] \u_decoder/fir_filter/Q_data_add_2_buff ;
  wire   [14:0] \u_decoder/fir_filter/Q_data_add_1 ;
  wire   [14:0] \u_decoder/fir_filter/Q_data_add_1_buff ;
  wire   [20:0] \u_decoder/fir_filter/I_data_mult_8_buff ;
  wire   [15:0] \u_decoder/fir_filter/I_data_mult_7_buff ;
  wire   [15:0] \u_decoder/fir_filter/I_data_mult_6_buff ;
  wire   [15:0] \u_decoder/fir_filter/I_data_mult_5_buff ;
  wire   [15:0] \u_decoder/fir_filter/I_data_mult_4 ;
  wire   [15:0] \u_decoder/fir_filter/I_data_mult_4_buff ;
  wire   [15:0] \u_decoder/fir_filter/I_data_mult_3 ;
  wire   [15:0] \u_decoder/fir_filter/I_data_mult_3_buff ;
  wire   [15:0] \u_decoder/fir_filter/I_data_mult_2_buff ;
  wire   [15:0] \u_decoder/fir_filter/I_data_mult_1_buff ;
  wire   [11:0] \u_decoder/fir_filter/I_data_mult_0 ;
  wire   [14:0] \u_decoder/fir_filter/I_data_mult_0_buff ;
  wire   [20:0] \u_decoder/fir_filter/I_data_add_7 ;
  wire   [20:0] \u_decoder/fir_filter/I_data_add_7_buff ;
  wire   [20:0] \u_decoder/fir_filter/I_data_add_6 ;
  wire   [20:0] \u_decoder/fir_filter/I_data_add_6_buff ;
  wire   [20:0] \u_decoder/fir_filter/I_data_add_5 ;
  wire   [20:0] \u_decoder/fir_filter/I_data_add_5_buff ;
  wire   [20:0] \u_decoder/fir_filter/I_data_add_4 ;
  wire   [20:0] \u_decoder/fir_filter/I_data_add_4_buff ;
  wire   [20:0] \u_decoder/fir_filter/I_data_add_3 ;
  wire   [20:0] \u_decoder/fir_filter/I_data_add_3_buff ;
  wire   [20:0] \u_decoder/fir_filter/I_data_add_2 ;
  wire   [20:0] \u_decoder/fir_filter/I_data_add_2_buff ;
  wire   [14:0] \u_decoder/fir_filter/I_data_add_1 ;
  wire   [14:0] \u_decoder/fir_filter/I_data_add_1_buff ;
  wire   [14:11] \u_decoder/fir_filter/Q_data_add_0 ;
  wire   [14:11] \u_decoder/fir_filter/I_data_add_0 ;
  wire   [1:0] \u_decoder/fir_filter/state ;
  wire   [15:0] \u_cordic/my_rotation/next_delta ;
  wire   [15:0] \u_cordic/my_rotation/present_delta ;
  wire   [5:0] \u_cdr/dec1/cnt_r ;
  wire   [2:0] \u_decoder/iq_demod/cossin_dig/val_counter ;
  wire   [2:0] \u_decoder/iq_demod/cossin_dig/counter ;
  wire   [5:0] \u_cdr/div1/cnt_div/cnt ;
  wire   [5:0] \u_cdr/dec1/cnt_dec/cnt ;
  wire   [5:0] \u_cdr/phd1/cnt_phd/cnt ;
  wire   [5:2] \u_cdr/phd1/cnt_phd/add_65/carry ;
  wire   [5:2] \u_cdr/dec1/cnt_dec/add_65/carry ;
  wire   [5:2] \u_cdr/div1/cnt_div/add_65/carry ;
  wire   [5:2] \u_cdr/dec1/add_41/carry ;
  wire   [16:0] \u_cordic/my_rotation/sub_40/carry ;
  wire   [15:1] \u_cordic/my_rotation/add_43/carry ;
  wire   [7:1] \u_cordic/mycordic/r144/carry ;
  wire   [15:1] \u_cordic/mycordic/r173/carry ;
  wire   [8:0] \u_cordic/mycordic/sub_178/carry ;
  wire   [8:0] \u_cordic/mycordic/sub_182/carry ;
  wire   [7:1] \u_cordic/mycordic/add_189/carry ;
  wire   [8:0] \u_cordic/mycordic/sub_190/carry ;
  wire   [8:0] \u_cordic/mycordic/sub_194/carry ;
  wire   [7:1] \u_cordic/mycordic/add_195/carry ;
  wire   [7:1] \u_cordic/mycordic/add_200/carry ;
  wire   [8:0] \u_cordic/mycordic/sub_201/carry ;
  wire   [15:1] \u_cordic/mycordic/add_202/carry ;
  wire   [8:0] \u_cordic/mycordic/sub_205/carry ;
  wire   [7:1] \u_cordic/mycordic/add_206/carry ;
  wire   [16:0] \u_cordic/mycordic/sub_207/carry ;
  wire   [7:1] \u_cordic/mycordic/add_211/carry ;
  wire   [8:0] \u_cordic/mycordic/sub_212/carry ;
  wire   [8:0] \u_cordic/mycordic/sub_216/carry ;
  wire   [7:1] \u_cordic/mycordic/add_217/carry ;
  wire   [15:1] \u_cordic/mycordic/add_233/carry ;
  wire   [16:0] \u_cordic/mycordic/sub_236/carry ;
  wire   [15:1] \u_cordic/mycordic/add_262/carry ;
  wire   [8:0] \u_cordic/mycordic/sub_add_150_b0/carry ;
  wire   [8:0] \u_cordic/mycordic/sub_add_151_b0/carry ;
  wire   [14:1] \u_decoder/fir_filter/add_294/carry ;
  wire   [20:1] \u_decoder/fir_filter/add_295/carry ;
  wire   [20:1] \u_decoder/fir_filter/add_296/carry ;
  wire   [20:1] \u_decoder/fir_filter/add_297/carry ;
  wire   [20:1] \u_decoder/fir_filter/add_298/carry ;
  wire   [20:1] \u_decoder/fir_filter/add_299/carry ;
  wire   [20:1] \u_decoder/fir_filter/add_300/carry ;
  wire   [20:1] \u_decoder/fir_filter/add_301/carry ;
  wire   [14:1] \u_decoder/fir_filter/add_326/carry ;
  wire   [20:1] \u_decoder/fir_filter/add_327/carry ;
  wire   [20:1] \u_decoder/fir_filter/add_328/carry ;
  wire   [20:1] \u_decoder/fir_filter/add_329/carry ;
  wire   [20:1] \u_decoder/fir_filter/add_330/carry ;
  wire   [20:1] \u_decoder/fir_filter/add_331/carry ;
  wire   [20:1] \u_decoder/fir_filter/add_332/carry ;
  wire   [20:1] \u_decoder/fir_filter/add_333/carry ;
  wire   [8:0] \u_decoder/iq_demod/dp_cluster_0/sub_153/carry ;
  wire   [7:1] \u_decoder/iq_demod/dp_cluster_1/add_154/carry ;
  wire   [6:0] \u_outFIFO/r98/carry ;
  wire   [5:2] \u_outFIFO/add_255/carry ;
  wire   [4:2] \u_outFIFO/add_256/carry ;
  wire   [4:2] \u_outFIFO/add_260/carry ;
  wire   [4:2] \u_outFIFO/add_360/carry ;
  wire   [19:2] \u_coder/add_93/carry ;
  wire   [19:2] \u_coder/add_206/carry ;
  wire   [19:2] \u_coder/add_282/carry ;
  wire   [6:0] \u_inFIFO/r96/carry ;
  wire   [4:2] \u_inFIFO/add_252/carry ;
  wire   [4:2] \u_inFIFO/add_253/carry ;
  wire   [5:2] \u_inFIFO/add_263/carry ;
  wire   [4:2] \u_inFIFO/add_357/carry ;

  OAI222 \u_inFIFO/U154  ( .A(n984), .B(\u_inFIFO/n209 ), .C(
        \u_inFIFO/currentState [0]), .D(\u_inFIFO/n225 ), .Q(\u_inFIFO/n239 )
         );
  OAI212 \u_inFIFO/U153  ( .A(\u_inFIFO/n238 ), .B(n986), .C(n1486), .Q(
        \u_inFIFO/N42 ) );
  OAI212 \u_inFIFO/U150  ( .A(\u_inFIFO/n235 ), .B(n980), .C(n1486), .Q(
        \u_inFIFO/N43 ) );
  OAI212 \u_inFIFO/U134  ( .A(n1485), .B(\u_inFIFO/n78 ), .C(\u_inFIFO/n222 ), 
        .Q(\u_inFIFO/n253 ) );
  OAI212 \u_inFIFO/U128  ( .A(n1485), .B(\u_inFIFO/n86 ), .C(\u_inFIFO/n216 ), 
        .Q(\u_inFIFO/n252 ) );
  OAI212 \u_inFIFO/U126  ( .A(n1485), .B(\u_inFIFO/n82 ), .C(\u_inFIFO/n215 ), 
        .Q(\u_inFIFO/n251 ) );
  OAI212 \u_inFIFO/U124  ( .A(n1485), .B(\u_inFIFO/n83 ), .C(\u_inFIFO/n214 ), 
        .Q(\u_inFIFO/n250 ) );
  OAI212 \u_inFIFO/U122  ( .A(n1485), .B(\u_inFIFO/n84 ), .C(\u_inFIFO/n213 ), 
        .Q(\u_inFIFO/n249 ) );
  OAI212 \u_inFIFO/U120  ( .A(n1485), .B(\u_inFIFO/n85 ), .C(\u_inFIFO/n210 ), 
        .Q(\u_inFIFO/n248 ) );
  OAI222 \u_inFIFO/U117  ( .A(\u_inFIFO/n111 ), .B(\u_inFIFO/n94 ), .C(
        \u_inFIFO/N38 ), .D(\u_inFIFO/n110 ), .Q(\u_inFIFO/n247 ) );
  OAI222 \u_inFIFO/U115  ( .A(\u_inFIFO/n111 ), .B(\u_inFIFO/n93 ), .C(
        \u_inFIFO/n208 ), .D(\u_inFIFO/n110 ), .Q(\u_inFIFO/n246 ) );
  OAI212 \u_inFIFO/U96  ( .A(\u_inFIFO/n193 ), .B(n966), .C(n967), .Q(
        \u_inFIFO/n192 ) );
  OAI212 \u_inFIFO/U90  ( .A(\u_inFIFO/n191 ), .B(n966), .C(n967), .Q(
        \u_inFIFO/n190 ) );
  OAI212 \u_inFIFO/U87  ( .A(\u_inFIFO/n189 ), .B(n966), .C(n967), .Q(
        \u_inFIFO/n188 ) );
  OAI212 \u_inFIFO/U84  ( .A(\u_inFIFO/n187 ), .B(n966), .C(n967), .Q(
        \u_inFIFO/n186 ) );
  OAI212 \u_inFIFO/U81  ( .A(\u_inFIFO/n185 ), .B(n966), .C(n967), .Q(
        \u_inFIFO/n184 ) );
  OAI212 \u_inFIFO/U78  ( .A(\u_inFIFO/n183 ), .B(n966), .C(n967), .Q(
        \u_inFIFO/n182 ) );
  OAI212 \u_inFIFO/U75  ( .A(\u_inFIFO/n181 ), .B(n966), .C(n967), .Q(
        \u_inFIFO/n180 ) );
  OAI212 \u_inFIFO/U72  ( .A(\u_inFIFO/n178 ), .B(n966), .C(n967), .Q(
        \u_inFIFO/n177 ) );
  OAI212 \u_inFIFO/U69  ( .A(\u_inFIFO/n176 ), .B(n966), .C(n967), .Q(
        \u_inFIFO/n175 ) );
  OAI212 \u_inFIFO/U67  ( .A(\u_inFIFO/n174 ), .B(n966), .C(n967), .Q(
        \u_inFIFO/n173 ) );
  OAI212 \u_inFIFO/U65  ( .A(\u_inFIFO/n172 ), .B(n966), .C(n967), .Q(
        \u_inFIFO/n171 ) );
  OAI212 \u_inFIFO/U63  ( .A(\u_inFIFO/n170 ), .B(n966), .C(n967), .Q(
        \u_inFIFO/n169 ) );
  OAI212 \u_inFIFO/U61  ( .A(\u_inFIFO/n168 ), .B(n966), .C(n967), .Q(
        \u_inFIFO/n167 ) );
  OAI212 \u_inFIFO/U59  ( .A(\u_inFIFO/n166 ), .B(n966), .C(n967), .Q(
        \u_inFIFO/n165 ) );
  OAI212 \u_inFIFO/U57  ( .A(\u_inFIFO/n164 ), .B(n966), .C(n967), .Q(
        \u_inFIFO/n163 ) );
  OAI212 \u_inFIFO/U55  ( .A(\u_inFIFO/n161 ), .B(n966), .C(n967), .Q(
        \u_inFIFO/n160 ) );
  OAI212 \u_inFIFO/U52  ( .A(\u_inFIFO/n159 ), .B(n966), .C(n967), .Q(
        \u_inFIFO/n158 ) );
  OAI212 \u_inFIFO/U50  ( .A(\u_inFIFO/n157 ), .B(\u_inFIFO/n118 ), .C(n967), 
        .Q(\u_inFIFO/n156 ) );
  OAI212 \u_inFIFO/U48  ( .A(\u_inFIFO/n155 ), .B(\u_inFIFO/n118 ), .C(n967), 
        .Q(\u_inFIFO/n154 ) );
  OAI212 \u_inFIFO/U46  ( .A(\u_inFIFO/n153 ), .B(\u_inFIFO/n118 ), .C(n967), 
        .Q(\u_inFIFO/n152 ) );
  OAI212 \u_inFIFO/U44  ( .A(\u_inFIFO/n151 ), .B(n966), .C(n967), .Q(
        \u_inFIFO/n150 ) );
  OAI212 \u_inFIFO/U42  ( .A(\u_inFIFO/n149 ), .B(n966), .C(n967), .Q(
        \u_inFIFO/n148 ) );
  OAI212 \u_inFIFO/U40  ( .A(\u_inFIFO/n147 ), .B(n966), .C(n967), .Q(
        \u_inFIFO/n146 ) );
  OAI212 \u_inFIFO/U38  ( .A(\u_inFIFO/n144 ), .B(n966), .C(n967), .Q(
        \u_inFIFO/n143 ) );
  OAI212 \u_inFIFO/U35  ( .A(\u_inFIFO/n141 ), .B(\u_inFIFO/n118 ), .C(
        \u_inFIFO/n119 ), .Q(\u_inFIFO/n140 ) );
  OAI212 \u_inFIFO/U33  ( .A(\u_inFIFO/n138 ), .B(\u_inFIFO/n118 ), .C(
        \u_inFIFO/n119 ), .Q(\u_inFIFO/n137 ) );
  OAI212 \u_inFIFO/U31  ( .A(\u_inFIFO/n135 ), .B(\u_inFIFO/n118 ), .C(
        \u_inFIFO/n119 ), .Q(\u_inFIFO/n134 ) );
  OAI212 \u_inFIFO/U29  ( .A(\u_inFIFO/n132 ), .B(\u_inFIFO/n118 ), .C(
        \u_inFIFO/n119 ), .Q(\u_inFIFO/n131 ) );
  OAI212 \u_inFIFO/U27  ( .A(\u_inFIFO/n129 ), .B(\u_inFIFO/n118 ), .C(
        \u_inFIFO/n119 ), .Q(\u_inFIFO/n128 ) );
  OAI212 \u_inFIFO/U25  ( .A(\u_inFIFO/n126 ), .B(\u_inFIFO/n118 ), .C(
        \u_inFIFO/n119 ), .Q(\u_inFIFO/n125 ) );
  OAI212 \u_inFIFO/U23  ( .A(\u_inFIFO/n123 ), .B(\u_inFIFO/n118 ), .C(
        \u_inFIFO/n119 ), .Q(\u_inFIFO/n122 ) );
  OAI212 \u_inFIFO/U21  ( .A(\u_inFIFO/n117 ), .B(\u_inFIFO/n118 ), .C(n967), 
        .Q(\u_inFIFO/n112 ) );
  OAI222 \u_inFIFO/U20  ( .A(n233), .B(\u_inFIFO/n110 ), .C(\u_inFIFO/n96 ), 
        .D(\u_inFIFO/n111 ), .Q(\u_inFIFO/n245 ) );
  OAI222 \u_coder/U200  ( .A(\u_coder/N1149 ), .B(\u_coder/n148 ), .C(
        \u_coder/n234 ), .D(\u_coder/n313 ), .Q(\u_coder/n374 ) );
  OAI212 \u_coder/U187  ( .A(\u_coder/IorQ ), .B(\u_coder/n307 ), .C(
        \u_coder/n308 ), .Q(\u_coder/n373 ) );
  OAI222 \u_coder/U184  ( .A(\u_coder/N1143 ), .B(\u_coder/n147 ), .C(
        \u_coder/n189 ), .D(\u_coder/n306 ), .Q(\u_coder/n372 ) );
  OAI212 \u_coder/U157  ( .A(\u_coder/n200 ), .B(n2275), .C(\u_coder/n256 ), 
        .Q(\u_coder/n282 ) );
  OAI222 \u_coder/U155  ( .A(n809), .B(\u_coder/n90 ), .C(n808), .D(n368), .Q(
        \u_coder/n371 ) );
  OAI222 \u_coder/U154  ( .A(\u_coder/n138 ), .B(n809), .C(\u_coder/n283 ), 
        .D(n777), .Q(\u_coder/n370 ) );
  OAI222 \u_coder/U153  ( .A(\u_coder/n137 ), .B(n809), .C(n808), .D(n1745), 
        .Q(\u_coder/n369 ) );
  OAI222 \u_coder/U152  ( .A(\u_coder/n135 ), .B(n809), .C(\u_coder/n283 ), 
        .D(n1744), .Q(\u_coder/n368 ) );
  OAI222 \u_coder/U151  ( .A(\u_coder/n134 ), .B(n809), .C(n808), .D(n1743), 
        .Q(\u_coder/n367 ) );
  OAI222 \u_coder/U150  ( .A(n809), .B(\u_coder/n131 ), .C(\u_coder/n283 ), 
        .D(n1742), .Q(\u_coder/n366 ) );
  OAI222 \u_coder/U149  ( .A(n809), .B(\u_coder/n130 ), .C(n808), .D(n1741), 
        .Q(\u_coder/n365 ) );
  OAI222 \u_coder/U148  ( .A(n809), .B(\u_coder/n129 ), .C(\u_coder/n283 ), 
        .D(n1740), .Q(\u_coder/n364 ) );
  OAI222 \u_coder/U147  ( .A(n809), .B(\u_coder/n128 ), .C(n808), .D(n1739), 
        .Q(\u_coder/n363 ) );
  OAI222 \u_coder/U146  ( .A(n809), .B(\u_coder/n127 ), .C(\u_coder/n283 ), 
        .D(n1738), .Q(\u_coder/n362 ) );
  OAI222 \u_coder/U145  ( .A(n809), .B(\u_coder/n126 ), .C(n808), .D(n1737), 
        .Q(\u_coder/n361 ) );
  OAI222 \u_coder/U144  ( .A(n809), .B(\u_coder/n125 ), .C(\u_coder/n283 ), 
        .D(n1736), .Q(\u_coder/n360 ) );
  OAI222 \u_coder/U143  ( .A(n809), .B(\u_coder/n124 ), .C(n808), .D(n1735), 
        .Q(\u_coder/n359 ) );
  OAI222 \u_coder/U142  ( .A(n809), .B(\u_coder/n123 ), .C(\u_coder/n283 ), 
        .D(n1734), .Q(\u_coder/n358 ) );
  OAI222 \u_coder/U141  ( .A(n809), .B(\u_coder/n122 ), .C(n808), .D(n1733), 
        .Q(\u_coder/n357 ) );
  OAI222 \u_coder/U140  ( .A(n809), .B(\u_coder/n121 ), .C(\u_coder/n283 ), 
        .D(n1732), .Q(\u_coder/n356 ) );
  OAI222 \u_coder/U139  ( .A(n809), .B(\u_coder/n120 ), .C(n808), .D(n1731), 
        .Q(\u_coder/n355 ) );
  OAI222 \u_coder/U138  ( .A(n809), .B(\u_coder/n119 ), .C(\u_coder/n283 ), 
        .D(n1730), .Q(\u_coder/n354 ) );
  OAI222 \u_coder/U137  ( .A(n809), .B(\u_coder/n118 ), .C(n808), .D(n1729), 
        .Q(\u_coder/n353 ) );
  OAI222 \u_coder/U136  ( .A(n809), .B(\u_coder/n117 ), .C(\u_coder/n283 ), 
        .D(n1728), .Q(\u_coder/n352 ) );
  OAI212 \u_coder/U133  ( .A(\u_coder/n278 ), .B(\u_coder/n161 ), .C(
        \u_coder/n279 ), .Q(\u_coder/n276 ) );
  OAI222 \u_coder/U131  ( .A(\u_coder/n276 ), .B(\u_coder/n277 ), .C(n1713), 
        .D(n2687), .Q(\u_coder/n351 ) );
  OAI222 \u_coder/U124  ( .A(\u_coder/n141 ), .B(\u_coder/n273 ), .C(
        \u_coder/n195 ), .D(\u_coder/n186 ), .Q(\u_coder/n350 ) );
  OAI222 \u_coder/U123  ( .A(\u_coder/n140 ), .B(\u_coder/n274 ), .C(
        \u_coder/n141 ), .D(n1660), .Q(\u_coder/n349 ) );
  OAI212 \u_coder/U120  ( .A(\u_coder/n196 ), .B(\u_coder/n266 ), .C(n1724), 
        .Q(\u_coder/n272 ) );
  OAI212 \u_coder/U110  ( .A(\u_coder/n263 ), .B(\u_coder/n161 ), .C(
        \u_coder/n264 ), .Q(\u_coder/n345 ) );
  OAI222 \u_coder/U99  ( .A(\u_coder/n144 ), .B(n1473), .C(\u_coder/n212 ), 
        .D(\u_coder/n230 ), .Q(\u_coder/n343 ) );
  OAI212 \u_coder/U96  ( .A(n1749), .B(\u_coder/n247 ), .C(n1756), .Q(
        \u_coder/n253 ) );
  OAI212 \u_coder/U86  ( .A(\u_coder/n244 ), .B(\u_coder/n200 ), .C(
        \u_coder/n245 ), .Q(\u_coder/n339 ) );
  OAI212 \u_coder/U73  ( .A(\u_coder/n211 ), .B(n1711), .C(\u_coder/n239 ), 
        .Q(\u_coder/n238 ) );
  OAI212 \u_coder/U72  ( .A(\u_coder/n201 ), .B(n1750), .C(\u_coder/n238 ), 
        .Q(\u_coder/n236 ) );
  OAI212 \u_coder/U64  ( .A(\u_coder/n138 ), .B(\u_coder/n137 ), .C(
        \u_coder/j [2]), .Q(\u_coder/n222 ) );
  OAI212 \u_coder/U59  ( .A(\u_coder/n217 ), .B(\u_coder/n209 ), .C(
        \u_coder/n221 ), .Q(\u_coder/n215 ) );
  OAI222 \u_coder/U58  ( .A(\u_coder/n217 ), .B(n1707), .C(n1727), .D(n1706), 
        .Q(\u_coder/n216 ) );
  OAI212 \u_coder/U52  ( .A(\u_coder/n207 ), .B(\u_coder/n209 ), .C(
        \u_coder/n210 ), .Q(\u_coder/n204 ) );
  OAI222 \u_coder/U51  ( .A(\u_coder/n207 ), .B(n1707), .C(\u_coder/n208 ), 
        .D(n1706), .Q(\u_coder/n206 ) );
  OAI222 \u_coder/U47  ( .A(n1707), .B(n1661), .C(\u_coder/n200 ), .D(
        \u_coder/n201 ), .Q(\u_coder/n199 ) );
  OAI212 \u_coder/U35  ( .A(n1709), .B(\u_coder/n176 ), .C(\u_coder/n194 ), 
        .Q(\u_coder/n193 ) );
  OAI212 \u_coder/U34  ( .A(\u_coder/n156 ), .B(n1719), .C(\u_coder/n193 ), 
        .Q(\u_coder/n192 ) );
  OAI212 \u_coder/U31  ( .A(\u_coder/n161 ), .B(\u_coder/n188 ), .C(n978), .Q(
        \u_coder/n187 ) );
  OAI212 \u_coder/U27  ( .A(\u_coder/n89 ), .B(\u_coder/n88 ), .C(
        \u_coder/i [2]), .Q(\u_coder/n179 ) );
  OAI222 \u_coder/U20  ( .A(n1715), .B(n1708), .C(\u_coder/n166 ), .D(
        \u_coder/n167 ), .Q(\u_coder/n174 ) );
  OAI222 \u_coder/U18  ( .A(\u_coder/n171 ), .B(n1660), .C(\u_coder/n172 ), 
        .D(\u_coder/n161 ), .Q(\u_coder/n170 ) );
  OAI222 \u_coder/U14  ( .A(\u_coder/n165 ), .B(n1708), .C(\u_coder/n166 ), 
        .D(\u_coder/n167 ), .Q(\u_coder/n164 ) );
  OAI222 \u_coder/U12  ( .A(\u_coder/n159 ), .B(n1660), .C(\u_coder/n160 ), 
        .D(\u_coder/n161 ), .Q(\u_coder/n158 ) );
  OAI212 \u_coder/U5  ( .A(\u_coder/n152 ), .B(\u_coder/n146 ), .C(
        \u_coder/n153 ), .Q(\u_coder/n333 ) );
  OAI212 \u_cordic/U24  ( .A(\u_cordic/n13 ), .B(n1663), .C(n1777), .Q(
        \u_cordic/n34 ) );
  OAI212 \u_cordic/U5  ( .A(\u_cordic/present_state [1]), .B(n1778), .C(
        \sig_MUX_inMUX14[0] ), .Q(\u_cordic/n16 ) );
  OAI222 \u_cdr/U35  ( .A(n294), .B(\u_cdr/n43 ), .C(n1785), .D(\u_cdr/n46 ), 
        .Q(\u_cdr/n58 ) );
  OAI222 \u_cdr/U34  ( .A(n3), .B(\u_cdr/n43 ), .C(n358), .D(\u_cdr/n46 ), .Q(
        \u_cdr/n57 ) );
  OAI222 \u_cdr/U33  ( .A(n295), .B(\u_cdr/n43 ), .C(n359), .D(\u_cdr/n46 ), 
        .Q(\u_cdr/n56 ) );
  OAI222 \u_cdr/U32  ( .A(\u_cdr/n43 ), .B(n36), .C(\u_cdr/n45 ), .D(
        \u_cdr/n46 ), .Q(\u_cdr/n55 ) );
  OAI212 \u_cdr/U25  ( .A(\u_cdr/n42 ), .B(n986), .C(\u_cdr/n43 ), .Q(
        \u_cdr/n26 ) );
  OAI222 \u_cdr/U23  ( .A(\u_cdr/cnt_d [0]), .B(\u_cdr/n23 ), .C(\u_cdr/n41 ), 
        .D(\u_cdr/n15 ), .Q(\u_cdr/n54 ) );
  OAI222 \u_cdr/U22  ( .A(n981), .B(\u_cdr/n14 ), .C(\u_cdr/n23 ), .D(
        \u_cdr/n15 ), .Q(\u_cdr/n53 ) );
  OAI212 \u_cdr/U15  ( .A(\u_cdr/cnt [0]), .B(n1470), .C(\u_cdr/n34 ), .Q(
        \u_cdr/n33 ) );
  OAI212 \u_cdr/U12  ( .A(\u_cdr/n35 ), .B(\u_cdr/n16 ), .C(\u_cdr/n36 ), .Q(
        \u_cdr/n51 ) );
  OAI212 \u_cdr/U10  ( .A(n1469), .B(\u_cdr/n17 ), .C(\u_cdr/n31 ), .Q(
        \u_cdr/n50 ) );
  OAI212 \u_cdr/U5  ( .A(\u_cdr/n25 ), .B(\u_cdr/n26 ), .C(\u_cdr/dir ), .Q(
        \u_cdr/n24 ) );
  OAI212 \u_outFIFO/U495  ( .A(\u_outFIFO/currentState [1]), .B(
        \u_outFIFO/n525 ), .C(\u_outFIFO/n544 ), .Q(\u_outFIFO/n549 ) );
  OAI212 \u_outFIFO/U494  ( .A(\u_outFIFO/n548 ), .B(n982), .C(n1585), .Q(
        \u_outFIFO/N41 ) );
  OAI212 \u_outFIFO/U488  ( .A(\u_outFIFO/n543 ), .B(n985), .C(
        \u_outFIFO/n544 ), .Q(\u_outFIFO/N42 ) );
  OAI222 \u_outFIFO/U487  ( .A(\u_outFIFO/N473 ), .B(n1788), .C(n1792), .D(
        n1789), .Q(\u_outFIFO/n542 ) );
  OAI212 \u_outFIFO/U485  ( .A(\u_outFIFO/n541 ), .B(n986), .C(n1585), .Q(
        \u_outFIFO/N43 ) );
  OAI222 \u_outFIFO/U478  ( .A(\u_outFIFO/n194 ), .B(n1468), .C(
        \u_outFIFO/n533 ), .D(\u_outFIFO/i_FIFO [0]), .Q(\u_outFIFO/n690 ) );
  OAI222 \u_outFIFO/U477  ( .A(\u_outFIFO/n193 ), .B(n1468), .C(
        \u_outFIFO/n533 ), .D(n1799), .Q(\u_outFIFO/n689 ) );
  OAI222 \u_outFIFO/U476  ( .A(\u_outFIFO/n192 ), .B(n1468), .C(
        \u_outFIFO/n533 ), .D(n1798), .Q(\u_outFIFO/n688 ) );
  OAI222 \u_outFIFO/U475  ( .A(\u_outFIFO/n191 ), .B(n1468), .C(
        \u_outFIFO/n533 ), .D(n1797), .Q(\u_outFIFO/n687 ) );
  OAI222 \u_outFIFO/U474  ( .A(\u_outFIFO/n185 ), .B(n1468), .C(
        \u_outFIFO/n533 ), .D(n380), .Q(\u_outFIFO/n686 ) );
  AOI212 \u_outFIFO/U470  ( .A(\u_outFIFO/n206 ), .B(\u_outFIFO/n530 ), .C(
        \u_outFIFO/n527 ), .Q(\u_outFIFO/n512 ) );
  OAI212 \u_outFIFO/U466  ( .A(\u_outFIFO/n512 ), .B(\u_outFIFO/n178 ), .C(
        \u_outFIFO/n528 ), .Q(\u_outFIFO/n685 ) );
  OAI212 \u_outFIFO/U457  ( .A(\u_outFIFO/n512 ), .B(\u_outFIFO/n184 ), .C(
        \u_outFIFO/n518 ), .Q(\u_outFIFO/n684 ) );
  OAI212 \u_outFIFO/U455  ( .A(\u_outFIFO/n512 ), .B(\u_outFIFO/n183 ), .C(
        \u_outFIFO/n517 ), .Q(\u_outFIFO/n683 ) );
  OAI212 \u_outFIFO/U453  ( .A(\u_outFIFO/n512 ), .B(\u_outFIFO/n182 ), .C(
        \u_outFIFO/n516 ), .Q(\u_outFIFO/n682 ) );
  OAI212 \u_outFIFO/U451  ( .A(\u_outFIFO/n512 ), .B(\u_outFIFO/n181 ), .C(
        \u_outFIFO/n515 ), .Q(\u_outFIFO/n681 ) );
  OAI212 \u_outFIFO/U449  ( .A(\u_outFIFO/n512 ), .B(\u_outFIFO/n180 ), .C(
        \u_outFIFO/n513 ), .Q(\u_outFIFO/n680 ) );
  OAI222 \u_outFIFO/U443  ( .A(\u_outFIFO/n195 ), .B(n958), .C(
        \u_outFIFO/n510 ), .D(\u_outFIFO/n502 ), .Q(\u_outFIFO/n679 ) );
  OAI212 \u_outFIFO/U431  ( .A(n806), .B(\u_outFIFO/n444 ), .C(n830), .Q(
        \u_outFIFO/n501 ) );
  OAI212 \u_outFIFO/U429  ( .A(n1459), .B(n948), .C(\u_outFIFO/FIFO[31][3] ), 
        .Q(\u_outFIFO/n500 ) );
  OAI212 \u_outFIFO/U428  ( .A(n1459), .B(n946), .C(\u_outFIFO/n500 ), .Q(
        \u_outFIFO/n678 ) );
  OAI212 \u_outFIFO/U426  ( .A(n806), .B(\u_outFIFO/n441 ), .C(n830), .Q(
        \u_outFIFO/n499 ) );
  OAI212 \u_outFIFO/U425  ( .A(n1458), .B(n948), .C(\u_outFIFO/FIFO[31][2] ), 
        .Q(\u_outFIFO/n498 ) );
  OAI212 \u_outFIFO/U424  ( .A(n1458), .B(n946), .C(\u_outFIFO/n498 ), .Q(
        \u_outFIFO/n677 ) );
  OAI212 \u_outFIFO/U422  ( .A(n806), .B(\u_outFIFO/n438 ), .C(n830), .Q(
        \u_outFIFO/n497 ) );
  OAI212 \u_outFIFO/U421  ( .A(n1457), .B(n948), .C(\u_outFIFO/FIFO[31][1] ), 
        .Q(\u_outFIFO/n496 ) );
  OAI212 \u_outFIFO/U420  ( .A(n1457), .B(n944), .C(\u_outFIFO/n496 ), .Q(
        \u_outFIFO/n676 ) );
  OAI212 \u_outFIFO/U418  ( .A(n806), .B(\u_outFIFO/n435 ), .C(n830), .Q(
        \u_outFIFO/n494 ) );
  OAI212 \u_outFIFO/U417  ( .A(n1456), .B(n948), .C(\u_outFIFO/FIFO[31][0] ), 
        .Q(\u_outFIFO/n493 ) );
  OAI212 \u_outFIFO/U416  ( .A(n1456), .B(n944), .C(\u_outFIFO/n493 ), .Q(
        \u_outFIFO/n675 ) );
  OAI212 \u_outFIFO/U414  ( .A(n803), .B(\u_outFIFO/n444 ), .C(n830), .Q(
        \u_outFIFO/n492 ) );
  OAI212 \u_outFIFO/U413  ( .A(n1455), .B(n948), .C(\u_outFIFO/FIFO[30][3] ), 
        .Q(\u_outFIFO/n491 ) );
  OAI212 \u_outFIFO/U412  ( .A(n1455), .B(n946), .C(\u_outFIFO/n491 ), .Q(
        \u_outFIFO/n674 ) );
  OAI212 \u_outFIFO/U411  ( .A(n803), .B(\u_outFIFO/n441 ), .C(n830), .Q(
        \u_outFIFO/n490 ) );
  OAI212 \u_outFIFO/U410  ( .A(n1454), .B(n948), .C(\u_outFIFO/FIFO[30][2] ), 
        .Q(\u_outFIFO/n489 ) );
  OAI212 \u_outFIFO/U409  ( .A(n1454), .B(n946), .C(\u_outFIFO/n489 ), .Q(
        \u_outFIFO/n673 ) );
  OAI212 \u_outFIFO/U408  ( .A(n803), .B(\u_outFIFO/n438 ), .C(n830), .Q(
        \u_outFIFO/n488 ) );
  OAI212 \u_outFIFO/U407  ( .A(n1453), .B(n948), .C(\u_outFIFO/FIFO[30][1] ), 
        .Q(\u_outFIFO/n487 ) );
  OAI212 \u_outFIFO/U406  ( .A(n1453), .B(n945), .C(\u_outFIFO/n487 ), .Q(
        \u_outFIFO/n672 ) );
  OAI212 \u_outFIFO/U405  ( .A(n803), .B(\u_outFIFO/n435 ), .C(n830), .Q(
        \u_outFIFO/n486 ) );
  OAI212 \u_outFIFO/U404  ( .A(n1452), .B(n948), .C(\u_outFIFO/FIFO[30][0] ), 
        .Q(\u_outFIFO/n485 ) );
  OAI212 \u_outFIFO/U403  ( .A(n1452), .B(n945), .C(\u_outFIFO/n485 ), .Q(
        \u_outFIFO/n671 ) );
  OAI212 \u_outFIFO/U401  ( .A(n801), .B(\u_outFIFO/n444 ), .C(n829), .Q(
        \u_outFIFO/n484 ) );
  OAI212 \u_outFIFO/U400  ( .A(n1451), .B(n948), .C(\u_outFIFO/FIFO[29][3] ), 
        .Q(\u_outFIFO/n483 ) );
  OAI212 \u_outFIFO/U399  ( .A(n1451), .B(n945), .C(\u_outFIFO/n483 ), .Q(
        \u_outFIFO/n670 ) );
  OAI212 \u_outFIFO/U398  ( .A(n801), .B(\u_outFIFO/n441 ), .C(n829), .Q(
        \u_outFIFO/n482 ) );
  OAI212 \u_outFIFO/U397  ( .A(n1450), .B(n948), .C(\u_outFIFO/FIFO[29][2] ), 
        .Q(\u_outFIFO/n481 ) );
  OAI212 \u_outFIFO/U396  ( .A(n1450), .B(n944), .C(\u_outFIFO/n481 ), .Q(
        \u_outFIFO/n669 ) );
  OAI212 \u_outFIFO/U395  ( .A(n801), .B(\u_outFIFO/n438 ), .C(n829), .Q(
        \u_outFIFO/n480 ) );
  OAI212 \u_outFIFO/U394  ( .A(n1449), .B(n948), .C(\u_outFIFO/FIFO[29][1] ), 
        .Q(\u_outFIFO/n479 ) );
  OAI212 \u_outFIFO/U393  ( .A(n1449), .B(n944), .C(\u_outFIFO/n479 ), .Q(
        \u_outFIFO/n668 ) );
  OAI212 \u_outFIFO/U392  ( .A(n801), .B(\u_outFIFO/n435 ), .C(n829), .Q(
        \u_outFIFO/n478 ) );
  OAI212 \u_outFIFO/U391  ( .A(n1448), .B(n948), .C(\u_outFIFO/FIFO[29][0] ), 
        .Q(\u_outFIFO/n477 ) );
  OAI212 \u_outFIFO/U390  ( .A(n1448), .B(n944), .C(\u_outFIFO/n477 ), .Q(
        \u_outFIFO/n667 ) );
  OAI212 \u_outFIFO/U388  ( .A(n799), .B(\u_outFIFO/n444 ), .C(n829), .Q(
        \u_outFIFO/n476 ) );
  OAI212 \u_outFIFO/U387  ( .A(n1447), .B(n948), .C(\u_outFIFO/FIFO[28][3] ), 
        .Q(\u_outFIFO/n475 ) );
  OAI212 \u_outFIFO/U386  ( .A(n1447), .B(n945), .C(\u_outFIFO/n475 ), .Q(
        \u_outFIFO/n666 ) );
  OAI212 \u_outFIFO/U385  ( .A(n799), .B(\u_outFIFO/n441 ), .C(n829), .Q(
        \u_outFIFO/n474 ) );
  OAI212 \u_outFIFO/U384  ( .A(n1446), .B(n949), .C(\u_outFIFO/FIFO[28][2] ), 
        .Q(\u_outFIFO/n473 ) );
  OAI212 \u_outFIFO/U383  ( .A(n1446), .B(n944), .C(\u_outFIFO/n473 ), .Q(
        \u_outFIFO/n665 ) );
  OAI212 \u_outFIFO/U382  ( .A(n799), .B(\u_outFIFO/n438 ), .C(n829), .Q(
        \u_outFIFO/n472 ) );
  OAI212 \u_outFIFO/U381  ( .A(n1445), .B(n949), .C(\u_outFIFO/FIFO[28][1] ), 
        .Q(\u_outFIFO/n471 ) );
  OAI212 \u_outFIFO/U380  ( .A(n1445), .B(n946), .C(\u_outFIFO/n471 ), .Q(
        \u_outFIFO/n664 ) );
  OAI212 \u_outFIFO/U379  ( .A(n799), .B(\u_outFIFO/n435 ), .C(n829), .Q(
        \u_outFIFO/n470 ) );
  OAI212 \u_outFIFO/U378  ( .A(n1444), .B(n949), .C(\u_outFIFO/FIFO[28][0] ), 
        .Q(\u_outFIFO/n469 ) );
  OAI212 \u_outFIFO/U377  ( .A(n1444), .B(n945), .C(\u_outFIFO/n469 ), .Q(
        \u_outFIFO/n663 ) );
  OAI212 \u_outFIFO/U375  ( .A(n797), .B(\u_outFIFO/n444 ), .C(n828), .Q(
        \u_outFIFO/n468 ) );
  OAI212 \u_outFIFO/U374  ( .A(n1443), .B(n949), .C(\u_outFIFO/FIFO[27][3] ), 
        .Q(\u_outFIFO/n467 ) );
  OAI212 \u_outFIFO/U373  ( .A(n1443), .B(n945), .C(\u_outFIFO/n467 ), .Q(
        \u_outFIFO/n662 ) );
  OAI212 \u_outFIFO/U372  ( .A(n797), .B(\u_outFIFO/n441 ), .C(n828), .Q(
        \u_outFIFO/n466 ) );
  OAI212 \u_outFIFO/U371  ( .A(n1442), .B(n949), .C(\u_outFIFO/FIFO[27][2] ), 
        .Q(\u_outFIFO/n465 ) );
  OAI212 \u_outFIFO/U370  ( .A(n1442), .B(n944), .C(\u_outFIFO/n465 ), .Q(
        \u_outFIFO/n661 ) );
  OAI212 \u_outFIFO/U369  ( .A(n797), .B(\u_outFIFO/n438 ), .C(n828), .Q(
        \u_outFIFO/n464 ) );
  OAI212 \u_outFIFO/U368  ( .A(n1441), .B(n949), .C(\u_outFIFO/FIFO[27][1] ), 
        .Q(\u_outFIFO/n463 ) );
  OAI212 \u_outFIFO/U367  ( .A(n1441), .B(n946), .C(\u_outFIFO/n463 ), .Q(
        \u_outFIFO/n660 ) );
  OAI212 \u_outFIFO/U366  ( .A(n797), .B(\u_outFIFO/n435 ), .C(n828), .Q(
        \u_outFIFO/n462 ) );
  OAI212 \u_outFIFO/U365  ( .A(n1440), .B(n949), .C(\u_outFIFO/FIFO[27][0] ), 
        .Q(\u_outFIFO/n461 ) );
  OAI212 \u_outFIFO/U364  ( .A(n1440), .B(n945), .C(\u_outFIFO/n461 ), .Q(
        \u_outFIFO/n659 ) );
  OAI212 \u_outFIFO/U362  ( .A(n795), .B(\u_outFIFO/n444 ), .C(n828), .Q(
        \u_outFIFO/n460 ) );
  OAI212 \u_outFIFO/U361  ( .A(n1439), .B(n949), .C(\u_outFIFO/FIFO[26][3] ), 
        .Q(\u_outFIFO/n459 ) );
  OAI212 \u_outFIFO/U360  ( .A(n1439), .B(n944), .C(\u_outFIFO/n459 ), .Q(
        \u_outFIFO/n658 ) );
  OAI212 \u_outFIFO/U359  ( .A(n795), .B(\u_outFIFO/n441 ), .C(n828), .Q(
        \u_outFIFO/n458 ) );
  OAI212 \u_outFIFO/U358  ( .A(n1438), .B(n949), .C(\u_outFIFO/FIFO[26][2] ), 
        .Q(\u_outFIFO/n457 ) );
  OAI212 \u_outFIFO/U357  ( .A(n1438), .B(n944), .C(\u_outFIFO/n457 ), .Q(
        \u_outFIFO/n657 ) );
  OAI212 \u_outFIFO/U356  ( .A(n795), .B(\u_outFIFO/n438 ), .C(n828), .Q(
        \u_outFIFO/n456 ) );
  OAI212 \u_outFIFO/U355  ( .A(n1437), .B(n949), .C(\u_outFIFO/FIFO[26][1] ), 
        .Q(\u_outFIFO/n455 ) );
  OAI212 \u_outFIFO/U354  ( .A(n1437), .B(n946), .C(\u_outFIFO/n455 ), .Q(
        \u_outFIFO/n656 ) );
  OAI212 \u_outFIFO/U353  ( .A(n795), .B(\u_outFIFO/n435 ), .C(n828), .Q(
        \u_outFIFO/n454 ) );
  OAI212 \u_outFIFO/U352  ( .A(n1436), .B(n949), .C(\u_outFIFO/FIFO[26][0] ), 
        .Q(\u_outFIFO/n453 ) );
  OAI212 \u_outFIFO/U351  ( .A(n1436), .B(n945), .C(\u_outFIFO/n453 ), .Q(
        \u_outFIFO/n655 ) );
  OAI212 \u_outFIFO/U349  ( .A(n793), .B(\u_outFIFO/n444 ), .C(n827), .Q(
        \u_outFIFO/n452 ) );
  OAI212 \u_outFIFO/U348  ( .A(n1435), .B(n949), .C(\u_outFIFO/FIFO[25][3] ), 
        .Q(\u_outFIFO/n451 ) );
  OAI212 \u_outFIFO/U347  ( .A(n1435), .B(n946), .C(\u_outFIFO/n451 ), .Q(
        \u_outFIFO/n654 ) );
  OAI212 \u_outFIFO/U346  ( .A(n793), .B(\u_outFIFO/n441 ), .C(n827), .Q(
        \u_outFIFO/n450 ) );
  OAI212 \u_outFIFO/U345  ( .A(n1434), .B(n949), .C(\u_outFIFO/FIFO[25][2] ), 
        .Q(\u_outFIFO/n449 ) );
  OAI212 \u_outFIFO/U344  ( .A(n1434), .B(n944), .C(\u_outFIFO/n449 ), .Q(
        \u_outFIFO/n653 ) );
  OAI212 \u_outFIFO/U343  ( .A(n793), .B(\u_outFIFO/n438 ), .C(n827), .Q(
        \u_outFIFO/n448 ) );
  OAI212 \u_outFIFO/U342  ( .A(n1433), .B(n950), .C(\u_outFIFO/FIFO[25][1] ), 
        .Q(\u_outFIFO/n447 ) );
  OAI212 \u_outFIFO/U341  ( .A(n1433), .B(n944), .C(\u_outFIFO/n447 ), .Q(
        \u_outFIFO/n652 ) );
  OAI212 \u_outFIFO/U340  ( .A(n793), .B(\u_outFIFO/n435 ), .C(n827), .Q(
        \u_outFIFO/n446 ) );
  OAI212 \u_outFIFO/U339  ( .A(n1432), .B(n950), .C(\u_outFIFO/FIFO[25][0] ), 
        .Q(\u_outFIFO/n445 ) );
  OAI212 \u_outFIFO/U338  ( .A(n1432), .B(n944), .C(\u_outFIFO/n445 ), .Q(
        \u_outFIFO/n651 ) );
  OAI212 \u_outFIFO/U336  ( .A(n791), .B(\u_outFIFO/n444 ), .C(n827), .Q(
        \u_outFIFO/n443 ) );
  OAI212 \u_outFIFO/U335  ( .A(n1431), .B(n950), .C(\u_outFIFO/FIFO[24][3] ), 
        .Q(\u_outFIFO/n442 ) );
  OAI212 \u_outFIFO/U334  ( .A(n1431), .B(n944), .C(\u_outFIFO/n442 ), .Q(
        \u_outFIFO/n650 ) );
  OAI212 \u_outFIFO/U333  ( .A(n791), .B(\u_outFIFO/n441 ), .C(n827), .Q(
        \u_outFIFO/n440 ) );
  OAI212 \u_outFIFO/U332  ( .A(n1430), .B(n950), .C(\u_outFIFO/FIFO[24][2] ), 
        .Q(\u_outFIFO/n439 ) );
  OAI212 \u_outFIFO/U331  ( .A(n1430), .B(n944), .C(\u_outFIFO/n439 ), .Q(
        \u_outFIFO/n649 ) );
  OAI212 \u_outFIFO/U330  ( .A(n791), .B(\u_outFIFO/n438 ), .C(n827), .Q(
        \u_outFIFO/n437 ) );
  OAI212 \u_outFIFO/U329  ( .A(n1429), .B(n950), .C(\u_outFIFO/FIFO[24][1] ), 
        .Q(\u_outFIFO/n436 ) );
  OAI212 \u_outFIFO/U328  ( .A(n1429), .B(n944), .C(\u_outFIFO/n436 ), .Q(
        \u_outFIFO/n648 ) );
  OAI212 \u_outFIFO/U327  ( .A(n791), .B(\u_outFIFO/n435 ), .C(n827), .Q(
        \u_outFIFO/n434 ) );
  OAI212 \u_outFIFO/U326  ( .A(n1428), .B(n950), .C(\u_outFIFO/FIFO[24][0] ), 
        .Q(\u_outFIFO/n433 ) );
  OAI212 \u_outFIFO/U325  ( .A(n1428), .B(n944), .C(\u_outFIFO/n433 ), .Q(
        \u_outFIFO/n647 ) );
  OAI212 \u_outFIFO/U322  ( .A(n807), .B(\u_outFIFO/n375 ), .C(n826), .Q(
        \u_outFIFO/n432 ) );
  OAI212 \u_outFIFO/U321  ( .A(n1427), .B(n950), .C(\u_outFIFO/FIFO[23][3] ), 
        .Q(\u_outFIFO/n431 ) );
  OAI212 \u_outFIFO/U320  ( .A(n1427), .B(n944), .C(\u_outFIFO/n431 ), .Q(
        \u_outFIFO/n646 ) );
  OAI212 \u_outFIFO/U318  ( .A(n807), .B(\u_outFIFO/n372 ), .C(n826), .Q(
        \u_outFIFO/n430 ) );
  OAI212 \u_outFIFO/U317  ( .A(n1426), .B(n950), .C(\u_outFIFO/FIFO[23][2] ), 
        .Q(\u_outFIFO/n429 ) );
  OAI212 \u_outFIFO/U316  ( .A(n1426), .B(n944), .C(\u_outFIFO/n429 ), .Q(
        \u_outFIFO/n645 ) );
  OAI212 \u_outFIFO/U314  ( .A(n807), .B(\u_outFIFO/n369 ), .C(n826), .Q(
        \u_outFIFO/n428 ) );
  OAI212 \u_outFIFO/U313  ( .A(n1425), .B(n950), .C(\u_outFIFO/FIFO[23][1] ), 
        .Q(\u_outFIFO/n427 ) );
  OAI212 \u_outFIFO/U312  ( .A(n1425), .B(n944), .C(\u_outFIFO/n427 ), .Q(
        \u_outFIFO/n644 ) );
  OAI212 \u_outFIFO/U310  ( .A(n807), .B(\u_outFIFO/n366 ), .C(n826), .Q(
        \u_outFIFO/n425 ) );
  OAI212 \u_outFIFO/U309  ( .A(n1424), .B(n950), .C(\u_outFIFO/FIFO[23][0] ), 
        .Q(\u_outFIFO/n424 ) );
  OAI212 \u_outFIFO/U308  ( .A(n1424), .B(n944), .C(\u_outFIFO/n424 ), .Q(
        \u_outFIFO/n643 ) );
  OAI212 \u_outFIFO/U307  ( .A(n804), .B(\u_outFIFO/n375 ), .C(n826), .Q(
        \u_outFIFO/n423 ) );
  OAI212 \u_outFIFO/U306  ( .A(n1423), .B(n950), .C(\u_outFIFO/FIFO[22][3] ), 
        .Q(\u_outFIFO/n422 ) );
  OAI212 \u_outFIFO/U305  ( .A(n1423), .B(n944), .C(\u_outFIFO/n422 ), .Q(
        \u_outFIFO/n642 ) );
  OAI212 \u_outFIFO/U304  ( .A(n804), .B(\u_outFIFO/n372 ), .C(n826), .Q(
        \u_outFIFO/n421 ) );
  OAI212 \u_outFIFO/U303  ( .A(n1422), .B(n950), .C(\u_outFIFO/FIFO[22][2] ), 
        .Q(\u_outFIFO/n420 ) );
  OAI212 \u_outFIFO/U302  ( .A(n1422), .B(n944), .C(\u_outFIFO/n420 ), .Q(
        \u_outFIFO/n641 ) );
  OAI212 \u_outFIFO/U301  ( .A(n804), .B(\u_outFIFO/n369 ), .C(n826), .Q(
        \u_outFIFO/n419 ) );
  OAI212 \u_outFIFO/U300  ( .A(n1421), .B(n950), .C(\u_outFIFO/FIFO[22][1] ), 
        .Q(\u_outFIFO/n418 ) );
  OAI212 \u_outFIFO/U299  ( .A(n1421), .B(n944), .C(\u_outFIFO/n418 ), .Q(
        \u_outFIFO/n640 ) );
  OAI212 \u_outFIFO/U298  ( .A(n804), .B(\u_outFIFO/n366 ), .C(n826), .Q(
        \u_outFIFO/n417 ) );
  OAI212 \u_outFIFO/U297  ( .A(n1420), .B(n951), .C(\u_outFIFO/FIFO[22][0] ), 
        .Q(\u_outFIFO/n416 ) );
  OAI212 \u_outFIFO/U296  ( .A(n1420), .B(n946), .C(\u_outFIFO/n416 ), .Q(
        \u_outFIFO/n639 ) );
  OAI212 \u_outFIFO/U295  ( .A(n802), .B(\u_outFIFO/n375 ), .C(n825), .Q(
        \u_outFIFO/n415 ) );
  OAI212 \u_outFIFO/U294  ( .A(n1419), .B(n951), .C(\u_outFIFO/FIFO[21][3] ), 
        .Q(\u_outFIFO/n414 ) );
  OAI212 \u_outFIFO/U293  ( .A(n1419), .B(n945), .C(\u_outFIFO/n414 ), .Q(
        \u_outFIFO/n638 ) );
  OAI212 \u_outFIFO/U292  ( .A(n802), .B(\u_outFIFO/n372 ), .C(n825), .Q(
        \u_outFIFO/n413 ) );
  OAI212 \u_outFIFO/U291  ( .A(n1418), .B(n951), .C(\u_outFIFO/FIFO[21][2] ), 
        .Q(\u_outFIFO/n412 ) );
  OAI212 \u_outFIFO/U290  ( .A(n1418), .B(n945), .C(\u_outFIFO/n412 ), .Q(
        \u_outFIFO/n637 ) );
  OAI212 \u_outFIFO/U289  ( .A(n802), .B(\u_outFIFO/n369 ), .C(n825), .Q(
        \u_outFIFO/n411 ) );
  OAI212 \u_outFIFO/U288  ( .A(n1417), .B(n951), .C(\u_outFIFO/FIFO[21][1] ), 
        .Q(\u_outFIFO/n410 ) );
  OAI212 \u_outFIFO/U287  ( .A(n1417), .B(n944), .C(\u_outFIFO/n410 ), .Q(
        \u_outFIFO/n636 ) );
  OAI212 \u_outFIFO/U286  ( .A(n802), .B(\u_outFIFO/n366 ), .C(n825), .Q(
        \u_outFIFO/n409 ) );
  OAI212 \u_outFIFO/U285  ( .A(n1416), .B(n951), .C(\u_outFIFO/FIFO[21][0] ), 
        .Q(\u_outFIFO/n408 ) );
  OAI212 \u_outFIFO/U284  ( .A(n1416), .B(n944), .C(\u_outFIFO/n408 ), .Q(
        \u_outFIFO/n635 ) );
  OAI212 \u_outFIFO/U283  ( .A(n800), .B(\u_outFIFO/n375 ), .C(n825), .Q(
        \u_outFIFO/n407 ) );
  OAI212 \u_outFIFO/U282  ( .A(n1415), .B(n951), .C(\u_outFIFO/FIFO[20][3] ), 
        .Q(\u_outFIFO/n406 ) );
  OAI212 \u_outFIFO/U281  ( .A(n1415), .B(n946), .C(\u_outFIFO/n406 ), .Q(
        \u_outFIFO/n634 ) );
  OAI212 \u_outFIFO/U280  ( .A(n800), .B(\u_outFIFO/n372 ), .C(n825), .Q(
        \u_outFIFO/n405 ) );
  OAI212 \u_outFIFO/U279  ( .A(n1414), .B(n951), .C(\u_outFIFO/FIFO[20][2] ), 
        .Q(\u_outFIFO/n404 ) );
  OAI212 \u_outFIFO/U278  ( .A(n1414), .B(n945), .C(\u_outFIFO/n404 ), .Q(
        \u_outFIFO/n633 ) );
  OAI212 \u_outFIFO/U277  ( .A(n800), .B(\u_outFIFO/n369 ), .C(n825), .Q(
        \u_outFIFO/n403 ) );
  OAI212 \u_outFIFO/U276  ( .A(n1413), .B(n951), .C(\u_outFIFO/FIFO[20][1] ), 
        .Q(\u_outFIFO/n402 ) );
  OAI212 \u_outFIFO/U275  ( .A(n1413), .B(n944), .C(\u_outFIFO/n402 ), .Q(
        \u_outFIFO/n632 ) );
  OAI212 \u_outFIFO/U274  ( .A(n800), .B(\u_outFIFO/n366 ), .C(n825), .Q(
        \u_outFIFO/n401 ) );
  OAI212 \u_outFIFO/U273  ( .A(n1412), .B(n951), .C(\u_outFIFO/FIFO[20][0] ), 
        .Q(\u_outFIFO/n400 ) );
  OAI212 \u_outFIFO/U272  ( .A(n1412), .B(n944), .C(\u_outFIFO/n400 ), .Q(
        \u_outFIFO/n631 ) );
  OAI212 \u_outFIFO/U271  ( .A(n798), .B(\u_outFIFO/n375 ), .C(n824), .Q(
        \u_outFIFO/n399 ) );
  OAI212 \u_outFIFO/U270  ( .A(n1411), .B(n951), .C(\u_outFIFO/FIFO[19][3] ), 
        .Q(\u_outFIFO/n398 ) );
  OAI212 \u_outFIFO/U269  ( .A(n1411), .B(n945), .C(\u_outFIFO/n398 ), .Q(
        \u_outFIFO/n630 ) );
  OAI212 \u_outFIFO/U268  ( .A(n798), .B(\u_outFIFO/n372 ), .C(n824), .Q(
        \u_outFIFO/n397 ) );
  OAI212 \u_outFIFO/U267  ( .A(n1410), .B(n951), .C(\u_outFIFO/FIFO[19][2] ), 
        .Q(\u_outFIFO/n396 ) );
  OAI212 \u_outFIFO/U266  ( .A(n1410), .B(n946), .C(\u_outFIFO/n396 ), .Q(
        \u_outFIFO/n629 ) );
  OAI212 \u_outFIFO/U265  ( .A(n798), .B(\u_outFIFO/n369 ), .C(n824), .Q(
        \u_outFIFO/n395 ) );
  OAI212 \u_outFIFO/U264  ( .A(n1409), .B(n951), .C(\u_outFIFO/FIFO[19][1] ), 
        .Q(\u_outFIFO/n394 ) );
  OAI212 \u_outFIFO/U263  ( .A(n1409), .B(n945), .C(\u_outFIFO/n394 ), .Q(
        \u_outFIFO/n628 ) );
  OAI212 \u_outFIFO/U262  ( .A(n798), .B(\u_outFIFO/n366 ), .C(n824), .Q(
        \u_outFIFO/n393 ) );
  OAI212 \u_outFIFO/U261  ( .A(n1408), .B(n951), .C(\u_outFIFO/FIFO[19][0] ), 
        .Q(\u_outFIFO/n392 ) );
  OAI212 \u_outFIFO/U260  ( .A(n1408), .B(n946), .C(\u_outFIFO/n392 ), .Q(
        \u_outFIFO/n627 ) );
  OAI212 \u_outFIFO/U259  ( .A(n796), .B(\u_outFIFO/n375 ), .C(n824), .Q(
        \u_outFIFO/n391 ) );
  OAI212 \u_outFIFO/U258  ( .A(n1407), .B(n952), .C(\u_outFIFO/FIFO[18][3] ), 
        .Q(\u_outFIFO/n390 ) );
  OAI212 \u_outFIFO/U257  ( .A(n1407), .B(n944), .C(\u_outFIFO/n390 ), .Q(
        \u_outFIFO/n626 ) );
  OAI212 \u_outFIFO/U256  ( .A(n796), .B(\u_outFIFO/n372 ), .C(n824), .Q(
        \u_outFIFO/n389 ) );
  OAI212 \u_outFIFO/U255  ( .A(n1406), .B(n952), .C(\u_outFIFO/FIFO[18][2] ), 
        .Q(\u_outFIFO/n388 ) );
  OAI212 \u_outFIFO/U254  ( .A(n1406), .B(n946), .C(\u_outFIFO/n388 ), .Q(
        \u_outFIFO/n625 ) );
  OAI212 \u_outFIFO/U253  ( .A(n796), .B(\u_outFIFO/n369 ), .C(n824), .Q(
        \u_outFIFO/n387 ) );
  OAI212 \u_outFIFO/U252  ( .A(n1405), .B(n952), .C(\u_outFIFO/FIFO[18][1] ), 
        .Q(\u_outFIFO/n386 ) );
  OAI212 \u_outFIFO/U251  ( .A(n1405), .B(n946), .C(\u_outFIFO/n386 ), .Q(
        \u_outFIFO/n624 ) );
  OAI212 \u_outFIFO/U250  ( .A(n796), .B(\u_outFIFO/n366 ), .C(n824), .Q(
        \u_outFIFO/n385 ) );
  OAI212 \u_outFIFO/U249  ( .A(n1404), .B(n952), .C(\u_outFIFO/FIFO[18][0] ), 
        .Q(\u_outFIFO/n384 ) );
  OAI212 \u_outFIFO/U248  ( .A(n1404), .B(n946), .C(\u_outFIFO/n384 ), .Q(
        \u_outFIFO/n623 ) );
  OAI212 \u_outFIFO/U247  ( .A(n794), .B(\u_outFIFO/n375 ), .C(n823), .Q(
        \u_outFIFO/n383 ) );
  OAI212 \u_outFIFO/U246  ( .A(n1403), .B(n952), .C(\u_outFIFO/FIFO[17][3] ), 
        .Q(\u_outFIFO/n382 ) );
  OAI212 \u_outFIFO/U245  ( .A(n1403), .B(n945), .C(\u_outFIFO/n382 ), .Q(
        \u_outFIFO/n622 ) );
  OAI212 \u_outFIFO/U244  ( .A(n794), .B(\u_outFIFO/n372 ), .C(n823), .Q(
        \u_outFIFO/n381 ) );
  OAI212 \u_outFIFO/U243  ( .A(n1402), .B(n952), .C(\u_outFIFO/FIFO[17][2] ), 
        .Q(\u_outFIFO/n380 ) );
  OAI212 \u_outFIFO/U242  ( .A(n1402), .B(n946), .C(\u_outFIFO/n380 ), .Q(
        \u_outFIFO/n621 ) );
  OAI212 \u_outFIFO/U241  ( .A(n794), .B(\u_outFIFO/n369 ), .C(n823), .Q(
        \u_outFIFO/n379 ) );
  OAI212 \u_outFIFO/U240  ( .A(n1401), .B(n952), .C(\u_outFIFO/FIFO[17][1] ), 
        .Q(\u_outFIFO/n378 ) );
  OAI212 \u_outFIFO/U239  ( .A(n1401), .B(n944), .C(\u_outFIFO/n378 ), .Q(
        \u_outFIFO/n620 ) );
  OAI212 \u_outFIFO/U238  ( .A(n794), .B(\u_outFIFO/n366 ), .C(n823), .Q(
        \u_outFIFO/n377 ) );
  OAI212 \u_outFIFO/U237  ( .A(n1400), .B(n952), .C(\u_outFIFO/FIFO[17][0] ), 
        .Q(\u_outFIFO/n376 ) );
  OAI212 \u_outFIFO/U236  ( .A(n1400), .B(n945), .C(\u_outFIFO/n376 ), .Q(
        \u_outFIFO/n619 ) );
  OAI212 \u_outFIFO/U235  ( .A(n791), .B(\u_outFIFO/n375 ), .C(n823), .Q(
        \u_outFIFO/n374 ) );
  OAI212 \u_outFIFO/U234  ( .A(n1399), .B(n952), .C(\u_outFIFO/FIFO[16][3] ), 
        .Q(\u_outFIFO/n373 ) );
  OAI212 \u_outFIFO/U233  ( .A(n1399), .B(n945), .C(\u_outFIFO/n373 ), .Q(
        \u_outFIFO/n618 ) );
  OAI212 \u_outFIFO/U232  ( .A(n791), .B(\u_outFIFO/n372 ), .C(n823), .Q(
        \u_outFIFO/n371 ) );
  OAI212 \u_outFIFO/U231  ( .A(n1398), .B(n952), .C(\u_outFIFO/FIFO[16][2] ), 
        .Q(\u_outFIFO/n370 ) );
  OAI212 \u_outFIFO/U230  ( .A(n1398), .B(n946), .C(\u_outFIFO/n370 ), .Q(
        \u_outFIFO/n617 ) );
  OAI212 \u_outFIFO/U229  ( .A(n791), .B(\u_outFIFO/n369 ), .C(n823), .Q(
        \u_outFIFO/n368 ) );
  OAI212 \u_outFIFO/U228  ( .A(n1397), .B(n952), .C(\u_outFIFO/FIFO[16][1] ), 
        .Q(\u_outFIFO/n367 ) );
  OAI212 \u_outFIFO/U227  ( .A(n1397), .B(n945), .C(\u_outFIFO/n367 ), .Q(
        \u_outFIFO/n616 ) );
  OAI212 \u_outFIFO/U226  ( .A(n791), .B(\u_outFIFO/n366 ), .C(n823), .Q(
        \u_outFIFO/n365 ) );
  OAI212 \u_outFIFO/U225  ( .A(n1396), .B(n952), .C(\u_outFIFO/FIFO[16][0] ), 
        .Q(\u_outFIFO/n364 ) );
  OAI212 \u_outFIFO/U224  ( .A(n1396), .B(n945), .C(\u_outFIFO/n364 ), .Q(
        \u_outFIFO/n615 ) );
  OAI212 \u_outFIFO/U221  ( .A(n807), .B(\u_outFIFO/n306 ), .C(n822), .Q(
        \u_outFIFO/n363 ) );
  OAI212 \u_outFIFO/U220  ( .A(n1395), .B(n952), .C(\u_outFIFO/FIFO[15][3] ), 
        .Q(\u_outFIFO/n362 ) );
  OAI212 \u_outFIFO/U219  ( .A(n1395), .B(n944), .C(\u_outFIFO/n362 ), .Q(
        \u_outFIFO/n614 ) );
  OAI212 \u_outFIFO/U217  ( .A(n807), .B(\u_outFIFO/n303 ), .C(n822), .Q(
        \u_outFIFO/n361 ) );
  OAI212 \u_outFIFO/U216  ( .A(n1394), .B(\u_outFIFO/n215 ), .C(
        \u_outFIFO/FIFO[15][2] ), .Q(\u_outFIFO/n360 ) );
  OAI212 \u_outFIFO/U215  ( .A(n1394), .B(\u_outFIFO/n213 ), .C(
        \u_outFIFO/n360 ), .Q(\u_outFIFO/n613 ) );
  OAI212 \u_outFIFO/U213  ( .A(n807), .B(\u_outFIFO/n300 ), .C(n822), .Q(
        \u_outFIFO/n359 ) );
  OAI212 \u_outFIFO/U212  ( .A(n1393), .B(\u_outFIFO/n215 ), .C(
        \u_outFIFO/FIFO[15][1] ), .Q(\u_outFIFO/n358 ) );
  OAI212 \u_outFIFO/U211  ( .A(n1393), .B(\u_outFIFO/n213 ), .C(
        \u_outFIFO/n358 ), .Q(\u_outFIFO/n612 ) );
  OAI212 \u_outFIFO/U209  ( .A(n807), .B(\u_outFIFO/n297 ), .C(n822), .Q(
        \u_outFIFO/n356 ) );
  OAI212 \u_outFIFO/U208  ( .A(n1392), .B(n950), .C(\u_outFIFO/FIFO[15][0] ), 
        .Q(\u_outFIFO/n355 ) );
  OAI212 \u_outFIFO/U207  ( .A(n1392), .B(\u_outFIFO/n213 ), .C(
        \u_outFIFO/n355 ), .Q(\u_outFIFO/n611 ) );
  OAI212 \u_outFIFO/U206  ( .A(n804), .B(\u_outFIFO/n306 ), .C(n822), .Q(
        \u_outFIFO/n354 ) );
  OAI212 \u_outFIFO/U205  ( .A(n1391), .B(n949), .C(\u_outFIFO/FIFO[14][3] ), 
        .Q(\u_outFIFO/n353 ) );
  OAI212 \u_outFIFO/U204  ( .A(n1391), .B(\u_outFIFO/n213 ), .C(
        \u_outFIFO/n353 ), .Q(\u_outFIFO/n610 ) );
  OAI212 \u_outFIFO/U203  ( .A(n804), .B(\u_outFIFO/n303 ), .C(n822), .Q(
        \u_outFIFO/n352 ) );
  OAI212 \u_outFIFO/U202  ( .A(n1390), .B(n948), .C(\u_outFIFO/FIFO[14][2] ), 
        .Q(\u_outFIFO/n351 ) );
  OAI212 \u_outFIFO/U201  ( .A(n1390), .B(n805), .C(\u_outFIFO/n351 ), .Q(
        \u_outFIFO/n609 ) );
  OAI212 \u_outFIFO/U200  ( .A(n804), .B(\u_outFIFO/n300 ), .C(n822), .Q(
        \u_outFIFO/n350 ) );
  OAI212 \u_outFIFO/U199  ( .A(n1389), .B(n950), .C(\u_outFIFO/FIFO[14][1] ), 
        .Q(\u_outFIFO/n349 ) );
  OAI212 \u_outFIFO/U198  ( .A(n1389), .B(n947), .C(\u_outFIFO/n349 ), .Q(
        \u_outFIFO/n608 ) );
  OAI212 \u_outFIFO/U197  ( .A(n804), .B(\u_outFIFO/n297 ), .C(n822), .Q(
        \u_outFIFO/n348 ) );
  OAI212 \u_outFIFO/U196  ( .A(n1388), .B(n949), .C(\u_outFIFO/FIFO[14][0] ), 
        .Q(\u_outFIFO/n347 ) );
  OAI212 \u_outFIFO/U195  ( .A(n1388), .B(n944), .C(\u_outFIFO/n347 ), .Q(
        \u_outFIFO/n607 ) );
  OAI212 \u_outFIFO/U194  ( .A(n802), .B(\u_outFIFO/n306 ), .C(n821), .Q(
        \u_outFIFO/n346 ) );
  OAI212 \u_outFIFO/U193  ( .A(n1387), .B(n948), .C(\u_outFIFO/FIFO[13][3] ), 
        .Q(\u_outFIFO/n345 ) );
  OAI212 \u_outFIFO/U192  ( .A(n1387), .B(n946), .C(\u_outFIFO/n345 ), .Q(
        \u_outFIFO/n606 ) );
  OAI212 \u_outFIFO/U191  ( .A(n802), .B(\u_outFIFO/n303 ), .C(n821), .Q(
        \u_outFIFO/n344 ) );
  OAI212 \u_outFIFO/U190  ( .A(n1386), .B(n950), .C(\u_outFIFO/FIFO[13][2] ), 
        .Q(\u_outFIFO/n343 ) );
  OAI212 \u_outFIFO/U189  ( .A(n1386), .B(n945), .C(\u_outFIFO/n343 ), .Q(
        \u_outFIFO/n605 ) );
  OAI212 \u_outFIFO/U188  ( .A(n802), .B(\u_outFIFO/n300 ), .C(n821), .Q(
        \u_outFIFO/n342 ) );
  OAI212 \u_outFIFO/U187  ( .A(n1385), .B(n949), .C(\u_outFIFO/FIFO[13][1] ), 
        .Q(\u_outFIFO/n341 ) );
  OAI212 \u_outFIFO/U186  ( .A(n1385), .B(n944), .C(\u_outFIFO/n341 ), .Q(
        \u_outFIFO/n604 ) );
  OAI212 \u_outFIFO/U185  ( .A(n802), .B(\u_outFIFO/n297 ), .C(n821), .Q(
        \u_outFIFO/n340 ) );
  OAI212 \u_outFIFO/U184  ( .A(n1384), .B(n948), .C(\u_outFIFO/FIFO[13][0] ), 
        .Q(\u_outFIFO/n339 ) );
  OAI212 \u_outFIFO/U183  ( .A(n1384), .B(n946), .C(\u_outFIFO/n339 ), .Q(
        \u_outFIFO/n603 ) );
  OAI212 \u_outFIFO/U182  ( .A(n800), .B(\u_outFIFO/n306 ), .C(n821), .Q(
        \u_outFIFO/n338 ) );
  OAI212 \u_outFIFO/U181  ( .A(n1383), .B(n952), .C(\u_outFIFO/FIFO[12][3] ), 
        .Q(\u_outFIFO/n337 ) );
  OAI212 \u_outFIFO/U180  ( .A(n1383), .B(n945), .C(\u_outFIFO/n337 ), .Q(
        \u_outFIFO/n602 ) );
  OAI212 \u_outFIFO/U179  ( .A(n800), .B(\u_outFIFO/n303 ), .C(n821), .Q(
        \u_outFIFO/n336 ) );
  OAI212 \u_outFIFO/U178  ( .A(n1382), .B(n951), .C(\u_outFIFO/FIFO[12][2] ), 
        .Q(\u_outFIFO/n335 ) );
  OAI212 \u_outFIFO/U177  ( .A(n1382), .B(n944), .C(\u_outFIFO/n335 ), .Q(
        \u_outFIFO/n601 ) );
  OAI212 \u_outFIFO/U176  ( .A(n800), .B(\u_outFIFO/n300 ), .C(n821), .Q(
        \u_outFIFO/n334 ) );
  OAI212 \u_outFIFO/U175  ( .A(n1381), .B(n953), .C(\u_outFIFO/FIFO[12][1] ), 
        .Q(\u_outFIFO/n333 ) );
  OAI212 \u_outFIFO/U174  ( .A(n1381), .B(n946), .C(\u_outFIFO/n333 ), .Q(
        \u_outFIFO/n600 ) );
  OAI212 \u_outFIFO/U173  ( .A(n800), .B(\u_outFIFO/n297 ), .C(n821), .Q(
        \u_outFIFO/n332 ) );
  OAI212 \u_outFIFO/U172  ( .A(n1380), .B(n953), .C(\u_outFIFO/FIFO[12][0] ), 
        .Q(\u_outFIFO/n331 ) );
  OAI212 \u_outFIFO/U171  ( .A(n1380), .B(n944), .C(\u_outFIFO/n331 ), .Q(
        \u_outFIFO/n599 ) );
  OAI212 \u_outFIFO/U170  ( .A(n798), .B(\u_outFIFO/n306 ), .C(n820), .Q(
        \u_outFIFO/n330 ) );
  OAI212 \u_outFIFO/U169  ( .A(n1379), .B(n953), .C(\u_outFIFO/FIFO[11][3] ), 
        .Q(\u_outFIFO/n329 ) );
  OAI212 \u_outFIFO/U168  ( .A(n1379), .B(n945), .C(\u_outFIFO/n329 ), .Q(
        \u_outFIFO/n598 ) );
  OAI212 \u_outFIFO/U167  ( .A(n798), .B(\u_outFIFO/n303 ), .C(n820), .Q(
        \u_outFIFO/n328 ) );
  OAI212 \u_outFIFO/U166  ( .A(n1378), .B(n953), .C(\u_outFIFO/FIFO[11][2] ), 
        .Q(\u_outFIFO/n327 ) );
  OAI212 \u_outFIFO/U165  ( .A(n1378), .B(n946), .C(\u_outFIFO/n327 ), .Q(
        \u_outFIFO/n597 ) );
  OAI212 \u_outFIFO/U164  ( .A(n798), .B(\u_outFIFO/n300 ), .C(n820), .Q(
        \u_outFIFO/n326 ) );
  OAI212 \u_outFIFO/U163  ( .A(n1377), .B(n953), .C(\u_outFIFO/FIFO[11][1] ), 
        .Q(\u_outFIFO/n325 ) );
  OAI212 \u_outFIFO/U162  ( .A(n1377), .B(n945), .C(\u_outFIFO/n325 ), .Q(
        \u_outFIFO/n596 ) );
  OAI212 \u_outFIFO/U161  ( .A(n798), .B(\u_outFIFO/n297 ), .C(n820), .Q(
        \u_outFIFO/n324 ) );
  OAI212 \u_outFIFO/U160  ( .A(n1376), .B(n953), .C(\u_outFIFO/FIFO[11][0] ), 
        .Q(\u_outFIFO/n323 ) );
  OAI212 \u_outFIFO/U159  ( .A(n1376), .B(n944), .C(\u_outFIFO/n323 ), .Q(
        \u_outFIFO/n595 ) );
  OAI212 \u_outFIFO/U158  ( .A(n796), .B(\u_outFIFO/n306 ), .C(n820), .Q(
        \u_outFIFO/n322 ) );
  OAI212 \u_outFIFO/U157  ( .A(n1375), .B(n953), .C(\u_outFIFO/FIFO[10][3] ), 
        .Q(\u_outFIFO/n321 ) );
  OAI212 \u_outFIFO/U156  ( .A(n1375), .B(n946), .C(\u_outFIFO/n321 ), .Q(
        \u_outFIFO/n594 ) );
  OAI212 \u_outFIFO/U155  ( .A(n796), .B(\u_outFIFO/n303 ), .C(n820), .Q(
        \u_outFIFO/n320 ) );
  OAI212 \u_outFIFO/U154  ( .A(n1374), .B(n953), .C(\u_outFIFO/FIFO[10][2] ), 
        .Q(\u_outFIFO/n319 ) );
  OAI212 \u_outFIFO/U153  ( .A(n1374), .B(n945), .C(\u_outFIFO/n319 ), .Q(
        \u_outFIFO/n593 ) );
  OAI212 \u_outFIFO/U152  ( .A(n796), .B(\u_outFIFO/n300 ), .C(n820), .Q(
        \u_outFIFO/n318 ) );
  OAI212 \u_outFIFO/U151  ( .A(n1373), .B(n953), .C(\u_outFIFO/FIFO[10][1] ), 
        .Q(\u_outFIFO/n317 ) );
  OAI212 \u_outFIFO/U150  ( .A(n1373), .B(n944), .C(\u_outFIFO/n317 ), .Q(
        \u_outFIFO/n592 ) );
  OAI212 \u_outFIFO/U149  ( .A(n796), .B(\u_outFIFO/n297 ), .C(n820), .Q(
        \u_outFIFO/n316 ) );
  OAI212 \u_outFIFO/U148  ( .A(n1372), .B(n953), .C(\u_outFIFO/FIFO[10][0] ), 
        .Q(\u_outFIFO/n315 ) );
  OAI212 \u_outFIFO/U147  ( .A(n1372), .B(n944), .C(\u_outFIFO/n315 ), .Q(
        \u_outFIFO/n591 ) );
  OAI212 \u_outFIFO/U146  ( .A(n794), .B(\u_outFIFO/n306 ), .C(n819), .Q(
        \u_outFIFO/n314 ) );
  OAI212 \u_outFIFO/U145  ( .A(n1371), .B(n953), .C(\u_outFIFO/FIFO[9][3] ), 
        .Q(\u_outFIFO/n313 ) );
  OAI212 \u_outFIFO/U144  ( .A(n1371), .B(n946), .C(\u_outFIFO/n313 ), .Q(
        \u_outFIFO/n590 ) );
  OAI212 \u_outFIFO/U143  ( .A(n794), .B(\u_outFIFO/n303 ), .C(n819), .Q(
        \u_outFIFO/n312 ) );
  OAI212 \u_outFIFO/U142  ( .A(n1370), .B(n953), .C(\u_outFIFO/FIFO[9][2] ), 
        .Q(\u_outFIFO/n311 ) );
  OAI212 \u_outFIFO/U141  ( .A(n1370), .B(n945), .C(\u_outFIFO/n311 ), .Q(
        \u_outFIFO/n589 ) );
  OAI212 \u_outFIFO/U140  ( .A(n794), .B(\u_outFIFO/n300 ), .C(n819), .Q(
        \u_outFIFO/n310 ) );
  OAI212 \u_outFIFO/U139  ( .A(n1369), .B(n953), .C(\u_outFIFO/FIFO[9][1] ), 
        .Q(\u_outFIFO/n309 ) );
  OAI212 \u_outFIFO/U138  ( .A(n1369), .B(n946), .C(\u_outFIFO/n309 ), .Q(
        \u_outFIFO/n588 ) );
  OAI212 \u_outFIFO/U137  ( .A(n794), .B(\u_outFIFO/n297 ), .C(n819), .Q(
        \u_outFIFO/n308 ) );
  OAI212 \u_outFIFO/U136  ( .A(n1368), .B(n950), .C(\u_outFIFO/FIFO[9][0] ), 
        .Q(\u_outFIFO/n307 ) );
  OAI212 \u_outFIFO/U135  ( .A(n1368), .B(n945), .C(\u_outFIFO/n307 ), .Q(
        \u_outFIFO/n587 ) );
  OAI212 \u_outFIFO/U134  ( .A(n792), .B(\u_outFIFO/n306 ), .C(n819), .Q(
        \u_outFIFO/n305 ) );
  OAI212 \u_outFIFO/U133  ( .A(n1367), .B(n949), .C(\u_outFIFO/FIFO[8][3] ), 
        .Q(\u_outFIFO/n304 ) );
  OAI212 \u_outFIFO/U132  ( .A(n1367), .B(n945), .C(\u_outFIFO/n304 ), .Q(
        \u_outFIFO/n586 ) );
  OAI212 \u_outFIFO/U131  ( .A(n792), .B(\u_outFIFO/n303 ), .C(n819), .Q(
        \u_outFIFO/n302 ) );
  OAI212 \u_outFIFO/U130  ( .A(n1366), .B(n948), .C(\u_outFIFO/FIFO[8][2] ), 
        .Q(\u_outFIFO/n301 ) );
  OAI212 \u_outFIFO/U129  ( .A(n1366), .B(n945), .C(\u_outFIFO/n301 ), .Q(
        \u_outFIFO/n585 ) );
  OAI212 \u_outFIFO/U128  ( .A(n792), .B(\u_outFIFO/n300 ), .C(n819), .Q(
        \u_outFIFO/n299 ) );
  OAI212 \u_outFIFO/U127  ( .A(n1365), .B(n952), .C(\u_outFIFO/FIFO[8][1] ), 
        .Q(\u_outFIFO/n298 ) );
  OAI212 \u_outFIFO/U126  ( .A(n1365), .B(n945), .C(\u_outFIFO/n298 ), .Q(
        \u_outFIFO/n584 ) );
  OAI212 \u_outFIFO/U125  ( .A(n792), .B(\u_outFIFO/n297 ), .C(n819), .Q(
        \u_outFIFO/n296 ) );
  OAI212 \u_outFIFO/U124  ( .A(n1364), .B(n951), .C(\u_outFIFO/FIFO[8][0] ), 
        .Q(\u_outFIFO/n295 ) );
  OAI212 \u_outFIFO/U123  ( .A(n1364), .B(n945), .C(\u_outFIFO/n295 ), .Q(
        \u_outFIFO/n583 ) );
  OAI212 \u_outFIFO/U120  ( .A(\u_outFIFO/n227 ), .B(n806), .C(n818), .Q(
        \u_outFIFO/n293 ) );
  OAI212 \u_outFIFO/U119  ( .A(n1363), .B(n952), .C(\u_outFIFO/FIFO[7][3] ), 
        .Q(\u_outFIFO/n292 ) );
  OAI212 \u_outFIFO/U118  ( .A(n1363), .B(n945), .C(\u_outFIFO/n292 ), .Q(
        \u_outFIFO/n582 ) );
  OAI212 \u_outFIFO/U116  ( .A(\u_outFIFO/n224 ), .B(n806), .C(n818), .Q(
        \u_outFIFO/n290 ) );
  OAI212 \u_outFIFO/U115  ( .A(n1362), .B(n951), .C(\u_outFIFO/FIFO[7][2] ), 
        .Q(\u_outFIFO/n289 ) );
  OAI212 \u_outFIFO/U114  ( .A(n1362), .B(n945), .C(\u_outFIFO/n289 ), .Q(
        \u_outFIFO/n581 ) );
  OAI212 \u_outFIFO/U112  ( .A(\u_outFIFO/n221 ), .B(n806), .C(n818), .Q(
        \u_outFIFO/n287 ) );
  OAI212 \u_outFIFO/U111  ( .A(n1361), .B(n952), .C(\u_outFIFO/FIFO[7][1] ), 
        .Q(\u_outFIFO/n286 ) );
  OAI212 \u_outFIFO/U110  ( .A(n1361), .B(n945), .C(\u_outFIFO/n286 ), .Q(
        \u_outFIFO/n580 ) );
  OAI212 \u_outFIFO/U108  ( .A(\u_outFIFO/n218 ), .B(n806), .C(n818), .Q(
        \u_outFIFO/n283 ) );
  OAI212 \u_outFIFO/U107  ( .A(n1360), .B(n951), .C(\u_outFIFO/FIFO[7][0] ), 
        .Q(\u_outFIFO/n282 ) );
  OAI212 \u_outFIFO/U106  ( .A(n1360), .B(n945), .C(\u_outFIFO/n282 ), .Q(
        \u_outFIFO/n579 ) );
  OAI212 \u_outFIFO/U105  ( .A(\u_outFIFO/n227 ), .B(n803), .C(n818), .Q(
        \u_outFIFO/n281 ) );
  OAI212 \u_outFIFO/U104  ( .A(n1359), .B(n954), .C(\u_outFIFO/FIFO[6][3] ), 
        .Q(\u_outFIFO/n280 ) );
  OAI212 \u_outFIFO/U103  ( .A(n1359), .B(n945), .C(\u_outFIFO/n280 ), .Q(
        \u_outFIFO/n578 ) );
  OAI212 \u_outFIFO/U102  ( .A(\u_outFIFO/n224 ), .B(n803), .C(n818), .Q(
        \u_outFIFO/n279 ) );
  OAI212 \u_outFIFO/U101  ( .A(n1358), .B(n953), .C(\u_outFIFO/FIFO[6][2] ), 
        .Q(\u_outFIFO/n278 ) );
  OAI212 \u_outFIFO/U100  ( .A(n1358), .B(n945), .C(\u_outFIFO/n278 ), .Q(
        \u_outFIFO/n577 ) );
  OAI212 \u_outFIFO/U99  ( .A(\u_outFIFO/n221 ), .B(n803), .C(n818), .Q(
        \u_outFIFO/n277 ) );
  OAI212 \u_outFIFO/U98  ( .A(n1357), .B(n952), .C(\u_outFIFO/FIFO[6][1] ), 
        .Q(\u_outFIFO/n276 ) );
  OAI212 \u_outFIFO/U97  ( .A(n1357), .B(n945), .C(\u_outFIFO/n276 ), .Q(
        \u_outFIFO/n576 ) );
  OAI212 \u_outFIFO/U96  ( .A(\u_outFIFO/n218 ), .B(n803), .C(n818), .Q(
        \u_outFIFO/n274 ) );
  OAI212 \u_outFIFO/U95  ( .A(n1356), .B(n954), .C(\u_outFIFO/FIFO[6][0] ), 
        .Q(\u_outFIFO/n273 ) );
  OAI212 \u_outFIFO/U94  ( .A(n1356), .B(n945), .C(\u_outFIFO/n273 ), .Q(
        \u_outFIFO/n575 ) );
  OAI212 \u_outFIFO/U93  ( .A(\u_outFIFO/n227 ), .B(n801), .C(n817), .Q(
        \u_outFIFO/n272 ) );
  OAI212 \u_outFIFO/U92  ( .A(n1355), .B(n954), .C(\u_outFIFO/FIFO[5][3] ), 
        .Q(\u_outFIFO/n271 ) );
  OAI212 \u_outFIFO/U91  ( .A(n1355), .B(n946), .C(\u_outFIFO/n271 ), .Q(
        \u_outFIFO/n574 ) );
  OAI212 \u_outFIFO/U90  ( .A(\u_outFIFO/n224 ), .B(n801), .C(n817), .Q(
        \u_outFIFO/n270 ) );
  OAI212 \u_outFIFO/U89  ( .A(n1354), .B(n954), .C(\u_outFIFO/FIFO[5][2] ), 
        .Q(\u_outFIFO/n269 ) );
  OAI212 \u_outFIFO/U88  ( .A(n1354), .B(n946), .C(\u_outFIFO/n269 ), .Q(
        \u_outFIFO/n573 ) );
  OAI212 \u_outFIFO/U87  ( .A(\u_outFIFO/n221 ), .B(n801), .C(n817), .Q(
        \u_outFIFO/n268 ) );
  OAI212 \u_outFIFO/U86  ( .A(n1353), .B(n954), .C(\u_outFIFO/FIFO[5][1] ), 
        .Q(\u_outFIFO/n267 ) );
  OAI212 \u_outFIFO/U85  ( .A(n1353), .B(n946), .C(\u_outFIFO/n267 ), .Q(
        \u_outFIFO/n572 ) );
  OAI212 \u_outFIFO/U84  ( .A(\u_outFIFO/n218 ), .B(n801), .C(n817), .Q(
        \u_outFIFO/n265 ) );
  OAI212 \u_outFIFO/U83  ( .A(n1352), .B(n954), .C(\u_outFIFO/FIFO[5][0] ), 
        .Q(\u_outFIFO/n264 ) );
  OAI212 \u_outFIFO/U82  ( .A(n1352), .B(n946), .C(\u_outFIFO/n264 ), .Q(
        \u_outFIFO/n571 ) );
  OAI212 \u_outFIFO/U81  ( .A(\u_outFIFO/n227 ), .B(n799), .C(n817), .Q(
        \u_outFIFO/n263 ) );
  OAI212 \u_outFIFO/U80  ( .A(n1351), .B(n954), .C(\u_outFIFO/FIFO[4][3] ), 
        .Q(\u_outFIFO/n262 ) );
  OAI212 \u_outFIFO/U79  ( .A(n1351), .B(n946), .C(\u_outFIFO/n262 ), .Q(
        \u_outFIFO/n570 ) );
  OAI212 \u_outFIFO/U78  ( .A(\u_outFIFO/n224 ), .B(n799), .C(n817), .Q(
        \u_outFIFO/n261 ) );
  OAI212 \u_outFIFO/U77  ( .A(n1350), .B(n954), .C(\u_outFIFO/FIFO[4][2] ), 
        .Q(\u_outFIFO/n260 ) );
  OAI212 \u_outFIFO/U76  ( .A(n1350), .B(n946), .C(\u_outFIFO/n260 ), .Q(
        \u_outFIFO/n569 ) );
  OAI212 \u_outFIFO/U75  ( .A(\u_outFIFO/n221 ), .B(n799), .C(n817), .Q(
        \u_outFIFO/n259 ) );
  OAI212 \u_outFIFO/U74  ( .A(n1349), .B(n954), .C(\u_outFIFO/FIFO[4][1] ), 
        .Q(\u_outFIFO/n258 ) );
  OAI212 \u_outFIFO/U73  ( .A(n1349), .B(n946), .C(\u_outFIFO/n258 ), .Q(
        \u_outFIFO/n568 ) );
  OAI212 \u_outFIFO/U72  ( .A(\u_outFIFO/n218 ), .B(n799), .C(n817), .Q(
        \u_outFIFO/n256 ) );
  OAI212 \u_outFIFO/U71  ( .A(n1348), .B(n954), .C(\u_outFIFO/FIFO[4][0] ), 
        .Q(\u_outFIFO/n255 ) );
  OAI212 \u_outFIFO/U70  ( .A(n1348), .B(n946), .C(\u_outFIFO/n255 ), .Q(
        \u_outFIFO/n567 ) );
  OAI212 \u_outFIFO/U69  ( .A(\u_outFIFO/n227 ), .B(n797), .C(n816), .Q(
        \u_outFIFO/n254 ) );
  OAI212 \u_outFIFO/U68  ( .A(n1347), .B(n954), .C(\u_outFIFO/FIFO[3][3] ), 
        .Q(\u_outFIFO/n253 ) );
  OAI212 \u_outFIFO/U67  ( .A(n1347), .B(n946), .C(\u_outFIFO/n253 ), .Q(
        \u_outFIFO/n566 ) );
  OAI212 \u_outFIFO/U66  ( .A(\u_outFIFO/n224 ), .B(n797), .C(n816), .Q(
        \u_outFIFO/n252 ) );
  OAI212 \u_outFIFO/U65  ( .A(n1346), .B(n954), .C(\u_outFIFO/FIFO[3][2] ), 
        .Q(\u_outFIFO/n251 ) );
  OAI212 \u_outFIFO/U64  ( .A(n1346), .B(n946), .C(\u_outFIFO/n251 ), .Q(
        \u_outFIFO/n565 ) );
  OAI212 \u_outFIFO/U63  ( .A(\u_outFIFO/n221 ), .B(n797), .C(n816), .Q(
        \u_outFIFO/n250 ) );
  OAI212 \u_outFIFO/U62  ( .A(n1345), .B(n954), .C(\u_outFIFO/FIFO[3][1] ), 
        .Q(\u_outFIFO/n249 ) );
  OAI212 \u_outFIFO/U61  ( .A(n1345), .B(n946), .C(\u_outFIFO/n249 ), .Q(
        \u_outFIFO/n564 ) );
  OAI212 \u_outFIFO/U60  ( .A(\u_outFIFO/n218 ), .B(n797), .C(n816), .Q(
        \u_outFIFO/n247 ) );
  OAI212 \u_outFIFO/U59  ( .A(n1344), .B(n954), .C(\u_outFIFO/FIFO[3][0] ), 
        .Q(\u_outFIFO/n246 ) );
  OAI212 \u_outFIFO/U58  ( .A(n1344), .B(n946), .C(\u_outFIFO/n246 ), .Q(
        \u_outFIFO/n563 ) );
  OAI212 \u_outFIFO/U57  ( .A(\u_outFIFO/n227 ), .B(n795), .C(n816), .Q(
        \u_outFIFO/n245 ) );
  OAI212 \u_outFIFO/U56  ( .A(n1343), .B(n954), .C(\u_outFIFO/FIFO[2][3] ), 
        .Q(\u_outFIFO/n244 ) );
  OAI212 \u_outFIFO/U55  ( .A(n1343), .B(n946), .C(\u_outFIFO/n244 ), .Q(
        \u_outFIFO/n562 ) );
  OAI212 \u_outFIFO/U54  ( .A(\u_outFIFO/n224 ), .B(n795), .C(n816), .Q(
        \u_outFIFO/n243 ) );
  OAI212 \u_outFIFO/U53  ( .A(n1342), .B(n953), .C(\u_outFIFO/FIFO[2][2] ), 
        .Q(\u_outFIFO/n242 ) );
  OAI212 \u_outFIFO/U52  ( .A(n1342), .B(n947), .C(\u_outFIFO/n242 ), .Q(
        \u_outFIFO/n561 ) );
  OAI212 \u_outFIFO/U51  ( .A(\u_outFIFO/n221 ), .B(n795), .C(n816), .Q(
        \u_outFIFO/n241 ) );
  OAI212 \u_outFIFO/U50  ( .A(n1341), .B(n950), .C(\u_outFIFO/FIFO[2][1] ), 
        .Q(\u_outFIFO/n240 ) );
  OAI212 \u_outFIFO/U49  ( .A(n1341), .B(n947), .C(\u_outFIFO/n240 ), .Q(
        \u_outFIFO/n560 ) );
  OAI212 \u_outFIFO/U48  ( .A(\u_outFIFO/n218 ), .B(n795), .C(n816), .Q(
        \u_outFIFO/n238 ) );
  OAI212 \u_outFIFO/U47  ( .A(n1340), .B(n954), .C(\u_outFIFO/FIFO[2][0] ), 
        .Q(\u_outFIFO/n237 ) );
  OAI212 \u_outFIFO/U46  ( .A(n1340), .B(n947), .C(\u_outFIFO/n237 ), .Q(
        \u_outFIFO/n559 ) );
  OAI212 \u_outFIFO/U45  ( .A(\u_outFIFO/n227 ), .B(n793), .C(n815), .Q(
        \u_outFIFO/n236 ) );
  OAI212 \u_outFIFO/U44  ( .A(n1339), .B(n953), .C(\u_outFIFO/FIFO[1][3] ), 
        .Q(\u_outFIFO/n235 ) );
  OAI212 \u_outFIFO/U43  ( .A(n1339), .B(n947), .C(\u_outFIFO/n235 ), .Q(
        \u_outFIFO/n558 ) );
  OAI212 \u_outFIFO/U42  ( .A(\u_outFIFO/n224 ), .B(n793), .C(n815), .Q(
        \u_outFIFO/n234 ) );
  OAI212 \u_outFIFO/U41  ( .A(n1338), .B(n953), .C(\u_outFIFO/FIFO[1][2] ), 
        .Q(\u_outFIFO/n233 ) );
  OAI212 \u_outFIFO/U40  ( .A(n1338), .B(n947), .C(\u_outFIFO/n233 ), .Q(
        \u_outFIFO/n557 ) );
  OAI212 \u_outFIFO/U39  ( .A(\u_outFIFO/n221 ), .B(n793), .C(n815), .Q(
        \u_outFIFO/n232 ) );
  OAI212 \u_outFIFO/U38  ( .A(n1337), .B(n949), .C(\u_outFIFO/FIFO[1][1] ), 
        .Q(\u_outFIFO/n231 ) );
  OAI212 \u_outFIFO/U37  ( .A(n1337), .B(n947), .C(\u_outFIFO/n231 ), .Q(
        \u_outFIFO/n556 ) );
  OAI212 \u_outFIFO/U36  ( .A(\u_outFIFO/n218 ), .B(n793), .C(n815), .Q(
        \u_outFIFO/n229 ) );
  OAI212 \u_outFIFO/U35  ( .A(n1336), .B(n954), .C(\u_outFIFO/FIFO[1][0] ), 
        .Q(\u_outFIFO/n228 ) );
  OAI212 \u_outFIFO/U34  ( .A(n1336), .B(n947), .C(\u_outFIFO/n228 ), .Q(
        \u_outFIFO/n555 ) );
  OAI212 \u_outFIFO/U33  ( .A(n792), .B(\u_outFIFO/n227 ), .C(n815), .Q(
        \u_outFIFO/n226 ) );
  OAI212 \u_outFIFO/U32  ( .A(n1335), .B(n951), .C(\u_outFIFO/FIFO[0][3] ), 
        .Q(\u_outFIFO/n225 ) );
  OAI212 \u_outFIFO/U31  ( .A(n1335), .B(n947), .C(\u_outFIFO/n225 ), .Q(
        \u_outFIFO/n554 ) );
  OAI212 \u_outFIFO/U30  ( .A(n792), .B(\u_outFIFO/n224 ), .C(n815), .Q(
        \u_outFIFO/n223 ) );
  OAI212 \u_outFIFO/U29  ( .A(n1334), .B(n953), .C(\u_outFIFO/FIFO[0][2] ), 
        .Q(\u_outFIFO/n222 ) );
  OAI212 \u_outFIFO/U28  ( .A(n1334), .B(n947), .C(\u_outFIFO/n222 ), .Q(
        \u_outFIFO/n553 ) );
  OAI212 \u_outFIFO/U27  ( .A(n792), .B(\u_outFIFO/n221 ), .C(n815), .Q(
        \u_outFIFO/n220 ) );
  OAI212 \u_outFIFO/U26  ( .A(n1333), .B(n948), .C(\u_outFIFO/FIFO[0][1] ), 
        .Q(\u_outFIFO/n219 ) );
  OAI212 \u_outFIFO/U25  ( .A(n1333), .B(n947), .C(\u_outFIFO/n219 ), .Q(
        \u_outFIFO/n552 ) );
  OAI212 \u_outFIFO/U24  ( .A(n792), .B(\u_outFIFO/n218 ), .C(n815), .Q(
        \u_outFIFO/n216 ) );
  OAI212 \u_outFIFO/U23  ( .A(n1332), .B(n954), .C(\u_outFIFO/FIFO[0][0] ), 
        .Q(\u_outFIFO/n214 ) );
  OAI212 \u_outFIFO/U22  ( .A(n1332), .B(n947), .C(\u_outFIFO/n214 ), .Q(
        \u_outFIFO/n551 ) );
  OAI222 \u_mux8/U1  ( .A(\u_mux8/n3 ), .B(n1688), .C(in_MUX_inSEL6[1]), .D(
        \u_mux8/n4 ), .Q(sig_MUX_outMUX8) );
  OAI212 \u_decoder/iq_demod/U30  ( .A(\u_decoder/iq_demod/n59 ), .B(
        sig_DEMUX_outDEMUX1[0]), .C(n1961), .Q(\u_decoder/iq_demod/n71 ) );
  OAI212 \u_decoder/fir_filter/U900  ( .A(n860), .B(n318), .C(
        \u_decoder/fir_filter/n1145 ), .Q(\u_decoder/fir_filter/n1447 ) );
  OAI212 \u_decoder/fir_filter/U898  ( .A(n883), .B(n324), .C(
        \u_decoder/fir_filter/n1144 ), .Q(\u_decoder/fir_filter/n1446 ) );
  OAI212 \u_decoder/fir_filter/U896  ( .A(n875), .B(n58), .C(
        \u_decoder/fir_filter/n1143 ), .Q(\u_decoder/fir_filter/n1445 ) );
  OAI212 \u_decoder/fir_filter/U894  ( .A(n875), .B(n1854), .C(
        \u_decoder/fir_filter/n1142 ), .Q(\u_decoder/fir_filter/n1444 ) );
  OAI212 \u_decoder/fir_filter/U892  ( .A(n875), .B(n108), .C(
        \u_decoder/fir_filter/n1141 ), .Q(\u_decoder/fir_filter/n1443 ) );
  OAI212 \u_decoder/fir_filter/U890  ( .A(n875), .B(n344), .C(
        \u_decoder/fir_filter/n1140 ), .Q(\u_decoder/fir_filter/n1442 ) );
  OAI212 \u_decoder/fir_filter/U888  ( .A(n875), .B(n2442), .C(
        \u_decoder/fir_filter/n1139 ), .Q(\u_decoder/fir_filter/n1441 ) );
  OAI212 \u_decoder/fir_filter/U886  ( .A(n876), .B(
        \u_decoder/fir_filter/dp_cluster_0/r164/PROD1[4] ), .C(
        \u_decoder/fir_filter/n1138 ), .Q(\u_decoder/fir_filter/n1440 ) );
  OAI212 \u_decoder/fir_filter/U884  ( .A(n876), .B(n1859), .C(
        \u_decoder/fir_filter/n1137 ), .Q(\u_decoder/fir_filter/n1439 ) );
  OAI212 \u_decoder/fir_filter/U882  ( .A(n876), .B(n366), .C(
        \u_decoder/fir_filter/n1136 ), .Q(\u_decoder/fir_filter/n1438 ) );
  OAI212 \u_decoder/fir_filter/U880  ( .A(n876), .B(n59), .C(
        \u_decoder/fir_filter/n1135 ), .Q(\u_decoder/fir_filter/n1437 ) );
  OAI212 \u_decoder/fir_filter/U878  ( .A(n876), .B(n51), .C(
        \u_decoder/fir_filter/n1134 ), .Q(\u_decoder/fir_filter/n1436 ) );
  OAI212 \u_decoder/fir_filter/U869  ( .A(n876), .B(n316), .C(
        \u_decoder/fir_filter/n1130 ), .Q(\u_decoder/fir_filter/n1432 ) );
  OAI212 \u_decoder/fir_filter/U867  ( .A(n876), .B(n322), .C(
        \u_decoder/fir_filter/n1129 ), .Q(\u_decoder/fir_filter/n1431 ) );
  OAI212 \u_decoder/fir_filter/U865  ( .A(n877), .B(n328), .C(
        \u_decoder/fir_filter/n1128 ), .Q(\u_decoder/fir_filter/n1430 ) );
  OAI212 \u_decoder/fir_filter/U863  ( .A(n877), .B(n334), .C(
        \u_decoder/fir_filter/n1127 ), .Q(\u_decoder/fir_filter/n1429 ) );
  OAI212 \u_decoder/fir_filter/U861  ( .A(n877), .B(n66), .C(
        \u_decoder/fir_filter/n1126 ), .Q(\u_decoder/fir_filter/n1428 ) );
  OAI212 \u_decoder/fir_filter/U859  ( .A(n877), .B(n346), .C(
        \u_decoder/fir_filter/n1125 ), .Q(\u_decoder/fir_filter/n1427 ) );
  OAI212 \u_decoder/fir_filter/U857  ( .A(n877), .B(n2457), .C(
        \u_decoder/fir_filter/n1124 ), .Q(\u_decoder/fir_filter/n1426 ) );
  OAI212 \u_decoder/fir_filter/U855  ( .A(n877), .B(
        \u_decoder/fir_filter/dp_cluster_0/r165/PROD1[5] ), .C(
        \u_decoder/fir_filter/n1123 ), .Q(\u_decoder/fir_filter/n1425 ) );
  OAI212 \u_decoder/fir_filter/U853  ( .A(n877), .B(n1807), .C(
        \u_decoder/fir_filter/n1122 ), .Q(\u_decoder/fir_filter/n1424 ) );
  OAI212 \u_decoder/fir_filter/U851  ( .A(n878), .B(n362), .C(
        \u_decoder/fir_filter/n1121 ), .Q(\u_decoder/fir_filter/n1423 ) );
  OAI212 \u_decoder/fir_filter/U849  ( .A(n878), .B(n53), .C(
        \u_decoder/fir_filter/n1120 ), .Q(\u_decoder/fir_filter/n1422 ) );
  OAI212 \u_decoder/fir_filter/U847  ( .A(n878), .B(n59), .C(
        \u_decoder/fir_filter/n1119 ), .Q(\u_decoder/fir_filter/n1421 ) );
  OAI212 \u_decoder/fir_filter/U845  ( .A(n878), .B(n51), .C(
        \u_decoder/fir_filter/n1118 ), .Q(\u_decoder/fir_filter/n1420 ) );
  OAI212 \u_decoder/fir_filter/U836  ( .A(n878), .B(n348), .C(
        \u_decoder/fir_filter/n1114 ), .Q(\u_decoder/fir_filter/n1416 ) );
  OAI212 \u_decoder/fir_filter/U834  ( .A(n878), .B(n340), .C(
        \u_decoder/fir_filter/n1113 ), .Q(\u_decoder/fir_filter/n1415 ) );
  OAI212 \u_decoder/fir_filter/U832  ( .A(n878), .B(n326), .C(
        \u_decoder/fir_filter/n1112 ), .Q(\u_decoder/fir_filter/n1414 ) );
  OAI212 \u_decoder/fir_filter/U830  ( .A(n879), .B(n327), .C(
        \u_decoder/fir_filter/n1111 ), .Q(\u_decoder/fir_filter/n1413 ) );
  OAI212 \u_decoder/fir_filter/U828  ( .A(n879), .B(n1813), .C(
        \u_decoder/fir_filter/n1110 ), .Q(\u_decoder/fir_filter/n1412 ) );
  OAI212 \u_decoder/fir_filter/U826  ( .A(n879), .B(n355), .C(
        \u_decoder/fir_filter/n1109 ), .Q(\u_decoder/fir_filter/n1411 ) );
  OAI212 \u_decoder/fir_filter/U824  ( .A(n879), .B(n1815), .C(
        \u_decoder/fir_filter/n1108 ), .Q(\u_decoder/fir_filter/n1410 ) );
  OAI212 \u_decoder/fir_filter/U822  ( .A(n879), .B(n1816), .C(
        \u_decoder/fir_filter/n1107 ), .Q(\u_decoder/fir_filter/n1409 ) );
  OAI212 \u_decoder/fir_filter/U820  ( .A(n879), .B(n1817), .C(
        \u_decoder/fir_filter/n1106 ), .Q(\u_decoder/fir_filter/n1408 ) );
  OAI212 \u_decoder/fir_filter/U818  ( .A(n879), .B(n360), .C(
        \u_decoder/fir_filter/n1105 ), .Q(\u_decoder/fir_filter/n1407 ) );
  OAI212 \u_decoder/fir_filter/U816  ( .A(n880), .B(n59), .C(
        \u_decoder/fir_filter/n1104 ), .Q(\u_decoder/fir_filter/n1406 ) );
  OAI212 \u_decoder/fir_filter/U814  ( .A(n880), .B(n51), .C(
        \u_decoder/fir_filter/n1103 ), .Q(\u_decoder/fir_filter/n1405 ) );
  OAI212 \u_decoder/fir_filter/U808  ( .A(n880), .B(n48), .C(
        \u_decoder/fir_filter/n1100 ), .Q(\u_decoder/fir_filter/n1402 ) );
  OAI212 \u_decoder/fir_filter/U806  ( .A(n880), .B(n336), .C(
        \u_decoder/fir_filter/n1099 ), .Q(\u_decoder/fir_filter/n1401 ) );
  OAI212 \u_decoder/fir_filter/U804  ( .A(n880), .B(n50), .C(
        \u_decoder/fir_filter/n1098 ), .Q(\u_decoder/fir_filter/n1400 ) );
  OAI212 \u_decoder/fir_filter/U802  ( .A(n880), .B(n56), .C(
        \u_decoder/fir_filter/n1097 ), .Q(\u_decoder/fir_filter/n1399 ) );
  OAI212 \u_decoder/fir_filter/U800  ( .A(n880), .B(n1844), .C(
        \u_decoder/fir_filter/n1096 ), .Q(\u_decoder/fir_filter/n1398 ) );
  OAI212 \u_decoder/fir_filter/U798  ( .A(n881), .B(n332), .C(
        \u_decoder/fir_filter/n1095 ), .Q(\u_decoder/fir_filter/n1397 ) );
  OAI212 \u_decoder/fir_filter/U796  ( .A(n881), .B(n1846), .C(
        \u_decoder/fir_filter/n1094 ), .Q(\u_decoder/fir_filter/n1396 ) );
  OAI212 \u_decoder/fir_filter/U794  ( .A(n881), .B(n354), .C(
        \u_decoder/fir_filter/n1093 ), .Q(\u_decoder/fir_filter/n1395 ) );
  OAI212 \u_decoder/fir_filter/U792  ( .A(n881), .B(n1847), .C(
        \u_decoder/fir_filter/n1092 ), .Q(\u_decoder/fir_filter/n1394 ) );
  OAI212 \u_decoder/fir_filter/U790  ( .A(n881), .B(n1848), .C(
        \u_decoder/fir_filter/n1091 ), .Q(\u_decoder/fir_filter/n1393 ) );
  OAI212 \u_decoder/fir_filter/U788  ( .A(n881), .B(n1849), .C(
        \u_decoder/fir_filter/n1090 ), .Q(\u_decoder/fir_filter/n1392 ) );
  OAI212 \u_decoder/fir_filter/U786  ( .A(n881), .B(n1850), .C(
        \u_decoder/fir_filter/n1089 ), .Q(\u_decoder/fir_filter/n1391 ) );
  OAI212 \u_decoder/fir_filter/U784  ( .A(n882), .B(n1851), .C(
        \u_decoder/fir_filter/n1088 ), .Q(\u_decoder/fir_filter/n1390 ) );
  OAI212 \u_decoder/fir_filter/U782  ( .A(n882), .B(n364), .C(
        \u_decoder/fir_filter/n1087 ), .Q(\u_decoder/fir_filter/n1389 ) );
  OAI212 \u_decoder/fir_filter/U780  ( .A(n882), .B(n51), .C(
        \u_decoder/fir_filter/n1086 ), .Q(\u_decoder/fir_filter/n1388 ) );
  OAI212 \u_decoder/fir_filter/U760  ( .A(n882), .B(n48), .C(
        \u_decoder/fir_filter/n1068 ), .Q(\u_decoder/fir_filter/n1386 ) );
  OAI212 \u_decoder/fir_filter/U758  ( .A(n882), .B(n336), .C(
        \u_decoder/fir_filter/n1067 ), .Q(\u_decoder/fir_filter/n1385 ) );
  OAI212 \u_decoder/fir_filter/U756  ( .A(n882), .B(n50), .C(
        \u_decoder/fir_filter/n1066 ), .Q(\u_decoder/fir_filter/n1384 ) );
  OAI212 \u_decoder/fir_filter/U754  ( .A(n882), .B(n56), .C(
        \u_decoder/fir_filter/n1065 ), .Q(\u_decoder/fir_filter/n1383 ) );
  OAI212 \u_decoder/fir_filter/U752  ( .A(n883), .B(n1844), .C(
        \u_decoder/fir_filter/n1064 ), .Q(\u_decoder/fir_filter/n1382 ) );
  OAI212 \u_decoder/fir_filter/U750  ( .A(n883), .B(n332), .C(
        \u_decoder/fir_filter/n1063 ), .Q(\u_decoder/fir_filter/n1381 ) );
  OAI212 \u_decoder/fir_filter/U748  ( .A(n883), .B(n1846), .C(
        \u_decoder/fir_filter/n1062 ), .Q(\u_decoder/fir_filter/n1380 ) );
  OAI212 \u_decoder/fir_filter/U746  ( .A(n883), .B(n354), .C(
        \u_decoder/fir_filter/n1061 ), .Q(\u_decoder/fir_filter/n1379 ) );
  OAI212 \u_decoder/fir_filter/U744  ( .A(n883), .B(n1847), .C(
        \u_decoder/fir_filter/n1060 ), .Q(\u_decoder/fir_filter/n1378 ) );
  OAI212 \u_decoder/fir_filter/U742  ( .A(n883), .B(n1848), .C(
        \u_decoder/fir_filter/n1059 ), .Q(\u_decoder/fir_filter/n1377 ) );
  OAI212 \u_decoder/fir_filter/U740  ( .A(n884), .B(n1849), .C(
        \u_decoder/fir_filter/n1058 ), .Q(\u_decoder/fir_filter/n1376 ) );
  OAI212 \u_decoder/fir_filter/U738  ( .A(n884), .B(n1850), .C(
        \u_decoder/fir_filter/n1057 ), .Q(\u_decoder/fir_filter/n1375 ) );
  OAI212 \u_decoder/fir_filter/U736  ( .A(n884), .B(n1851), .C(
        \u_decoder/fir_filter/n1056 ), .Q(\u_decoder/fir_filter/n1374 ) );
  OAI212 \u_decoder/fir_filter/U734  ( .A(n884), .B(n364), .C(
        \u_decoder/fir_filter/n1055 ), .Q(\u_decoder/fir_filter/n1373 ) );
  OAI212 \u_decoder/fir_filter/U732  ( .A(n884), .B(n51), .C(
        \u_decoder/fir_filter/n1054 ), .Q(\u_decoder/fir_filter/n1372 ) );
  OAI212 \u_decoder/fir_filter/U724  ( .A(n884), .B(n348), .C(
        \u_decoder/fir_filter/n1049 ), .Q(\u_decoder/fir_filter/n1368 ) );
  OAI212 \u_decoder/fir_filter/U722  ( .A(n884), .B(n340), .C(
        \u_decoder/fir_filter/n1048 ), .Q(\u_decoder/fir_filter/n1367 ) );
  OAI212 \u_decoder/fir_filter/U720  ( .A(n885), .B(n326), .C(
        \u_decoder/fir_filter/n1047 ), .Q(\u_decoder/fir_filter/n1366 ) );
  OAI212 \u_decoder/fir_filter/U718  ( .A(n885), .B(n327), .C(
        \u_decoder/fir_filter/n1046 ), .Q(\u_decoder/fir_filter/n1365 ) );
  OAI212 \u_decoder/fir_filter/U716  ( .A(n885), .B(n1813), .C(
        \u_decoder/fir_filter/n1045 ), .Q(\u_decoder/fir_filter/n1364 ) );
  OAI212 \u_decoder/fir_filter/U714  ( .A(n885), .B(n355), .C(
        \u_decoder/fir_filter/n1044 ), .Q(\u_decoder/fir_filter/n1363 ) );
  OAI212 \u_decoder/fir_filter/U712  ( .A(n885), .B(n1815), .C(
        \u_decoder/fir_filter/n1043 ), .Q(\u_decoder/fir_filter/n1362 ) );
  OAI212 \u_decoder/fir_filter/U710  ( .A(n885), .B(n1816), .C(
        \u_decoder/fir_filter/n1042 ), .Q(\u_decoder/fir_filter/n1361 ) );
  OAI212 \u_decoder/fir_filter/U708  ( .A(n885), .B(n1817), .C(
        \u_decoder/fir_filter/n1041 ), .Q(\u_decoder/fir_filter/n1360 ) );
  OAI212 \u_decoder/fir_filter/U706  ( .A(n886), .B(n360), .C(
        \u_decoder/fir_filter/n1040 ), .Q(\u_decoder/fir_filter/n1359 ) );
  OAI212 \u_decoder/fir_filter/U704  ( .A(n886), .B(n59), .C(
        \u_decoder/fir_filter/n1039 ), .Q(\u_decoder/fir_filter/n1358 ) );
  OAI212 \u_decoder/fir_filter/U702  ( .A(n886), .B(n51), .C(
        \u_decoder/fir_filter/n1038 ), .Q(\u_decoder/fir_filter/n1357 ) );
  OAI212 \u_decoder/fir_filter/U692  ( .A(n886), .B(n316), .C(
        \u_decoder/fir_filter/n1032 ), .Q(\u_decoder/fir_filter/n1352 ) );
  OAI212 \u_decoder/fir_filter/U690  ( .A(n886), .B(n322), .C(
        \u_decoder/fir_filter/n1031 ), .Q(\u_decoder/fir_filter/n1351 ) );
  OAI212 \u_decoder/fir_filter/U688  ( .A(n886), .B(n328), .C(
        \u_decoder/fir_filter/n1030 ), .Q(\u_decoder/fir_filter/n1350 ) );
  OAI212 \u_decoder/fir_filter/U686  ( .A(n886), .B(n334), .C(
        \u_decoder/fir_filter/n1029 ), .Q(\u_decoder/fir_filter/n1349 ) );
  OAI212 \u_decoder/fir_filter/U684  ( .A(n887), .B(n66), .C(
        \u_decoder/fir_filter/n1028 ), .Q(\u_decoder/fir_filter/n1348 ) );
  OAI212 \u_decoder/fir_filter/U682  ( .A(n887), .B(n346), .C(
        \u_decoder/fir_filter/n1027 ), .Q(\u_decoder/fir_filter/n1347 ) );
  OAI212 \u_decoder/fir_filter/U680  ( .A(n887), .B(n2457), .C(
        \u_decoder/fir_filter/n1026 ), .Q(\u_decoder/fir_filter/n1346 ) );
  OAI212 \u_decoder/fir_filter/U678  ( .A(n887), .B(
        \u_decoder/fir_filter/dp_cluster_0/r165/PROD1[5] ), .C(
        \u_decoder/fir_filter/n1025 ), .Q(\u_decoder/fir_filter/n1345 ) );
  OAI212 \u_decoder/fir_filter/U676  ( .A(n887), .B(n1807), .C(
        \u_decoder/fir_filter/n1024 ), .Q(\u_decoder/fir_filter/n1344 ) );
  OAI212 \u_decoder/fir_filter/U674  ( .A(n887), .B(n362), .C(
        \u_decoder/fir_filter/n1023 ), .Q(\u_decoder/fir_filter/n1343 ) );
  OAI212 \u_decoder/fir_filter/U672  ( .A(n887), .B(n53), .C(
        \u_decoder/fir_filter/n1022 ), .Q(\u_decoder/fir_filter/n1342 ) );
  OAI212 \u_decoder/fir_filter/U670  ( .A(n888), .B(n59), .C(
        \u_decoder/fir_filter/n1021 ), .Q(\u_decoder/fir_filter/n1341 ) );
  OAI212 \u_decoder/fir_filter/U668  ( .A(n888), .B(n51), .C(
        \u_decoder/fir_filter/n1020 ), .Q(\u_decoder/fir_filter/n1340 ) );
  OAI212 \u_decoder/fir_filter/U666  ( .A(n938), .B(
        \u_decoder/fir_filter/n412 ), .C(\u_decoder/fir_filter/n1019 ), .Q(
        \u_decoder/fir_filter/n1338 ) );
  OAI212 \u_decoder/fir_filter/U665  ( .A(n938), .B(
        \u_decoder/fir_filter/n413 ), .C(\u_decoder/fir_filter/n1019 ), .Q(
        \u_decoder/fir_filter/n1337 ) );
  OAI212 \u_decoder/fir_filter/U664  ( .A(n938), .B(
        \u_decoder/fir_filter/n414 ), .C(\u_decoder/fir_filter/n1019 ), .Q(
        \u_decoder/fir_filter/n1336 ) );
  OAI222 \u_decoder/fir_filter/U663  ( .A(n939), .B(
        \u_decoder/fir_filter/n415 ), .C(n860), .D(n318), .Q(
        \u_decoder/fir_filter/n1335 ) );
  OAI222 \u_decoder/fir_filter/U662  ( .A(n939), .B(
        \u_decoder/fir_filter/n416 ), .C(n859), .D(n324), .Q(
        \u_decoder/fir_filter/n1334 ) );
  OAI222 \u_decoder/fir_filter/U661  ( .A(n939), .B(
        \u_decoder/fir_filter/n417 ), .C(n860), .D(n58), .Q(
        \u_decoder/fir_filter/n1333 ) );
  OAI222 \u_decoder/fir_filter/U660  ( .A(n939), .B(
        \u_decoder/fir_filter/n418 ), .C(n860), .D(n1854), .Q(
        \u_decoder/fir_filter/n1332 ) );
  OAI222 \u_decoder/fir_filter/U659  ( .A(n939), .B(
        \u_decoder/fir_filter/n419 ), .C(n858), .D(n108), .Q(
        \u_decoder/fir_filter/n1331 ) );
  OAI222 \u_decoder/fir_filter/U658  ( .A(n939), .B(
        \u_decoder/fir_filter/n420 ), .C(n858), .D(n344), .Q(
        \u_decoder/fir_filter/n1330 ) );
  OAI222 \u_decoder/fir_filter/U657  ( .A(n940), .B(
        \u_decoder/fir_filter/n421 ), .C(n860), .D(n2442), .Q(
        \u_decoder/fir_filter/n1329 ) );
  OAI222 \u_decoder/fir_filter/U656  ( .A(n940), .B(
        \u_decoder/fir_filter/n422 ), .C(n858), .D(
        \u_decoder/fir_filter/dp_cluster_0/r164/PROD1[4] ), .Q(
        \u_decoder/fir_filter/n1328 ) );
  OAI222 \u_decoder/fir_filter/U655  ( .A(n940), .B(
        \u_decoder/fir_filter/n423 ), .C(n860), .D(n1859), .Q(
        \u_decoder/fir_filter/n1327 ) );
  OAI222 \u_decoder/fir_filter/U654  ( .A(n940), .B(
        \u_decoder/fir_filter/n424 ), .C(n857), .D(n366), .Q(
        \u_decoder/fir_filter/n1326 ) );
  OAI222 \u_decoder/fir_filter/U653  ( .A(n940), .B(
        \u_decoder/fir_filter/n425 ), .C(n858), .D(n59), .Q(
        \u_decoder/fir_filter/n1325 ) );
  OAI222 \u_decoder/fir_filter/U652  ( .A(n940), .B(
        \u_decoder/fir_filter/n426 ), .C(n859), .D(n51), .Q(
        \u_decoder/fir_filter/n1324 ) );
  OAI212 \u_decoder/fir_filter/U637  ( .A(n888), .B(
        \u_decoder/fir_filter/n412 ), .C(\u_decoder/fir_filter/n1011 ), .Q(
        \u_decoder/fir_filter/n1317 ) );
  OAI212 \u_decoder/fir_filter/U635  ( .A(n888), .B(
        \u_decoder/fir_filter/n413 ), .C(\u_decoder/fir_filter/n1010 ), .Q(
        \u_decoder/fir_filter/n1316 ) );
  OAI212 \u_decoder/fir_filter/U633  ( .A(n888), .B(
        \u_decoder/fir_filter/n414 ), .C(\u_decoder/fir_filter/n1009 ), .Q(
        \u_decoder/fir_filter/n1315 ) );
  OAI212 \u_decoder/fir_filter/U631  ( .A(n888), .B(
        \u_decoder/fir_filter/n415 ), .C(\u_decoder/fir_filter/n1008 ), .Q(
        \u_decoder/fir_filter/n1314 ) );
  OAI212 \u_decoder/fir_filter/U629  ( .A(n888), .B(
        \u_decoder/fir_filter/n416 ), .C(\u_decoder/fir_filter/n1007 ), .Q(
        \u_decoder/fir_filter/n1313 ) );
  OAI212 \u_decoder/fir_filter/U627  ( .A(n889), .B(
        \u_decoder/fir_filter/n417 ), .C(\u_decoder/fir_filter/n1006 ), .Q(
        \u_decoder/fir_filter/n1312 ) );
  OAI212 \u_decoder/fir_filter/U625  ( .A(n889), .B(
        \u_decoder/fir_filter/n418 ), .C(\u_decoder/fir_filter/n1005 ), .Q(
        \u_decoder/fir_filter/n1311 ) );
  OAI212 \u_decoder/fir_filter/U623  ( .A(n889), .B(
        \u_decoder/fir_filter/n419 ), .C(\u_decoder/fir_filter/n1004 ), .Q(
        \u_decoder/fir_filter/n1310 ) );
  OAI212 \u_decoder/fir_filter/U621  ( .A(n889), .B(
        \u_decoder/fir_filter/n420 ), .C(\u_decoder/fir_filter/n1003 ), .Q(
        \u_decoder/fir_filter/n1309 ) );
  OAI212 \u_decoder/fir_filter/U619  ( .A(n889), .B(
        \u_decoder/fir_filter/n421 ), .C(\u_decoder/fir_filter/n1002 ), .Q(
        \u_decoder/fir_filter/n1308 ) );
  OAI212 \u_decoder/fir_filter/U617  ( .A(n889), .B(
        \u_decoder/fir_filter/n422 ), .C(\u_decoder/fir_filter/n1001 ), .Q(
        \u_decoder/fir_filter/n1307 ) );
  OAI212 \u_decoder/fir_filter/U615  ( .A(n889), .B(
        \u_decoder/fir_filter/n423 ), .C(\u_decoder/fir_filter/n1000 ), .Q(
        \u_decoder/fir_filter/n1306 ) );
  OAI212 \u_decoder/fir_filter/U613  ( .A(n890), .B(
        \u_decoder/fir_filter/n424 ), .C(\u_decoder/fir_filter/n999 ), .Q(
        \u_decoder/fir_filter/n1305 ) );
  OAI212 \u_decoder/fir_filter/U611  ( .A(n890), .B(
        \u_decoder/fir_filter/n425 ), .C(\u_decoder/fir_filter/n998 ), .Q(
        \u_decoder/fir_filter/n1304 ) );
  OAI212 \u_decoder/fir_filter/U609  ( .A(n890), .B(
        \u_decoder/fir_filter/n426 ), .C(\u_decoder/fir_filter/n997 ), .Q(
        \u_decoder/fir_filter/n1303 ) );
  OAI212 \u_decoder/fir_filter/U455  ( .A(n890), .B(n319), .C(
        \u_decoder/fir_filter/n848 ), .Q(\u_decoder/fir_filter/n1299 ) );
  OAI212 \u_decoder/fir_filter/U453  ( .A(n890), .B(n325), .C(
        \u_decoder/fir_filter/n847 ), .Q(\u_decoder/fir_filter/n1298 ) );
  OAI212 \u_decoder/fir_filter/U451  ( .A(n890), .B(n57), .C(
        \u_decoder/fir_filter/n846 ), .Q(\u_decoder/fir_filter/n1297 ) );
  OAI212 \u_decoder/fir_filter/U449  ( .A(n890), .B(n1925), .C(
        \u_decoder/fir_filter/n845 ), .Q(\u_decoder/fir_filter/n1296 ) );
  OAI212 \u_decoder/fir_filter/U447  ( .A(n891), .B(n107), .C(
        \u_decoder/fir_filter/n844 ), .Q(\u_decoder/fir_filter/n1295 ) );
  OAI212 \u_decoder/fir_filter/U445  ( .A(n891), .B(n345), .C(
        \u_decoder/fir_filter/n843 ), .Q(\u_decoder/fir_filter/n1294 ) );
  OAI212 \u_decoder/fir_filter/U443  ( .A(n867), .B(n2355), .C(
        \u_decoder/fir_filter/n842 ), .Q(\u_decoder/fir_filter/n1293 ) );
  OAI212 \u_decoder/fir_filter/U441  ( .A(n861), .B(
        \u_decoder/fir_filter/dp_cluster_0/r177/PROD1[4] ), .C(
        \u_decoder/fir_filter/n841 ), .Q(\u_decoder/fir_filter/n1292 ) );
  OAI212 \u_decoder/fir_filter/U439  ( .A(n860), .B(n1930), .C(
        \u_decoder/fir_filter/n840 ), .Q(\u_decoder/fir_filter/n1291 ) );
  OAI212 \u_decoder/fir_filter/U437  ( .A(n863), .B(n367), .C(
        \u_decoder/fir_filter/n839 ), .Q(\u_decoder/fir_filter/n1290 ) );
  OAI212 \u_decoder/fir_filter/U435  ( .A(n863), .B(n60), .C(
        \u_decoder/fir_filter/n838 ), .Q(\u_decoder/fir_filter/n1289 ) );
  OAI212 \u_decoder/fir_filter/U433  ( .A(n861), .B(n52), .C(
        \u_decoder/fir_filter/n837 ), .Q(\u_decoder/fir_filter/n1288 ) );
  OAI212 \u_decoder/fir_filter/U424  ( .A(n861), .B(n317), .C(
        \u_decoder/fir_filter/n833 ), .Q(\u_decoder/fir_filter/n1284 ) );
  OAI212 \u_decoder/fir_filter/U422  ( .A(n862), .B(n323), .C(
        \u_decoder/fir_filter/n832 ), .Q(\u_decoder/fir_filter/n1283 ) );
  OAI212 \u_decoder/fir_filter/U420  ( .A(n861), .B(n331), .C(
        \u_decoder/fir_filter/n831 ), .Q(\u_decoder/fir_filter/n1282 ) );
  OAI212 \u_decoder/fir_filter/U418  ( .A(n861), .B(n335), .C(
        \u_decoder/fir_filter/n830 ), .Q(\u_decoder/fir_filter/n1281 ) );
  OAI212 \u_decoder/fir_filter/U416  ( .A(n862), .B(n65), .C(
        \u_decoder/fir_filter/n829 ), .Q(\u_decoder/fir_filter/n1280 ) );
  OAI212 \u_decoder/fir_filter/U414  ( .A(n862), .B(n347), .C(
        \u_decoder/fir_filter/n828 ), .Q(\u_decoder/fir_filter/n1279 ) );
  OAI212 \u_decoder/fir_filter/U412  ( .A(n861), .B(n2370), .C(
        \u_decoder/fir_filter/n827 ), .Q(\u_decoder/fir_filter/n1278 ) );
  OAI212 \u_decoder/fir_filter/U410  ( .A(n862), .B(
        \u_decoder/fir_filter/dp_cluster_0/r178/PROD1[5] ), .C(
        \u_decoder/fir_filter/n826 ), .Q(\u_decoder/fir_filter/n1277 ) );
  OAI212 \u_decoder/fir_filter/U408  ( .A(n861), .B(n1878), .C(
        \u_decoder/fir_filter/n825 ), .Q(\u_decoder/fir_filter/n1276 ) );
  OAI212 \u_decoder/fir_filter/U406  ( .A(n862), .B(n363), .C(
        \u_decoder/fir_filter/n824 ), .Q(\u_decoder/fir_filter/n1275 ) );
  OAI212 \u_decoder/fir_filter/U404  ( .A(n863), .B(n54), .C(
        \u_decoder/fir_filter/n823 ), .Q(\u_decoder/fir_filter/n1274 ) );
  OAI212 \u_decoder/fir_filter/U402  ( .A(n862), .B(n60), .C(
        \u_decoder/fir_filter/n822 ), .Q(\u_decoder/fir_filter/n1273 ) );
  OAI212 \u_decoder/fir_filter/U400  ( .A(n862), .B(n52), .C(
        \u_decoder/fir_filter/n821 ), .Q(\u_decoder/fir_filter/n1272 ) );
  OAI212 \u_decoder/fir_filter/U391  ( .A(n863), .B(n349), .C(
        \u_decoder/fir_filter/n817 ), .Q(\u_decoder/fir_filter/n1268 ) );
  OAI212 \u_decoder/fir_filter/U389  ( .A(n863), .B(n341), .C(
        \u_decoder/fir_filter/n816 ), .Q(\u_decoder/fir_filter/n1267 ) );
  OAI212 \u_decoder/fir_filter/U387  ( .A(n863), .B(n329), .C(
        \u_decoder/fir_filter/n815 ), .Q(\u_decoder/fir_filter/n1266 ) );
  OAI212 \u_decoder/fir_filter/U385  ( .A(n863), .B(n330), .C(
        \u_decoder/fir_filter/n814 ), .Q(\u_decoder/fir_filter/n1265 ) );
  OAI212 \u_decoder/fir_filter/U383  ( .A(n864), .B(n1884), .C(
        \u_decoder/fir_filter/n813 ), .Q(\u_decoder/fir_filter/n1264 ) );
  OAI212 \u_decoder/fir_filter/U381  ( .A(n864), .B(n357), .C(
        \u_decoder/fir_filter/n812 ), .Q(\u_decoder/fir_filter/n1263 ) );
  OAI212 \u_decoder/fir_filter/U379  ( .A(n864), .B(n1886), .C(
        \u_decoder/fir_filter/n811 ), .Q(\u_decoder/fir_filter/n1262 ) );
  OAI212 \u_decoder/fir_filter/U377  ( .A(n864), .B(n1887), .C(
        \u_decoder/fir_filter/n810 ), .Q(\u_decoder/fir_filter/n1261 ) );
  OAI212 \u_decoder/fir_filter/U375  ( .A(n864), .B(n1888), .C(
        \u_decoder/fir_filter/n809 ), .Q(\u_decoder/fir_filter/n1260 ) );
  OAI212 \u_decoder/fir_filter/U373  ( .A(n864), .B(n361), .C(
        \u_decoder/fir_filter/n808 ), .Q(\u_decoder/fir_filter/n1259 ) );
  OAI212 \u_decoder/fir_filter/U371  ( .A(n864), .B(n60), .C(
        \u_decoder/fir_filter/n807 ), .Q(\u_decoder/fir_filter/n1258 ) );
  OAI212 \u_decoder/fir_filter/U369  ( .A(n865), .B(n52), .C(
        \u_decoder/fir_filter/n806 ), .Q(\u_decoder/fir_filter/n1257 ) );
  OAI212 \u_decoder/fir_filter/U363  ( .A(n865), .B(n47), .C(
        \u_decoder/fir_filter/n803 ), .Q(\u_decoder/fir_filter/n1254 ) );
  OAI212 \u_decoder/fir_filter/U361  ( .A(n865), .B(n337), .C(
        \u_decoder/fir_filter/n802 ), .Q(\u_decoder/fir_filter/n1253 ) );
  OAI212 \u_decoder/fir_filter/U359  ( .A(n865), .B(n49), .C(
        \u_decoder/fir_filter/n801 ), .Q(\u_decoder/fir_filter/n1252 ) );
  OAI212 \u_decoder/fir_filter/U357  ( .A(n865), .B(n55), .C(
        \u_decoder/fir_filter/n800 ), .Q(\u_decoder/fir_filter/n1251 ) );
  OAI212 \u_decoder/fir_filter/U355  ( .A(n865), .B(n1915), .C(
        \u_decoder/fir_filter/n799 ), .Q(\u_decoder/fir_filter/n1250 ) );
  OAI212 \u_decoder/fir_filter/U353  ( .A(n865), .B(n333), .C(
        \u_decoder/fir_filter/n798 ), .Q(\u_decoder/fir_filter/n1249 ) );
  OAI212 \u_decoder/fir_filter/U351  ( .A(n866), .B(n1917), .C(
        \u_decoder/fir_filter/n797 ), .Q(\u_decoder/fir_filter/n1248 ) );
  OAI212 \u_decoder/fir_filter/U349  ( .A(n866), .B(n356), .C(
        \u_decoder/fir_filter/n796 ), .Q(\u_decoder/fir_filter/n1247 ) );
  OAI212 \u_decoder/fir_filter/U347  ( .A(n866), .B(n1918), .C(
        \u_decoder/fir_filter/n795 ), .Q(\u_decoder/fir_filter/n1246 ) );
  OAI212 \u_decoder/fir_filter/U345  ( .A(n866), .B(n1919), .C(
        \u_decoder/fir_filter/n794 ), .Q(\u_decoder/fir_filter/n1245 ) );
  OAI212 \u_decoder/fir_filter/U343  ( .A(n866), .B(n1920), .C(
        \u_decoder/fir_filter/n793 ), .Q(\u_decoder/fir_filter/n1244 ) );
  OAI212 \u_decoder/fir_filter/U341  ( .A(n866), .B(n1921), .C(
        \u_decoder/fir_filter/n792 ), .Q(\u_decoder/fir_filter/n1243 ) );
  OAI212 \u_decoder/fir_filter/U339  ( .A(n866), .B(n1922), .C(
        \u_decoder/fir_filter/n791 ), .Q(\u_decoder/fir_filter/n1242 ) );
  OAI212 \u_decoder/fir_filter/U337  ( .A(n867), .B(n365), .C(
        \u_decoder/fir_filter/n790 ), .Q(\u_decoder/fir_filter/n1241 ) );
  OAI212 \u_decoder/fir_filter/U335  ( .A(n867), .B(n52), .C(
        \u_decoder/fir_filter/n789 ), .Q(\u_decoder/fir_filter/n1240 ) );
  OAI212 \u_decoder/fir_filter/U315  ( .A(n867), .B(n47), .C(
        \u_decoder/fir_filter/n771 ), .Q(\u_decoder/fir_filter/n1238 ) );
  OAI212 \u_decoder/fir_filter/U313  ( .A(n867), .B(n337), .C(
        \u_decoder/fir_filter/n770 ), .Q(\u_decoder/fir_filter/n1237 ) );
  OAI212 \u_decoder/fir_filter/U311  ( .A(n867), .B(n49), .C(
        \u_decoder/fir_filter/n769 ), .Q(\u_decoder/fir_filter/n1236 ) );
  OAI212 \u_decoder/fir_filter/U309  ( .A(n867), .B(n55), .C(
        \u_decoder/fir_filter/n768 ), .Q(\u_decoder/fir_filter/n1235 ) );
  OAI212 \u_decoder/fir_filter/U307  ( .A(n868), .B(n1915), .C(
        \u_decoder/fir_filter/n767 ), .Q(\u_decoder/fir_filter/n1234 ) );
  OAI212 \u_decoder/fir_filter/U305  ( .A(n868), .B(n333), .C(
        \u_decoder/fir_filter/n766 ), .Q(\u_decoder/fir_filter/n1233 ) );
  OAI212 \u_decoder/fir_filter/U303  ( .A(n868), .B(n1917), .C(
        \u_decoder/fir_filter/n765 ), .Q(\u_decoder/fir_filter/n1232 ) );
  OAI212 \u_decoder/fir_filter/U301  ( .A(n868), .B(n356), .C(
        \u_decoder/fir_filter/n764 ), .Q(\u_decoder/fir_filter/n1231 ) );
  OAI212 \u_decoder/fir_filter/U299  ( .A(n868), .B(n1918), .C(
        \u_decoder/fir_filter/n763 ), .Q(\u_decoder/fir_filter/n1230 ) );
  OAI212 \u_decoder/fir_filter/U297  ( .A(n868), .B(n1919), .C(
        \u_decoder/fir_filter/n762 ), .Q(\u_decoder/fir_filter/n1229 ) );
  OAI212 \u_decoder/fir_filter/U295  ( .A(n868), .B(n1920), .C(
        \u_decoder/fir_filter/n761 ), .Q(\u_decoder/fir_filter/n1228 ) );
  OAI212 \u_decoder/fir_filter/U293  ( .A(n869), .B(n1921), .C(
        \u_decoder/fir_filter/n760 ), .Q(\u_decoder/fir_filter/n1227 ) );
  OAI212 \u_decoder/fir_filter/U291  ( .A(n869), .B(n1922), .C(
        \u_decoder/fir_filter/n759 ), .Q(\u_decoder/fir_filter/n1226 ) );
  OAI212 \u_decoder/fir_filter/U289  ( .A(n869), .B(n365), .C(
        \u_decoder/fir_filter/n758 ), .Q(\u_decoder/fir_filter/n1225 ) );
  OAI212 \u_decoder/fir_filter/U287  ( .A(n869), .B(n52), .C(
        \u_decoder/fir_filter/n757 ), .Q(\u_decoder/fir_filter/n1224 ) );
  OAI212 \u_decoder/fir_filter/U279  ( .A(n869), .B(n349), .C(
        \u_decoder/fir_filter/n752 ), .Q(\u_decoder/fir_filter/n1220 ) );
  OAI212 \u_decoder/fir_filter/U277  ( .A(n869), .B(n341), .C(
        \u_decoder/fir_filter/n751 ), .Q(\u_decoder/fir_filter/n1219 ) );
  OAI212 \u_decoder/fir_filter/U275  ( .A(n869), .B(n329), .C(
        \u_decoder/fir_filter/n750 ), .Q(\u_decoder/fir_filter/n1218 ) );
  OAI212 \u_decoder/fir_filter/U273  ( .A(n870), .B(n330), .C(
        \u_decoder/fir_filter/n749 ), .Q(\u_decoder/fir_filter/n1217 ) );
  OAI212 \u_decoder/fir_filter/U271  ( .A(n870), .B(n1884), .C(
        \u_decoder/fir_filter/n748 ), .Q(\u_decoder/fir_filter/n1216 ) );
  OAI212 \u_decoder/fir_filter/U269  ( .A(n870), .B(n357), .C(
        \u_decoder/fir_filter/n747 ), .Q(\u_decoder/fir_filter/n1215 ) );
  OAI212 \u_decoder/fir_filter/U267  ( .A(n870), .B(n1886), .C(
        \u_decoder/fir_filter/n746 ), .Q(\u_decoder/fir_filter/n1214 ) );
  OAI212 \u_decoder/fir_filter/U265  ( .A(n870), .B(n1887), .C(
        \u_decoder/fir_filter/n745 ), .Q(\u_decoder/fir_filter/n1213 ) );
  OAI212 \u_decoder/fir_filter/U263  ( .A(n870), .B(n1888), .C(
        \u_decoder/fir_filter/n744 ), .Q(\u_decoder/fir_filter/n1212 ) );
  OAI212 \u_decoder/fir_filter/U261  ( .A(n870), .B(n361), .C(
        \u_decoder/fir_filter/n743 ), .Q(\u_decoder/fir_filter/n1211 ) );
  OAI212 \u_decoder/fir_filter/U259  ( .A(n871), .B(n60), .C(
        \u_decoder/fir_filter/n742 ), .Q(\u_decoder/fir_filter/n1210 ) );
  OAI212 \u_decoder/fir_filter/U257  ( .A(n871), .B(n52), .C(
        \u_decoder/fir_filter/n741 ), .Q(\u_decoder/fir_filter/n1209 ) );
  OAI212 \u_decoder/fir_filter/U247  ( .A(n871), .B(n317), .C(
        \u_decoder/fir_filter/n735 ), .Q(\u_decoder/fir_filter/n1204 ) );
  OAI212 \u_decoder/fir_filter/U245  ( .A(n871), .B(n323), .C(
        \u_decoder/fir_filter/n734 ), .Q(\u_decoder/fir_filter/n1203 ) );
  OAI212 \u_decoder/fir_filter/U243  ( .A(n871), .B(n331), .C(
        \u_decoder/fir_filter/n733 ), .Q(\u_decoder/fir_filter/n1202 ) );
  OAI212 \u_decoder/fir_filter/U241  ( .A(n871), .B(n335), .C(
        \u_decoder/fir_filter/n732 ), .Q(\u_decoder/fir_filter/n1201 ) );
  OAI212 \u_decoder/fir_filter/U239  ( .A(n871), .B(n65), .C(
        \u_decoder/fir_filter/n731 ), .Q(\u_decoder/fir_filter/n1200 ) );
  OAI212 \u_decoder/fir_filter/U237  ( .A(n872), .B(n347), .C(
        \u_decoder/fir_filter/n730 ), .Q(\u_decoder/fir_filter/n1199 ) );
  OAI212 \u_decoder/fir_filter/U235  ( .A(n872), .B(n2370), .C(
        \u_decoder/fir_filter/n729 ), .Q(\u_decoder/fir_filter/n1198 ) );
  OAI212 \u_decoder/fir_filter/U233  ( .A(n872), .B(
        \u_decoder/fir_filter/dp_cluster_0/r178/PROD1[5] ), .C(
        \u_decoder/fir_filter/n728 ), .Q(\u_decoder/fir_filter/n1197 ) );
  OAI212 \u_decoder/fir_filter/U231  ( .A(n872), .B(n1878), .C(
        \u_decoder/fir_filter/n727 ), .Q(\u_decoder/fir_filter/n1196 ) );
  OAI212 \u_decoder/fir_filter/U229  ( .A(n872), .B(n363), .C(
        \u_decoder/fir_filter/n726 ), .Q(\u_decoder/fir_filter/n1195 ) );
  OAI212 \u_decoder/fir_filter/U227  ( .A(n872), .B(n54), .C(
        \u_decoder/fir_filter/n725 ), .Q(\u_decoder/fir_filter/n1194 ) );
  OAI212 \u_decoder/fir_filter/U225  ( .A(n872), .B(n60), .C(
        \u_decoder/fir_filter/n724 ), .Q(\u_decoder/fir_filter/n1193 ) );
  OAI212 \u_decoder/fir_filter/U223  ( .A(n873), .B(n52), .C(
        \u_decoder/fir_filter/n723 ), .Q(\u_decoder/fir_filter/n1192 ) );
  OAI212 \u_decoder/fir_filter/U221  ( .A(n939), .B(
        \u_decoder/fir_filter/n428 ), .C(\u_decoder/fir_filter/n722 ), .Q(
        \u_decoder/fir_filter/n1190 ) );
  OAI212 \u_decoder/fir_filter/U220  ( .A(n939), .B(
        \u_decoder/fir_filter/n429 ), .C(\u_decoder/fir_filter/n722 ), .Q(
        \u_decoder/fir_filter/n1189 ) );
  OAI212 \u_decoder/fir_filter/U219  ( .A(n939), .B(
        \u_decoder/fir_filter/n430 ), .C(\u_decoder/fir_filter/n722 ), .Q(
        \u_decoder/fir_filter/n1188 ) );
  OAI222 \u_decoder/fir_filter/U218  ( .A(n940), .B(
        \u_decoder/fir_filter/n431 ), .C(n859), .D(n319), .Q(
        \u_decoder/fir_filter/n1187 ) );
  OAI222 \u_decoder/fir_filter/U217  ( .A(n940), .B(
        \u_decoder/fir_filter/n432 ), .C(n858), .D(n325), .Q(
        \u_decoder/fir_filter/n1186 ) );
  OAI222 \u_decoder/fir_filter/U216  ( .A(n940), .B(
        \u_decoder/fir_filter/n433 ), .C(n859), .D(n57), .Q(
        \u_decoder/fir_filter/n1185 ) );
  OAI222 \u_decoder/fir_filter/U215  ( .A(n940), .B(
        \u_decoder/fir_filter/n434 ), .C(n859), .D(n1925), .Q(
        \u_decoder/fir_filter/n1184 ) );
  OAI222 \u_decoder/fir_filter/U214  ( .A(n941), .B(
        \u_decoder/fir_filter/n435 ), .C(n857), .D(n107), .Q(
        \u_decoder/fir_filter/n1183 ) );
  OAI222 \u_decoder/fir_filter/U213  ( .A(n941), .B(
        \u_decoder/fir_filter/n436 ), .C(n859), .D(n345), .Q(
        \u_decoder/fir_filter/n1182 ) );
  OAI222 \u_decoder/fir_filter/U212  ( .A(n941), .B(
        \u_decoder/fir_filter/n437 ), .C(n859), .D(n2355), .Q(
        \u_decoder/fir_filter/n1181 ) );
  OAI222 \u_decoder/fir_filter/U211  ( .A(n941), .B(
        \u_decoder/fir_filter/n438 ), .C(n857), .D(
        \u_decoder/fir_filter/dp_cluster_0/r177/PROD1[4] ), .Q(
        \u_decoder/fir_filter/n1180 ) );
  OAI222 \u_decoder/fir_filter/U210  ( .A(n941), .B(
        \u_decoder/fir_filter/n439 ), .C(n857), .D(n1930), .Q(
        \u_decoder/fir_filter/n1179 ) );
  OAI222 \u_decoder/fir_filter/U209  ( .A(n941), .B(
        \u_decoder/fir_filter/n440 ), .C(n858), .D(n367), .Q(
        \u_decoder/fir_filter/n1178 ) );
  OAI222 \u_decoder/fir_filter/U208  ( .A(n941), .B(
        \u_decoder/fir_filter/n441 ), .C(n857), .D(n60), .Q(
        \u_decoder/fir_filter/n1177 ) );
  OAI222 \u_decoder/fir_filter/U207  ( .A(n941), .B(
        \u_decoder/fir_filter/n442 ), .C(n858), .D(n52), .Q(
        \u_decoder/fir_filter/n1176 ) );
  OAI212 \u_decoder/fir_filter/U192  ( .A(n873), .B(
        \u_decoder/fir_filter/n428 ), .C(\u_decoder/fir_filter/n713 ), .Q(
        \u_decoder/fir_filter/n1169 ) );
  OAI212 \u_decoder/fir_filter/U190  ( .A(n873), .B(
        \u_decoder/fir_filter/n429 ), .C(\u_decoder/fir_filter/n712 ), .Q(
        \u_decoder/fir_filter/n1168 ) );
  OAI212 \u_decoder/fir_filter/U188  ( .A(n873), .B(
        \u_decoder/fir_filter/n430 ), .C(\u_decoder/fir_filter/n711 ), .Q(
        \u_decoder/fir_filter/n1167 ) );
  OAI212 \u_decoder/fir_filter/U186  ( .A(n873), .B(
        \u_decoder/fir_filter/n431 ), .C(\u_decoder/fir_filter/n710 ), .Q(
        \u_decoder/fir_filter/n1166 ) );
  OAI212 \u_decoder/fir_filter/U184  ( .A(n873), .B(
        \u_decoder/fir_filter/n432 ), .C(\u_decoder/fir_filter/n709 ), .Q(
        \u_decoder/fir_filter/n1165 ) );
  OAI212 \u_decoder/fir_filter/U182  ( .A(n873), .B(
        \u_decoder/fir_filter/n433 ), .C(\u_decoder/fir_filter/n708 ), .Q(
        \u_decoder/fir_filter/n1164 ) );
  OAI212 \u_decoder/fir_filter/U180  ( .A(n874), .B(
        \u_decoder/fir_filter/n434 ), .C(\u_decoder/fir_filter/n707 ), .Q(
        \u_decoder/fir_filter/n1163 ) );
  OAI212 \u_decoder/fir_filter/U178  ( .A(n874), .B(
        \u_decoder/fir_filter/n435 ), .C(\u_decoder/fir_filter/n706 ), .Q(
        \u_decoder/fir_filter/n1162 ) );
  OAI212 \u_decoder/fir_filter/U176  ( .A(n874), .B(
        \u_decoder/fir_filter/n436 ), .C(\u_decoder/fir_filter/n705 ), .Q(
        \u_decoder/fir_filter/n1161 ) );
  OAI212 \u_decoder/fir_filter/U174  ( .A(n874), .B(
        \u_decoder/fir_filter/n437 ), .C(\u_decoder/fir_filter/n704 ), .Q(
        \u_decoder/fir_filter/n1160 ) );
  OAI212 \u_decoder/fir_filter/U172  ( .A(n874), .B(
        \u_decoder/fir_filter/n438 ), .C(\u_decoder/fir_filter/n703 ), .Q(
        \u_decoder/fir_filter/n1159 ) );
  OAI212 \u_decoder/fir_filter/U170  ( .A(n874), .B(
        \u_decoder/fir_filter/n439 ), .C(\u_decoder/fir_filter/n702 ), .Q(
        \u_decoder/fir_filter/n1158 ) );
  OAI212 \u_decoder/fir_filter/U168  ( .A(n874), .B(
        \u_decoder/fir_filter/n440 ), .C(\u_decoder/fir_filter/n701 ), .Q(
        \u_decoder/fir_filter/n1157 ) );
  OAI212 \u_decoder/fir_filter/U166  ( .A(n875), .B(
        \u_decoder/fir_filter/n441 ), .C(\u_decoder/fir_filter/n700 ), .Q(
        \u_decoder/fir_filter/n1156 ) );
  OAI212 \u_decoder/fir_filter/U164  ( .A(n875), .B(
        \u_decoder/fir_filter/n442 ), .C(\u_decoder/fir_filter/n699 ), .Q(
        \u_decoder/fir_filter/n1155 ) );
  OAI222 \u_cdr/phd1/U10  ( .A(\u_cdr/phd1/n16 ), .B(\u_cdr/phd1/n9 ), .C(
        \u_cdr/phd1/n19 ), .D(\u_cdr/phd1/n18 ), .Q(\u_cdr/phd1/n21 ) );
  OAI222 \u_cdr/phd1/U8  ( .A(\u_cdr/phd1/n16 ), .B(\u_cdr/phd1/n10 ), .C(
        \u_cdr/phd1/n17 ), .D(\u_cdr/phd1/n18 ), .Q(\u_cdr/phd1/n20 ) );
  OAI222 \u_cdr/dec1/U9  ( .A(n308), .B(\u_cdr/dir ), .C(\u_cdr/dec1/n20 ), 
        .D(\u_cdr/dec1/w_en_dec ), .Q(\u_cdr/dec1/n25 ) );
  OAI212 \u_decoder/iq_demod/cossin_dig/U31  ( .A(
        \u_decoder/iq_demod/cossin_dig/n47 ), .B(
        \u_decoder/iq_demod/cossin_dig/N20 ), .C(
        \u_decoder/iq_demod/cossin_dig/counter [2]), .Q(
        \u_decoder/iq_demod/cossin_dig/n46 ) );
  OAI222 \u_decoder/iq_demod/cossin_dig/U20  ( .A(
        \u_decoder/iq_demod/cossin_dig/n21 ), .B(
        \u_decoder/iq_demod/cossin_dig/n41 ), .C(
        \u_decoder/iq_demod/cossin_dig/N55 ), .D(
        \u_decoder/iq_demod/cossin_dig/n40 ), .Q(
        \u_decoder/iq_demod/cossin_dig/n53 ) );
  OAI222 \u_decoder/iq_demod/cossin_dig/U18  ( .A(
        \u_decoder/iq_demod/cossin_dig/n19 ), .B(n1504), .C(
        \u_decoder/iq_demod/cossin_dig/n21 ), .D(
        \u_decoder/iq_demod/cossin_dig/n40 ), .Q(
        \u_decoder/iq_demod/cossin_dig/n52 ) );
  OAI212 \u_decoder/iq_demod/cossin_dig/U10  ( .A(
        \u_decoder/iq_demod/cossin_dig/N55 ), .B(
        \u_decoder/iq_demod/cossin_dig/n31 ), .C(
        \u_decoder/iq_demod/cossin_dig/n32 ), .Q(
        \u_decoder/iq_demod/cossin_dig/n51 ) );
  OAI222 \u_mux7/mux3/U1  ( .A(n2685), .B(n1688), .C(in_MUX_inSEL6[1]), .D(
        n2686), .Q(sig_MUX_outMUX7[3]) );
  OAI222 \u_mux7/mux2/U1  ( .A(n2683), .B(n1688), .C(in_MUX_inSEL6[1]), .D(
        n2684), .Q(sig_MUX_outMUX7[2]) );
  OAI222 \u_mux7/mux1/U1  ( .A(n2681), .B(n1688), .C(in_MUX_inSEL6[1]), .D(
        n2682), .Q(sig_MUX_outMUX7[1]) );
  OAI222 \u_mux7/mux0/U1  ( .A(n2679), .B(n1688), .C(in_MUX_inSEL6[1]), .D(
        n2680), .Q(sig_MUX_outMUX7[0]) );
  OAI222 \u_mux6/mux3/U1  ( .A(n2677), .B(n1688), .C(in_MUX_inSEL6[1]), .D(
        n2678), .Q(sig_MUX_outMUX6[3]) );
  OAI222 \u_mux6/mux2/U1  ( .A(n2675), .B(n1688), .C(in_MUX_inSEL6[1]), .D(
        n2676), .Q(sig_MUX_outMUX6[2]) );
  OAI222 \u_mux6/mux1/U1  ( .A(n2673), .B(n1688), .C(in_MUX_inSEL6[1]), .D(
        n2674), .Q(sig_MUX_outMUX6[1]) );
  OAI222 \u_mux6/mux0/U1  ( .A(n2671), .B(n1688), .C(in_MUX_inSEL6[1]), .D(
        n2672), .Q(sig_MUX_outMUX6[0]) );
  OAI222 \u_mux10/mux3/U1  ( .A(n2669), .B(n1690), .C(in_MUX_inSEL9[1]), .D(
        n2670), .Q(out_MUX_outMUX10[3]) );
  OAI222 \u_mux10/mux2/U1  ( .A(n2667), .B(n1690), .C(in_MUX_inSEL9[1]), .D(
        n2668), .Q(out_MUX_outMUX10[2]) );
  OAI222 \u_mux10/mux1/U1  ( .A(n2665), .B(n1690), .C(in_MUX_inSEL9[1]), .D(
        n2666), .Q(out_MUX_outMUX10[1]) );
  OAI222 \u_mux10/mux0/U1  ( .A(n2663), .B(n1690), .C(in_MUX_inSEL9[1]), .D(
        n2664), .Q(out_MUX_outMUX10[0]) );
  OAI222 \u_mux9/mux3/U1  ( .A(n2661), .B(n1690), .C(in_MUX_inSEL9[1]), .D(
        n2662), .Q(out_MUX_outMUX9[3]) );
  OAI222 \u_mux9/mux2/U1  ( .A(n2659), .B(n1690), .C(in_MUX_inSEL9[1]), .D(
        n2660), .Q(out_MUX_outMUX9[2]) );
  OAI222 \u_mux9/mux1/U1  ( .A(n2657), .B(n1690), .C(in_MUX_inSEL9[1]), .D(
        n2658), .Q(out_MUX_outMUX9[1]) );
  OAI222 \u_mux9/mux0/U1  ( .A(n2655), .B(n1690), .C(in_MUX_inSEL9[1]), .D(
        n2656), .Q(out_MUX_outMUX9[0]) );
  OAI222 \u_mux16/U1  ( .A(n2653), .B(n1694), .C(in_MUX_inSEL15[1]), .D(n2654), 
        .Q(out_MUX_outMUX16) );
  OAI222 \u_mux15/U1  ( .A(n2651), .B(n1694), .C(in_MUX_inSEL15[1]), .D(n2652), 
        .Q(out_MUX_outMUX15) );
  ADD22 \u_cdr/phd1/cnt_phd/add_65/U1_1_1  ( .A(\u_cdr/phd1/cnt_phd/cnt [1]), 
        .B(\u_cdr/phd1/cnt_phd/cnt [0]), .CO(
        \u_cdr/phd1/cnt_phd/add_65/carry [2]), .S(\u_cdr/phd1/cnt_phd/N80 ) );
  ADD22 \u_cdr/phd1/cnt_phd/add_65/U1_1_2  ( .A(\u_cdr/phd1/cnt_phd/cnt [2]), 
        .B(\u_cdr/phd1/cnt_phd/add_65/carry [2]), .CO(
        \u_cdr/phd1/cnt_phd/add_65/carry [3]), .S(\u_cdr/phd1/cnt_phd/N81 ) );
  ADD22 \u_cdr/phd1/cnt_phd/add_65/U1_1_3  ( .A(\u_cdr/phd1/cnt_phd/cnt [3]), 
        .B(\u_cdr/phd1/cnt_phd/add_65/carry [3]), .CO(
        \u_cdr/phd1/cnt_phd/add_65/carry [4]), .S(\u_cdr/phd1/cnt_phd/N82 ) );
  ADD22 \u_cdr/phd1/cnt_phd/add_65/U1_1_4  ( .A(\u_cdr/phd1/cnt_phd/cnt [4]), 
        .B(\u_cdr/phd1/cnt_phd/add_65/carry [4]), .CO(
        \u_cdr/phd1/cnt_phd/add_65/carry [5]), .S(\u_cdr/phd1/cnt_phd/N83 ) );
  ADD22 \u_cdr/dec1/cnt_dec/add_65/U1_1_1  ( .A(\u_cdr/dec1/cnt_dec/cnt [1]), 
        .B(\u_cdr/dec1/cnt_dec/cnt [0]), .CO(
        \u_cdr/dec1/cnt_dec/add_65/carry [2]), .S(\u_cdr/dec1/cnt_dec/N80 ) );
  ADD22 \u_cdr/dec1/cnt_dec/add_65/U1_1_2  ( .A(\u_cdr/dec1/cnt_dec/cnt [2]), 
        .B(\u_cdr/dec1/cnt_dec/add_65/carry [2]), .CO(
        \u_cdr/dec1/cnt_dec/add_65/carry [3]), .S(\u_cdr/dec1/cnt_dec/N81 ) );
  ADD22 \u_cdr/dec1/cnt_dec/add_65/U1_1_3  ( .A(\u_cdr/dec1/cnt_dec/cnt [3]), 
        .B(\u_cdr/dec1/cnt_dec/add_65/carry [3]), .CO(
        \u_cdr/dec1/cnt_dec/add_65/carry [4]), .S(\u_cdr/dec1/cnt_dec/N82 ) );
  ADD22 \u_cdr/dec1/cnt_dec/add_65/U1_1_4  ( .A(\u_cdr/dec1/cnt_dec/cnt [4]), 
        .B(\u_cdr/dec1/cnt_dec/add_65/carry [4]), .CO(
        \u_cdr/dec1/cnt_dec/add_65/carry [5]), .S(\u_cdr/dec1/cnt_dec/N83 ) );
  ADD22 \u_cdr/div1/cnt_div/add_65/U1_1_1  ( .A(\u_cdr/div1/cnt_div/cnt [1]), 
        .B(\u_cdr/div1/cnt_div/cnt [0]), .CO(
        \u_cdr/div1/cnt_div/add_65/carry [2]), .S(\u_cdr/div1/cnt_div/N80 ) );
  ADD22 \u_cdr/div1/cnt_div/add_65/U1_1_2  ( .A(\u_cdr/div1/cnt_div/cnt [2]), 
        .B(\u_cdr/div1/cnt_div/add_65/carry [2]), .CO(
        \u_cdr/div1/cnt_div/add_65/carry [3]), .S(\u_cdr/div1/cnt_div/N81 ) );
  ADD22 \u_cdr/div1/cnt_div/add_65/U1_1_3  ( .A(\u_cdr/div1/cnt_div/cnt [3]), 
        .B(\u_cdr/div1/cnt_div/add_65/carry [3]), .CO(
        \u_cdr/div1/cnt_div/add_65/carry [4]), .S(\u_cdr/div1/cnt_div/N82 ) );
  ADD22 \u_cdr/div1/cnt_div/add_65/U1_1_4  ( .A(\u_cdr/div1/cnt_div/cnt [4]), 
        .B(\u_cdr/div1/cnt_div/add_65/carry [4]), .CO(
        \u_cdr/div1/cnt_div/add_65/carry [5]), .S(\u_cdr/div1/cnt_div/N83 ) );
  ADD22 \u_cdr/dec1/add_41/U1_1_1  ( .A(\u_cdr/dec1/cnt_r [1]), .B(
        \u_cdr/dec1/cnt_r [0]), .CO(\u_cdr/dec1/add_41/carry [2]), .S(
        \u_cdr/dec1/N61 ) );
  ADD22 \u_cdr/dec1/add_41/U1_1_2  ( .A(\u_cdr/dec1/cnt_r [2]), .B(
        \u_cdr/dec1/add_41/carry [2]), .CO(\u_cdr/dec1/add_41/carry [3]), .S(
        \u_cdr/dec1/N62 ) );
  ADD22 \u_cdr/dec1/add_41/U1_1_3  ( .A(\u_cdr/dec1/cnt_r [3]), .B(
        \u_cdr/dec1/add_41/carry [3]), .CO(\u_cdr/dec1/add_41/carry [4]), .S(
        \u_cdr/dec1/N63 ) );
  ADD22 \u_cdr/dec1/add_41/U1_1_4  ( .A(\u_cdr/dec1/cnt_r [4]), .B(
        \u_cdr/dec1/add_41/carry [4]), .CO(\u_cdr/dec1/add_41/carry [5]), .S(
        \u_cdr/dec1/N64 ) );
  ADD32 \u_cordic/my_rotation/sub_40/U2_1  ( .A(
        \u_cordic/my_rotation/present_angle[0][1] ), .B(n68), .CI(
        \u_cordic/my_rotation/sub_40/carry [1]), .CO(
        \u_cordic/my_rotation/sub_40/carry [2]), .S(
        \u_cordic/my_rotation/next_delta [1]) );
  ADD32 \u_cordic/my_rotation/sub_40/U2_2  ( .A(
        \u_cordic/my_rotation/present_angle[0][2] ), .B(n111), .CI(
        \u_cordic/my_rotation/sub_40/carry [2]), .CO(
        \u_cordic/my_rotation/sub_40/carry [3]), .S(
        \u_cordic/my_rotation/next_delta [2]) );
  ADD32 \u_cordic/my_rotation/sub_40/U2_3  ( .A(
        \u_cordic/my_rotation/present_angle[0][3] ), .B(n110), .CI(
        \u_cordic/my_rotation/sub_40/carry [3]), .CO(
        \u_cordic/my_rotation/sub_40/carry [4]), .S(
        \u_cordic/my_rotation/next_delta [3]) );
  ADD32 \u_cordic/my_rotation/sub_40/U2_4  ( .A(
        \u_cordic/my_rotation/present_angle[0][4] ), .B(n127), .CI(
        \u_cordic/my_rotation/sub_40/carry [4]), .CO(
        \u_cordic/my_rotation/sub_40/carry [5]), .S(
        \u_cordic/my_rotation/next_delta [4]) );
  ADD32 \u_cordic/my_rotation/sub_40/U2_5  ( .A(
        \u_cordic/my_rotation/present_angle[0][5] ), .B(n141), .CI(
        \u_cordic/my_rotation/sub_40/carry [5]), .CO(
        \u_cordic/my_rotation/sub_40/carry [6]), .S(
        \u_cordic/my_rotation/next_delta [5]) );
  ADD32 \u_cordic/my_rotation/sub_40/U2_6  ( .A(
        \u_cordic/my_rotation/present_angle[0][6] ), .B(n140), .CI(
        \u_cordic/my_rotation/sub_40/carry [6]), .CO(
        \u_cordic/my_rotation/sub_40/carry [7]), .S(
        \u_cordic/my_rotation/next_delta [6]) );
  ADD32 \u_cordic/my_rotation/sub_40/U2_7  ( .A(
        \u_cordic/my_rotation/present_angle[0][7] ), .B(n163), .CI(
        \u_cordic/my_rotation/sub_40/carry [7]), .CO(
        \u_cordic/my_rotation/sub_40/carry [8]), .S(
        \u_cordic/my_rotation/next_delta [7]) );
  ADD32 \u_cordic/my_rotation/sub_40/U2_8  ( .A(
        \u_cordic/my_rotation/present_angle[0][8] ), .B(n195), .CI(
        \u_cordic/my_rotation/sub_40/carry [8]), .CO(
        \u_cordic/my_rotation/sub_40/carry [9]), .S(
        \u_cordic/my_rotation/next_delta [8]) );
  ADD32 \u_cordic/my_rotation/sub_40/U2_9  ( .A(
        \u_cordic/my_rotation/present_angle[0][9] ), .B(n194), .CI(
        \u_cordic/my_rotation/sub_40/carry [9]), .CO(
        \u_cordic/my_rotation/sub_40/carry [10]), .S(
        \u_cordic/my_rotation/next_delta [9]) );
  ADD32 \u_cordic/my_rotation/sub_40/U2_10  ( .A(
        \u_cordic/my_rotation/present_angle[0][10] ), .B(n228), .CI(
        \u_cordic/my_rotation/sub_40/carry [10]), .CO(
        \u_cordic/my_rotation/sub_40/carry [11]), .S(
        \u_cordic/my_rotation/next_delta [10]) );
  ADD32 \u_cordic/my_rotation/sub_40/U2_11  ( .A(
        \u_cordic/my_rotation/present_angle[0][11] ), .B(n256), .CI(
        \u_cordic/my_rotation/sub_40/carry [11]), .CO(
        \u_cordic/my_rotation/sub_40/carry [12]), .S(
        \u_cordic/my_rotation/next_delta [11]) );
  ADD32 \u_cordic/my_rotation/sub_40/U2_12  ( .A(
        \u_cordic/my_rotation/present_angle[0][12] ), .B(n255), .CI(
        \u_cordic/my_rotation/sub_40/carry [12]), .CO(
        \u_cordic/my_rotation/sub_40/carry [13]), .S(
        \u_cordic/my_rotation/next_delta [12]) );
  ADD32 \u_cordic/my_rotation/sub_40/U2_13  ( .A(
        \u_cordic/my_rotation/present_angle[0][13] ), .B(n275), .CI(
        \u_cordic/my_rotation/sub_40/carry [13]), .CO(
        \u_cordic/my_rotation/sub_40/carry [14]), .S(
        \u_cordic/my_rotation/next_delta [13]) );
  ADD32 \u_cordic/my_rotation/sub_40/U2_14  ( .A(
        \u_cordic/my_rotation/present_angle[0][14] ), .B(n296), .CI(
        \u_cordic/my_rotation/sub_40/carry [14]), .CO(
        \u_cordic/my_rotation/sub_40/carry [15]), .S(
        \u_cordic/my_rotation/next_delta [14]) );
  ADD32 \u_cordic/mycordic/r144/U1_4  ( .A(
        \u_cordic/mycordic/present_I_table[1][4] ), .B(
        \u_cordic/mycordic/present_Q_table[1][4] ), .CI(
        \u_cordic/mycordic/r144/carry [4]), .CO(
        \u_cordic/mycordic/r144/carry [5]), .S(\u_cordic/mycordic/N256 ) );
  ADD32 \u_cordic/mycordic/r144/U1_5  ( .A(
        \u_cordic/mycordic/present_I_table[1][5] ), .B(
        \u_cordic/mycordic/present_Q_table[1][5] ), .CI(
        \u_cordic/mycordic/r144/carry [5]), .CO(
        \u_cordic/mycordic/r144/carry [6]), .S(\u_cordic/mycordic/N257 ) );
  ADD32 \u_cordic/mycordic/r144/U1_6  ( .A(
        \u_cordic/mycordic/present_I_table[1][6] ), .B(
        \u_cordic/mycordic/present_Q_table[1][6] ), .CI(
        \u_cordic/mycordic/r144/carry [6]), .CO(
        \u_cordic/mycordic/r144/carry [7]), .S(\u_cordic/mycordic/N258 ) );
  ADD32 \u_cordic/mycordic/r144/U1_7  ( .A(
        \u_cordic/mycordic/present_I_table[1][7] ), .B(
        \u_cordic/mycordic/present_Q_table[1][7] ), .CI(
        \u_cordic/mycordic/r144/carry [7]), .S(\u_cordic/mycordic/N259 ) );
  ADD32 \u_cordic/mycordic/sub_178/U2_4  ( .A(
        \u_cordic/mycordic/present_Q_table[1][4] ), .B(n251), .CI(
        \u_cordic/mycordic/sub_178/carry [4]), .CO(
        \u_cordic/mycordic/sub_178/carry [5]), .S(\u_cordic/mycordic/N264 ) );
  ADD32 \u_cordic/mycordic/sub_178/U2_5  ( .A(
        \u_cordic/mycordic/present_Q_table[1][5] ), .B(n273), .CI(
        \u_cordic/mycordic/sub_178/carry [5]), .CO(
        \u_cordic/mycordic/sub_178/carry [6]), .S(\u_cordic/mycordic/N265 ) );
  ADD32 \u_cordic/mycordic/sub_178/U2_6  ( .A(
        \u_cordic/mycordic/present_Q_table[1][6] ), .B(n272), .CI(
        \u_cordic/mycordic/sub_178/carry [6]), .CO(
        \u_cordic/mycordic/sub_178/carry [7]), .S(\u_cordic/mycordic/N266 ) );
  ADD32 \u_cordic/mycordic/sub_182/U2_4  ( .A(
        \u_cordic/mycordic/present_I_table[1][4] ), .B(n253), .CI(
        \u_cordic/mycordic/sub_182/carry [4]), .CO(
        \u_cordic/mycordic/sub_182/carry [5]), .S(\u_cordic/mycordic/N288 ) );
  ADD32 \u_cordic/mycordic/sub_182/U2_5  ( .A(
        \u_cordic/mycordic/present_I_table[1][5] ), .B(n252), .CI(
        \u_cordic/mycordic/sub_182/carry [5]), .CO(
        \u_cordic/mycordic/sub_182/carry [6]), .S(\u_cordic/mycordic/N289 ) );
  ADD32 \u_cordic/mycordic/sub_182/U2_6  ( .A(
        \u_cordic/mycordic/present_I_table[1][6] ), .B(n274), .CI(
        \u_cordic/mycordic/sub_182/carry [6]), .CO(
        \u_cordic/mycordic/sub_182/carry [7]), .S(\u_cordic/mycordic/N290 ) );
  ADD32 \u_cordic/mycordic/add_189/U1_1  ( .A(
        \u_cordic/mycordic/present_I_table[2][1] ), .B(
        \u_cordic/mycordic/present_Q_table[2][2] ), .CI(
        \u_cordic/mycordic/add_189/carry [1]), .CO(
        \u_cordic/mycordic/add_189/carry [2]), .S(\u_cordic/mycordic/N317 ) );
  ADD32 \u_cordic/mycordic/add_189/U1_2  ( .A(
        \u_cordic/mycordic/present_I_table[2][2] ), .B(
        \u_cordic/mycordic/present_Q_table[2][3] ), .CI(
        \u_cordic/mycordic/add_189/carry [2]), .CO(
        \u_cordic/mycordic/add_189/carry [3]), .S(\u_cordic/mycordic/N318 ) );
  ADD32 \u_cordic/mycordic/add_189/U1_3  ( .A(
        \u_cordic/mycordic/present_I_table[2][3] ), .B(
        \u_cordic/mycordic/present_Q_table[2][4] ), .CI(
        \u_cordic/mycordic/add_189/carry [3]), .CO(
        \u_cordic/mycordic/add_189/carry [4]), .S(\u_cordic/mycordic/N319 ) );
  ADD32 \u_cordic/mycordic/add_189/U1_4  ( .A(
        \u_cordic/mycordic/present_I_table[2][4] ), .B(
        \u_cordic/mycordic/present_Q_table[2][5] ), .CI(
        \u_cordic/mycordic/add_189/carry [4]), .CO(
        \u_cordic/mycordic/add_189/carry [5]), .S(\u_cordic/mycordic/N320 ) );
  ADD32 \u_cordic/mycordic/add_189/U1_5  ( .A(
        \u_cordic/mycordic/present_I_table[2][5] ), .B(
        \u_cordic/mycordic/present_Q_table[2][6] ), .CI(
        \u_cordic/mycordic/add_189/carry [5]), .CO(
        \u_cordic/mycordic/add_189/carry [6]), .S(\u_cordic/mycordic/N321 ) );
  ADD32 \u_cordic/mycordic/add_189/U1_6  ( .A(
        \u_cordic/mycordic/present_I_table[2][6] ), .B(
        \u_cordic/mycordic/present_Q_table[2][7] ), .CI(
        \u_cordic/mycordic/add_189/carry [6]), .CO(
        \u_cordic/mycordic/add_189/carry [7]), .S(\u_cordic/mycordic/N322 ) );
  ADD32 \u_cordic/mycordic/sub_190/U2_1  ( .A(
        \u_cordic/mycordic/present_Q_table[2][1] ), .B(n192), .CI(
        \u_cordic/mycordic/sub_190/carry [1]), .CO(
        \u_cordic/mycordic/sub_190/carry [2]), .S(\u_cordic/mycordic/N325 ) );
  ADD32 \u_cordic/mycordic/sub_190/U2_2  ( .A(
        \u_cordic/mycordic/present_Q_table[2][2] ), .B(n191), .CI(
        \u_cordic/mycordic/sub_190/carry [2]), .CO(
        \u_cordic/mycordic/sub_190/carry [3]), .S(\u_cordic/mycordic/N326 ) );
  ADD32 \u_cordic/mycordic/sub_190/U2_3  ( .A(
        \u_cordic/mycordic/present_Q_table[2][3] ), .B(n222), .CI(
        \u_cordic/mycordic/sub_190/carry [3]), .CO(
        \u_cordic/mycordic/sub_190/carry [4]), .S(\u_cordic/mycordic/N327 ) );
  ADD32 \u_cordic/mycordic/sub_190/U2_4  ( .A(
        \u_cordic/mycordic/present_Q_table[2][4] ), .B(n249), .CI(
        \u_cordic/mycordic/sub_190/carry [4]), .CO(
        \u_cordic/mycordic/sub_190/carry [5]), .S(\u_cordic/mycordic/N328 ) );
  ADD32 \u_cordic/mycordic/sub_190/U2_5  ( .A(
        \u_cordic/mycordic/present_Q_table[2][5] ), .B(n248), .CI(
        \u_cordic/mycordic/sub_190/carry [5]), .CO(
        \u_cordic/mycordic/sub_190/carry [6]), .S(\u_cordic/mycordic/N329 ) );
  ADD32 \u_cordic/mycordic/sub_190/U2_6  ( .A(
        \u_cordic/mycordic/present_Q_table[2][6] ), .B(n270), .CI(
        \u_cordic/mycordic/sub_190/carry [6]), .CO(
        \u_cordic/mycordic/sub_190/carry [7]), .S(\u_cordic/mycordic/N330 ) );
  ADD32 \u_cordic/mycordic/sub_194/U2_1  ( .A(
        \u_cordic/mycordic/present_I_table[2][1] ), .B(n190), .CI(
        \u_cordic/mycordic/sub_194/carry [1]), .CO(
        \u_cordic/mycordic/sub_194/carry [2]), .S(\u_cordic/mycordic/N349 ) );
  ADD32 \u_cordic/mycordic/sub_194/U2_2  ( .A(
        \u_cordic/mycordic/present_I_table[2][2] ), .B(n189), .CI(
        \u_cordic/mycordic/sub_194/carry [2]), .CO(
        \u_cordic/mycordic/sub_194/carry [3]), .S(\u_cordic/mycordic/N350 ) );
  ADD32 \u_cordic/mycordic/sub_194/U2_3  ( .A(
        \u_cordic/mycordic/present_I_table[2][3] ), .B(n221), .CI(
        \u_cordic/mycordic/sub_194/carry [3]), .CO(
        \u_cordic/mycordic/sub_194/carry [4]), .S(\u_cordic/mycordic/N351 ) );
  ADD32 \u_cordic/mycordic/sub_194/U2_4  ( .A(
        \u_cordic/mycordic/present_I_table[2][4] ), .B(n247), .CI(
        \u_cordic/mycordic/sub_194/carry [4]), .CO(
        \u_cordic/mycordic/sub_194/carry [5]), .S(\u_cordic/mycordic/N352 ) );
  ADD32 \u_cordic/mycordic/sub_194/U2_5  ( .A(
        \u_cordic/mycordic/present_I_table[2][5] ), .B(n246), .CI(
        \u_cordic/mycordic/sub_194/carry [5]), .CO(
        \u_cordic/mycordic/sub_194/carry [6]), .S(\u_cordic/mycordic/N353 ) );
  ADD32 \u_cordic/mycordic/sub_194/U2_6  ( .A(
        \u_cordic/mycordic/present_I_table[2][6] ), .B(n268), .CI(
        \u_cordic/mycordic/sub_194/carry [6]), .CO(
        \u_cordic/mycordic/sub_194/carry [7]), .S(\u_cordic/mycordic/N354 ) );
  ADD32 \u_cordic/mycordic/add_195/U1_1  ( .A(
        \u_cordic/mycordic/present_Q_table[2][1] ), .B(
        \u_cordic/mycordic/present_I_table[2][2] ), .CI(
        \u_cordic/mycordic/add_195/carry [1]), .CO(
        \u_cordic/mycordic/add_195/carry [2]), .S(\u_cordic/mycordic/N357 ) );
  ADD32 \u_cordic/mycordic/add_195/U1_2  ( .A(
        \u_cordic/mycordic/present_Q_table[2][2] ), .B(
        \u_cordic/mycordic/present_I_table[2][3] ), .CI(
        \u_cordic/mycordic/add_195/carry [2]), .CO(
        \u_cordic/mycordic/add_195/carry [3]), .S(\u_cordic/mycordic/N358 ) );
  ADD32 \u_cordic/mycordic/add_195/U1_3  ( .A(
        \u_cordic/mycordic/present_Q_table[2][3] ), .B(
        \u_cordic/mycordic/present_I_table[2][4] ), .CI(
        \u_cordic/mycordic/add_195/carry [3]), .CO(
        \u_cordic/mycordic/add_195/carry [4]), .S(\u_cordic/mycordic/N359 ) );
  ADD32 \u_cordic/mycordic/add_195/U1_4  ( .A(
        \u_cordic/mycordic/present_Q_table[2][4] ), .B(
        \u_cordic/mycordic/present_I_table[2][5] ), .CI(
        \u_cordic/mycordic/add_195/carry [4]), .CO(
        \u_cordic/mycordic/add_195/carry [5]), .S(\u_cordic/mycordic/N360 ) );
  ADD32 \u_cordic/mycordic/add_195/U1_5  ( .A(
        \u_cordic/mycordic/present_Q_table[2][5] ), .B(
        \u_cordic/mycordic/present_I_table[2][6] ), .CI(
        \u_cordic/mycordic/add_195/carry [5]), .CO(
        \u_cordic/mycordic/add_195/carry [6]), .S(\u_cordic/mycordic/N361 ) );
  ADD32 \u_cordic/mycordic/add_195/U1_6  ( .A(
        \u_cordic/mycordic/present_Q_table[2][6] ), .B(
        \u_cordic/mycordic/present_I_table[2][7] ), .CI(
        \u_cordic/mycordic/add_195/carry [6]), .CO(
        \u_cordic/mycordic/add_195/carry [7]), .S(\u_cordic/mycordic/N362 ) );
  ADD32 \u_cordic/mycordic/add_200/U1_1  ( .A(
        \u_cordic/mycordic/present_I_table[3][1] ), .B(
        \u_cordic/mycordic/present_Q_table[3][3] ), .CI(
        \u_cordic/mycordic/add_200/carry [1]), .CO(
        \u_cordic/mycordic/add_200/carry [2]), .S(\u_cordic/mycordic/N381 ) );
  ADD32 \u_cordic/mycordic/add_200/U1_2  ( .A(
        \u_cordic/mycordic/present_I_table[3][2] ), .B(
        \u_cordic/mycordic/present_Q_table[3][4] ), .CI(
        \u_cordic/mycordic/add_200/carry [2]), .CO(
        \u_cordic/mycordic/add_200/carry [3]), .S(\u_cordic/mycordic/N382 ) );
  ADD32 \u_cordic/mycordic/add_200/U1_3  ( .A(
        \u_cordic/mycordic/present_I_table[3][3] ), .B(
        \u_cordic/mycordic/present_Q_table[3][5] ), .CI(
        \u_cordic/mycordic/add_200/carry [3]), .CO(
        \u_cordic/mycordic/add_200/carry [4]), .S(\u_cordic/mycordic/N383 ) );
  ADD32 \u_cordic/mycordic/add_200/U1_4  ( .A(
        \u_cordic/mycordic/present_I_table[3][4] ), .B(
        \u_cordic/mycordic/present_Q_table[3][6] ), .CI(
        \u_cordic/mycordic/add_200/carry [4]), .CO(
        \u_cordic/mycordic/add_200/carry [5]), .S(\u_cordic/mycordic/N384 ) );
  ADD32 \u_cordic/mycordic/add_200/U1_5  ( .A(
        \u_cordic/mycordic/present_I_table[3][5] ), .B(
        \u_cordic/mycordic/present_Q_table[3][7] ), .CI(
        \u_cordic/mycordic/add_200/carry [5]), .CO(
        \u_cordic/mycordic/add_200/carry [6]), .S(\u_cordic/mycordic/N385 ) );
  ADD32 \u_cordic/mycordic/add_200/U1_6  ( .A(
        \u_cordic/mycordic/present_I_table[3][6] ), .B(
        \u_cordic/mycordic/present_Q_table[3][7] ), .CI(
        \u_cordic/mycordic/add_200/carry [6]), .CO(
        \u_cordic/mycordic/add_200/carry [7]), .S(\u_cordic/mycordic/N386 ) );
  ADD32 \u_cordic/mycordic/sub_201/U2_1  ( .A(
        \u_cordic/mycordic/present_Q_table[3][1] ), .B(n188), .CI(
        \u_cordic/mycordic/sub_201/carry [1]), .CO(
        \u_cordic/mycordic/sub_201/carry [2]), .S(\u_cordic/mycordic/N389 ) );
  ADD32 \u_cordic/mycordic/sub_201/U2_2  ( .A(
        \u_cordic/mycordic/present_Q_table[3][2] ), .B(n187), .CI(
        \u_cordic/mycordic/sub_201/carry [2]), .CO(
        \u_cordic/mycordic/sub_201/carry [3]), .S(\u_cordic/mycordic/N390 ) );
  ADD32 \u_cordic/mycordic/sub_201/U2_3  ( .A(
        \u_cordic/mycordic/present_Q_table[3][3] ), .B(n220), .CI(
        \u_cordic/mycordic/sub_201/carry [3]), .CO(
        \u_cordic/mycordic/sub_201/carry [4]), .S(\u_cordic/mycordic/N391 ) );
  ADD32 \u_cordic/mycordic/sub_201/U2_4  ( .A(
        \u_cordic/mycordic/present_Q_table[3][4] ), .B(n245), .CI(
        \u_cordic/mycordic/sub_201/carry [4]), .CO(
        \u_cordic/mycordic/sub_201/carry [5]), .S(\u_cordic/mycordic/N392 ) );
  ADD32 \u_cordic/mycordic/sub_201/U2_5  ( .A(
        \u_cordic/mycordic/present_Q_table[3][5] ), .B(n243), .CI(
        \u_cordic/mycordic/sub_201/carry [5]), .CO(
        \u_cordic/mycordic/sub_201/carry [6]), .S(\u_cordic/mycordic/N393 ) );
  ADD32 \u_cordic/mycordic/sub_201/U2_6  ( .A(
        \u_cordic/mycordic/present_Q_table[3][6] ), .B(n243), .CI(
        \u_cordic/mycordic/sub_201/carry [6]), .CO(
        \u_cordic/mycordic/sub_201/carry [7]), .S(\u_cordic/mycordic/N394 ) );
  ADD32 \u_cordic/mycordic/sub_205/U2_1  ( .A(
        \u_cordic/mycordic/present_I_table[3][1] ), .B(n186), .CI(
        \u_cordic/mycordic/sub_205/carry [1]), .CO(
        \u_cordic/mycordic/sub_205/carry [2]), .S(\u_cordic/mycordic/N413 ) );
  ADD32 \u_cordic/mycordic/sub_205/U2_2  ( .A(
        \u_cordic/mycordic/present_I_table[3][2] ), .B(n185), .CI(
        \u_cordic/mycordic/sub_205/carry [2]), .CO(
        \u_cordic/mycordic/sub_205/carry [3]), .S(\u_cordic/mycordic/N414 ) );
  ADD32 \u_cordic/mycordic/sub_205/U2_3  ( .A(
        \u_cordic/mycordic/present_I_table[3][3] ), .B(n219), .CI(
        \u_cordic/mycordic/sub_205/carry [3]), .CO(
        \u_cordic/mycordic/sub_205/carry [4]), .S(\u_cordic/mycordic/N415 ) );
  ADD32 \u_cordic/mycordic/sub_205/U2_4  ( .A(
        \u_cordic/mycordic/present_I_table[3][4] ), .B(n244), .CI(
        \u_cordic/mycordic/sub_205/carry [4]), .CO(
        \u_cordic/mycordic/sub_205/carry [5]), .S(\u_cordic/mycordic/N416 ) );
  ADD32 \u_cordic/mycordic/sub_205/U2_5  ( .A(
        \u_cordic/mycordic/present_I_table[3][5] ), .B(n242), .CI(
        \u_cordic/mycordic/sub_205/carry [5]), .CO(
        \u_cordic/mycordic/sub_205/carry [6]), .S(\u_cordic/mycordic/N417 ) );
  ADD32 \u_cordic/mycordic/sub_205/U2_6  ( .A(
        \u_cordic/mycordic/present_I_table[3][6] ), .B(n242), .CI(
        \u_cordic/mycordic/sub_205/carry [6]), .CO(
        \u_cordic/mycordic/sub_205/carry [7]), .S(\u_cordic/mycordic/N418 ) );
  ADD32 \u_cordic/mycordic/add_206/U1_1  ( .A(
        \u_cordic/mycordic/present_Q_table[3][1] ), .B(
        \u_cordic/mycordic/present_I_table[3][3] ), .CI(
        \u_cordic/mycordic/add_206/carry [1]), .CO(
        \u_cordic/mycordic/add_206/carry [2]), .S(\u_cordic/mycordic/N421 ) );
  ADD32 \u_cordic/mycordic/add_206/U1_2  ( .A(
        \u_cordic/mycordic/present_Q_table[3][2] ), .B(
        \u_cordic/mycordic/present_I_table[3][4] ), .CI(
        \u_cordic/mycordic/add_206/carry [2]), .CO(
        \u_cordic/mycordic/add_206/carry [3]), .S(\u_cordic/mycordic/N422 ) );
  ADD32 \u_cordic/mycordic/add_206/U1_3  ( .A(
        \u_cordic/mycordic/present_Q_table[3][3] ), .B(
        \u_cordic/mycordic/present_I_table[3][5] ), .CI(
        \u_cordic/mycordic/add_206/carry [3]), .CO(
        \u_cordic/mycordic/add_206/carry [4]), .S(\u_cordic/mycordic/N423 ) );
  ADD32 \u_cordic/mycordic/add_206/U1_4  ( .A(
        \u_cordic/mycordic/present_Q_table[3][4] ), .B(
        \u_cordic/mycordic/present_I_table[3][6] ), .CI(
        \u_cordic/mycordic/add_206/carry [4]), .CO(
        \u_cordic/mycordic/add_206/carry [5]), .S(\u_cordic/mycordic/N424 ) );
  ADD32 \u_cordic/mycordic/add_206/U1_5  ( .A(
        \u_cordic/mycordic/present_Q_table[3][5] ), .B(
        \u_cordic/mycordic/present_I_table[3][7] ), .CI(
        \u_cordic/mycordic/add_206/carry [5]), .CO(
        \u_cordic/mycordic/add_206/carry [6]), .S(\u_cordic/mycordic/N425 ) );
  ADD32 \u_cordic/mycordic/add_206/U1_6  ( .A(
        \u_cordic/mycordic/present_Q_table[3][6] ), .B(
        \u_cordic/mycordic/present_I_table[3][7] ), .CI(
        \u_cordic/mycordic/add_206/carry [6]), .CO(
        \u_cordic/mycordic/add_206/carry [7]), .S(\u_cordic/mycordic/N426 ) );
  ADD32 \u_cordic/mycordic/add_211/U1_4  ( .A(
        \u_cordic/mycordic/present_I_table[4][4] ), .B(n749), .CI(n2217), .CO(
        \u_cordic/mycordic/add_211/carry [5]), .S(\u_cordic/mycordic/N444 ) );
  ADD32 \u_cordic/mycordic/add_211/U1_5  ( .A(
        \u_cordic/mycordic/present_I_table[4][5] ), .B(n749), .CI(
        \u_cordic/mycordic/add_211/carry [5]), .CO(
        \u_cordic/mycordic/add_211/carry [6]), .S(\u_cordic/mycordic/N445 ) );
  ADD32 \u_cordic/mycordic/add_211/U1_6  ( .A(
        \u_cordic/mycordic/present_I_table[4][6] ), .B(n749), .CI(
        \u_cordic/mycordic/add_211/carry [6]), .CO(
        \u_cordic/mycordic/add_211/carry [7]), .S(\u_cordic/mycordic/N446 ) );
  ADD32 \u_cordic/mycordic/sub_212/U2_1  ( .A(
        \u_cordic/mycordic/present_Q_table[4][1] ), .B(n184), .CI(
        \u_cordic/mycordic/sub_212/carry [1]), .CO(
        \u_cordic/mycordic/sub_212/carry [2]), .S(\u_cordic/mycordic/N449 ) );
  ADD32 \u_cordic/mycordic/sub_212/U2_2  ( .A(
        \u_cordic/mycordic/present_Q_table[4][2] ), .B(n183), .CI(
        \u_cordic/mycordic/sub_212/carry [2]), .CO(
        \u_cordic/mycordic/sub_212/carry [3]), .S(\u_cordic/mycordic/N450 ) );
  ADD32 \u_cordic/mycordic/sub_212/U2_3  ( .A(
        \u_cordic/mycordic/present_Q_table[4][3] ), .B(n218), .CI(
        \u_cordic/mycordic/sub_212/carry [3]), .CO(
        \u_cordic/mycordic/sub_212/carry [4]), .S(\u_cordic/mycordic/N451 ) );
  ADD32 \u_cordic/mycordic/sub_212/U2_4  ( .A(
        \u_cordic/mycordic/present_Q_table[4][4] ), .B(n214), .CI(
        \u_cordic/mycordic/sub_212/carry [4]), .CO(
        \u_cordic/mycordic/sub_212/carry [5]), .S(\u_cordic/mycordic/N452 ) );
  ADD32 \u_cordic/mycordic/sub_212/U2_5  ( .A(
        \u_cordic/mycordic/present_Q_table[4][5] ), .B(n214), .CI(
        \u_cordic/mycordic/sub_212/carry [5]), .CO(
        \u_cordic/mycordic/sub_212/carry [6]), .S(\u_cordic/mycordic/N453 ) );
  ADD32 \u_cordic/mycordic/sub_212/U2_6  ( .A(
        \u_cordic/mycordic/present_Q_table[4][6] ), .B(n214), .CI(
        \u_cordic/mycordic/sub_212/carry [6]), .CO(
        \u_cordic/mycordic/sub_212/carry [7]), .S(\u_cordic/mycordic/N454 ) );
  ADD32 \u_cordic/mycordic/sub_216/U2_4  ( .A(
        \u_cordic/mycordic/present_I_table[4][4] ), .B(n180), .CI(
        \u_cordic/mycordic/sub_216/carry [4]), .CO(
        \u_cordic/mycordic/sub_216/carry [5]), .S(\u_cordic/mycordic/N472 ) );
  ADD32 \u_cordic/mycordic/sub_216/U2_5  ( .A(
        \u_cordic/mycordic/present_I_table[4][5] ), .B(n180), .CI(
        \u_cordic/mycordic/sub_216/carry [5]), .CO(
        \u_cordic/mycordic/sub_216/carry [6]), .S(\u_cordic/mycordic/N473 ) );
  ADD32 \u_cordic/mycordic/sub_216/U2_6  ( .A(
        \u_cordic/mycordic/present_I_table[4][6] ), .B(n180), .CI(
        \u_cordic/mycordic/sub_216/carry [6]), .CO(
        \u_cordic/mycordic/sub_216/carry [7]), .S(\u_cordic/mycordic/N474 ) );
  ADD32 \u_cordic/mycordic/add_217/U1_1  ( .A(
        \u_cordic/mycordic/present_Q_table[4][1] ), .B(
        \u_cordic/mycordic/present_I_table[4][4] ), .CI(
        \u_cordic/mycordic/add_217/carry [1]), .CO(
        \u_cordic/mycordic/add_217/carry [2]), .S(\u_cordic/mycordic/N477 ) );
  ADD32 \u_cordic/mycordic/add_217/U1_2  ( .A(
        \u_cordic/mycordic/present_Q_table[4][2] ), .B(
        \u_cordic/mycordic/present_I_table[4][5] ), .CI(
        \u_cordic/mycordic/add_217/carry [2]), .CO(
        \u_cordic/mycordic/add_217/carry [3]), .S(\u_cordic/mycordic/N478 ) );
  ADD32 \u_cordic/mycordic/add_217/U1_3  ( .A(
        \u_cordic/mycordic/present_Q_table[4][3] ), .B(
        \u_cordic/mycordic/present_I_table[4][6] ), .CI(
        \u_cordic/mycordic/add_217/carry [3]), .CO(
        \u_cordic/mycordic/add_217/carry [4]), .S(\u_cordic/mycordic/N479 ) );
  ADD32 \u_cordic/mycordic/add_217/U1_4  ( .A(
        \u_cordic/mycordic/present_Q_table[4][4] ), .B(
        \u_cordic/mycordic/present_I_table[4][7] ), .CI(
        \u_cordic/mycordic/add_217/carry [4]), .CO(
        \u_cordic/mycordic/add_217/carry [5]), .S(\u_cordic/mycordic/N480 ) );
  ADD32 \u_cordic/mycordic/add_217/U1_5  ( .A(
        \u_cordic/mycordic/present_Q_table[4][5] ), .B(
        \u_cordic/mycordic/present_I_table[4][7] ), .CI(
        \u_cordic/mycordic/add_217/carry [5]), .CO(
        \u_cordic/mycordic/add_217/carry [6]), .S(\u_cordic/mycordic/N481 ) );
  ADD32 \u_cordic/mycordic/add_217/U1_6  ( .A(
        \u_cordic/mycordic/present_Q_table[4][6] ), .B(
        \u_cordic/mycordic/present_I_table[4][7] ), .CI(
        \u_cordic/mycordic/add_217/carry [6]), .CO(
        \u_cordic/mycordic/add_217/carry [7]), .S(\u_cordic/mycordic/N482 ) );
  ADD32 \u_decoder/fir_filter/add_294/U1_11  ( .A(
        \u_decoder/fir_filter/I_data_mult_0_buff [11]), .B(
        \u_decoder/fir_filter/I_data_add_1_buff [11]), .CI(
        \u_decoder/fir_filter/add_294/carry [11]), .CO(
        \u_decoder/fir_filter/add_294/carry [12]), .S(
        \u_decoder/fir_filter/I_data_add_0 [11]) );
  ADD32 \u_decoder/fir_filter/add_294/U1_12  ( .A(
        \u_decoder/fir_filter/I_data_mult_0_buff [12]), .B(
        \u_decoder/fir_filter/I_data_add_1_buff [12]), .CI(
        \u_decoder/fir_filter/add_294/carry [12]), .CO(
        \u_decoder/fir_filter/add_294/carry [13]), .S(
        \u_decoder/fir_filter/I_data_add_0 [12]) );
  ADD32 \u_decoder/fir_filter/add_294/U1_13  ( .A(
        \u_decoder/fir_filter/I_data_mult_0_buff [13]), .B(
        \u_decoder/fir_filter/I_data_add_1_buff [13]), .CI(
        \u_decoder/fir_filter/add_294/carry [13]), .CO(
        \u_decoder/fir_filter/add_294/carry [14]), .S(
        \u_decoder/fir_filter/I_data_add_0 [13]) );
  ADD32 \u_decoder/fir_filter/add_295/U1_1  ( .A(
        \u_decoder/fir_filter/I_data_mult_1_buff [1]), .B(
        \u_decoder/fir_filter/I_data_add_2_buff [1]), .CI(
        \u_decoder/fir_filter/add_295/carry [1]), .CO(
        \u_decoder/fir_filter/add_295/carry [2]), .S(
        \u_decoder/fir_filter/I_data_add_1 [1]) );
  ADD32 \u_decoder/fir_filter/add_295/U1_2  ( .A(
        \u_decoder/fir_filter/I_data_mult_1_buff [2]), .B(
        \u_decoder/fir_filter/I_data_add_2_buff [2]), .CI(
        \u_decoder/fir_filter/add_295/carry [2]), .CO(
        \u_decoder/fir_filter/add_295/carry [3]), .S(
        \u_decoder/fir_filter/I_data_add_1 [2]) );
  ADD32 \u_decoder/fir_filter/add_295/U1_3  ( .A(
        \u_decoder/fir_filter/I_data_mult_1_buff [3]), .B(
        \u_decoder/fir_filter/I_data_add_2_buff [3]), .CI(
        \u_decoder/fir_filter/add_295/carry [3]), .CO(
        \u_decoder/fir_filter/add_295/carry [4]), .S(
        \u_decoder/fir_filter/I_data_add_1 [3]) );
  ADD32 \u_decoder/fir_filter/add_295/U1_4  ( .A(
        \u_decoder/fir_filter/I_data_mult_1_buff [4]), .B(
        \u_decoder/fir_filter/I_data_add_2_buff [4]), .CI(
        \u_decoder/fir_filter/add_295/carry [4]), .CO(
        \u_decoder/fir_filter/add_295/carry [5]), .S(
        \u_decoder/fir_filter/I_data_add_1 [4]) );
  ADD32 \u_decoder/fir_filter/add_295/U1_5  ( .A(
        \u_decoder/fir_filter/I_data_mult_1_buff [5]), .B(
        \u_decoder/fir_filter/I_data_add_2_buff [5]), .CI(
        \u_decoder/fir_filter/add_295/carry [5]), .CO(
        \u_decoder/fir_filter/add_295/carry [6]), .S(
        \u_decoder/fir_filter/I_data_add_1 [5]) );
  ADD32 \u_decoder/fir_filter/add_295/U1_6  ( .A(
        \u_decoder/fir_filter/I_data_mult_1_buff [6]), .B(
        \u_decoder/fir_filter/I_data_add_2_buff [6]), .CI(
        \u_decoder/fir_filter/add_295/carry [6]), .CO(
        \u_decoder/fir_filter/add_295/carry [7]), .S(
        \u_decoder/fir_filter/I_data_add_1 [6]) );
  ADD32 \u_decoder/fir_filter/add_295/U1_7  ( .A(
        \u_decoder/fir_filter/I_data_mult_1_buff [7]), .B(
        \u_decoder/fir_filter/I_data_add_2_buff [7]), .CI(
        \u_decoder/fir_filter/add_295/carry [7]), .CO(
        \u_decoder/fir_filter/add_295/carry [8]), .S(
        \u_decoder/fir_filter/I_data_add_1 [7]) );
  ADD32 \u_decoder/fir_filter/add_295/U1_8  ( .A(
        \u_decoder/fir_filter/I_data_mult_1_buff [8]), .B(
        \u_decoder/fir_filter/I_data_add_2_buff [8]), .CI(
        \u_decoder/fir_filter/add_295/carry [8]), .CO(
        \u_decoder/fir_filter/add_295/carry [9]), .S(
        \u_decoder/fir_filter/I_data_add_1 [8]) );
  ADD32 \u_decoder/fir_filter/add_295/U1_9  ( .A(
        \u_decoder/fir_filter/I_data_mult_1_buff [9]), .B(
        \u_decoder/fir_filter/I_data_add_2_buff [9]), .CI(
        \u_decoder/fir_filter/add_295/carry [9]), .CO(
        \u_decoder/fir_filter/add_295/carry [10]), .S(
        \u_decoder/fir_filter/I_data_add_1 [9]) );
  ADD32 \u_decoder/fir_filter/add_295/U1_10  ( .A(
        \u_decoder/fir_filter/I_data_mult_1_buff [10]), .B(
        \u_decoder/fir_filter/I_data_add_2_buff [10]), .CI(
        \u_decoder/fir_filter/add_295/carry [10]), .CO(
        \u_decoder/fir_filter/add_295/carry [11]), .S(
        \u_decoder/fir_filter/I_data_add_1 [10]) );
  ADD32 \u_decoder/fir_filter/add_295/U1_11  ( .A(
        \u_decoder/fir_filter/I_data_mult_1_buff [11]), .B(
        \u_decoder/fir_filter/I_data_add_2_buff [11]), .CI(
        \u_decoder/fir_filter/add_295/carry [11]), .CO(
        \u_decoder/fir_filter/add_295/carry [12]), .S(
        \u_decoder/fir_filter/I_data_add_1 [11]) );
  ADD32 \u_decoder/fir_filter/add_295/U1_12  ( .A(
        \u_decoder/fir_filter/I_data_mult_1_buff [12]), .B(
        \u_decoder/fir_filter/I_data_add_2_buff [12]), .CI(
        \u_decoder/fir_filter/add_295/carry [12]), .CO(
        \u_decoder/fir_filter/add_295/carry [13]), .S(
        \u_decoder/fir_filter/I_data_add_1 [12]) );
  ADD32 \u_decoder/fir_filter/add_295/U1_13  ( .A(
        \u_decoder/fir_filter/I_data_mult_1_buff [13]), .B(
        \u_decoder/fir_filter/I_data_add_2_buff [13]), .CI(
        \u_decoder/fir_filter/add_295/carry [13]), .CO(
        \u_decoder/fir_filter/add_295/carry [14]), .S(
        \u_decoder/fir_filter/I_data_add_1 [13]) );
  ADD32 \u_decoder/fir_filter/add_296/U1_1  ( .A(
        \u_decoder/fir_filter/I_data_mult_2_buff [1]), .B(
        \u_decoder/fir_filter/I_data_add_3_buff [1]), .CI(
        \u_decoder/fir_filter/add_296/carry [1]), .CO(
        \u_decoder/fir_filter/add_296/carry [2]), .S(
        \u_decoder/fir_filter/I_data_add_2 [1]) );
  ADD32 \u_decoder/fir_filter/add_296/U1_2  ( .A(
        \u_decoder/fir_filter/I_data_mult_2_buff [2]), .B(
        \u_decoder/fir_filter/I_data_add_3_buff [2]), .CI(
        \u_decoder/fir_filter/add_296/carry [2]), .CO(
        \u_decoder/fir_filter/add_296/carry [3]), .S(
        \u_decoder/fir_filter/I_data_add_2 [2]) );
  ADD32 \u_decoder/fir_filter/add_296/U1_3  ( .A(
        \u_decoder/fir_filter/I_data_mult_2_buff [3]), .B(
        \u_decoder/fir_filter/I_data_add_3_buff [3]), .CI(
        \u_decoder/fir_filter/add_296/carry [3]), .CO(
        \u_decoder/fir_filter/add_296/carry [4]), .S(
        \u_decoder/fir_filter/I_data_add_2 [3]) );
  ADD32 \u_decoder/fir_filter/add_296/U1_4  ( .A(
        \u_decoder/fir_filter/I_data_mult_2_buff [4]), .B(
        \u_decoder/fir_filter/I_data_add_3_buff [4]), .CI(
        \u_decoder/fir_filter/add_296/carry [4]), .CO(
        \u_decoder/fir_filter/add_296/carry [5]), .S(
        \u_decoder/fir_filter/I_data_add_2 [4]) );
  ADD32 \u_decoder/fir_filter/add_296/U1_5  ( .A(
        \u_decoder/fir_filter/I_data_mult_2_buff [5]), .B(
        \u_decoder/fir_filter/I_data_add_3_buff [5]), .CI(
        \u_decoder/fir_filter/add_296/carry [5]), .CO(
        \u_decoder/fir_filter/add_296/carry [6]), .S(
        \u_decoder/fir_filter/I_data_add_2 [5]) );
  ADD32 \u_decoder/fir_filter/add_296/U1_6  ( .A(
        \u_decoder/fir_filter/I_data_mult_2_buff [6]), .B(
        \u_decoder/fir_filter/I_data_add_3_buff [6]), .CI(
        \u_decoder/fir_filter/add_296/carry [6]), .CO(
        \u_decoder/fir_filter/add_296/carry [7]), .S(
        \u_decoder/fir_filter/I_data_add_2 [6]) );
  ADD32 \u_decoder/fir_filter/add_296/U1_7  ( .A(
        \u_decoder/fir_filter/I_data_mult_2_buff [7]), .B(
        \u_decoder/fir_filter/I_data_add_3_buff [7]), .CI(
        \u_decoder/fir_filter/add_296/carry [7]), .CO(
        \u_decoder/fir_filter/add_296/carry [8]), .S(
        \u_decoder/fir_filter/I_data_add_2 [7]) );
  ADD32 \u_decoder/fir_filter/add_296/U1_8  ( .A(
        \u_decoder/fir_filter/I_data_mult_2_buff [8]), .B(
        \u_decoder/fir_filter/I_data_add_3_buff [8]), .CI(
        \u_decoder/fir_filter/add_296/carry [8]), .CO(
        \u_decoder/fir_filter/add_296/carry [9]), .S(
        \u_decoder/fir_filter/I_data_add_2 [8]) );
  ADD32 \u_decoder/fir_filter/add_296/U1_9  ( .A(
        \u_decoder/fir_filter/I_data_mult_2_buff [9]), .B(
        \u_decoder/fir_filter/I_data_add_3_buff [9]), .CI(
        \u_decoder/fir_filter/add_296/carry [9]), .CO(
        \u_decoder/fir_filter/add_296/carry [10]), .S(
        \u_decoder/fir_filter/I_data_add_2 [9]) );
  ADD32 \u_decoder/fir_filter/add_296/U1_10  ( .A(
        \u_decoder/fir_filter/I_data_mult_2_buff [10]), .B(
        \u_decoder/fir_filter/I_data_add_3_buff [10]), .CI(
        \u_decoder/fir_filter/add_296/carry [10]), .CO(
        \u_decoder/fir_filter/add_296/carry [11]), .S(
        \u_decoder/fir_filter/I_data_add_2 [10]) );
  ADD32 \u_decoder/fir_filter/add_296/U1_11  ( .A(
        \u_decoder/fir_filter/I_data_mult_2_buff [11]), .B(
        \u_decoder/fir_filter/I_data_add_3_buff [11]), .CI(
        \u_decoder/fir_filter/add_296/carry [11]), .CO(
        \u_decoder/fir_filter/add_296/carry [12]), .S(
        \u_decoder/fir_filter/I_data_add_2 [11]) );
  ADD32 \u_decoder/fir_filter/add_296/U1_12  ( .A(
        \u_decoder/fir_filter/I_data_mult_2_buff [12]), .B(
        \u_decoder/fir_filter/I_data_add_3_buff [12]), .CI(
        \u_decoder/fir_filter/add_296/carry [12]), .CO(
        \u_decoder/fir_filter/add_296/carry [13]), .S(
        \u_decoder/fir_filter/I_data_add_2 [12]) );
  ADD32 \u_decoder/fir_filter/add_296/U1_13  ( .A(
        \u_decoder/fir_filter/I_data_mult_2_buff [13]), .B(
        \u_decoder/fir_filter/I_data_add_3_buff [13]), .CI(
        \u_decoder/fir_filter/add_296/carry [13]), .CO(
        \u_decoder/fir_filter/add_296/carry [14]), .S(
        \u_decoder/fir_filter/I_data_add_2 [13]) );
  ADD32 \u_decoder/fir_filter/add_297/U1_1  ( .A(
        \u_decoder/fir_filter/I_data_mult_3_buff [1]), .B(
        \u_decoder/fir_filter/I_data_add_4_buff [1]), .CI(
        \u_decoder/fir_filter/add_297/carry [1]), .CO(
        \u_decoder/fir_filter/add_297/carry [2]), .S(
        \u_decoder/fir_filter/I_data_add_3 [1]) );
  ADD32 \u_decoder/fir_filter/add_297/U1_2  ( .A(
        \u_decoder/fir_filter/I_data_mult_3_buff [2]), .B(
        \u_decoder/fir_filter/I_data_add_4_buff [2]), .CI(
        \u_decoder/fir_filter/add_297/carry [2]), .CO(
        \u_decoder/fir_filter/add_297/carry [3]), .S(
        \u_decoder/fir_filter/I_data_add_3 [2]) );
  ADD32 \u_decoder/fir_filter/add_297/U1_3  ( .A(
        \u_decoder/fir_filter/I_data_mult_3_buff [3]), .B(
        \u_decoder/fir_filter/I_data_add_4_buff [3]), .CI(
        \u_decoder/fir_filter/add_297/carry [3]), .CO(
        \u_decoder/fir_filter/add_297/carry [4]), .S(
        \u_decoder/fir_filter/I_data_add_3 [3]) );
  ADD32 \u_decoder/fir_filter/add_297/U1_4  ( .A(
        \u_decoder/fir_filter/I_data_mult_3_buff [4]), .B(
        \u_decoder/fir_filter/I_data_add_4_buff [4]), .CI(
        \u_decoder/fir_filter/add_297/carry [4]), .CO(
        \u_decoder/fir_filter/add_297/carry [5]), .S(
        \u_decoder/fir_filter/I_data_add_3 [4]) );
  ADD32 \u_decoder/fir_filter/add_297/U1_5  ( .A(
        \u_decoder/fir_filter/I_data_mult_3_buff [5]), .B(
        \u_decoder/fir_filter/I_data_add_4_buff [5]), .CI(
        \u_decoder/fir_filter/add_297/carry [5]), .CO(
        \u_decoder/fir_filter/add_297/carry [6]), .S(
        \u_decoder/fir_filter/I_data_add_3 [5]) );
  ADD32 \u_decoder/fir_filter/add_297/U1_6  ( .A(
        \u_decoder/fir_filter/I_data_mult_3_buff [6]), .B(
        \u_decoder/fir_filter/I_data_add_4_buff [6]), .CI(
        \u_decoder/fir_filter/add_297/carry [6]), .CO(
        \u_decoder/fir_filter/add_297/carry [7]), .S(
        \u_decoder/fir_filter/I_data_add_3 [6]) );
  ADD32 \u_decoder/fir_filter/add_297/U1_7  ( .A(
        \u_decoder/fir_filter/I_data_mult_3_buff [7]), .B(
        \u_decoder/fir_filter/I_data_add_4_buff [7]), .CI(
        \u_decoder/fir_filter/add_297/carry [7]), .CO(
        \u_decoder/fir_filter/add_297/carry [8]), .S(
        \u_decoder/fir_filter/I_data_add_3 [7]) );
  ADD32 \u_decoder/fir_filter/add_297/U1_8  ( .A(
        \u_decoder/fir_filter/I_data_mult_3_buff [8]), .B(
        \u_decoder/fir_filter/I_data_add_4_buff [8]), .CI(
        \u_decoder/fir_filter/add_297/carry [8]), .CO(
        \u_decoder/fir_filter/add_297/carry [9]), .S(
        \u_decoder/fir_filter/I_data_add_3 [8]) );
  ADD32 \u_decoder/fir_filter/add_297/U1_9  ( .A(
        \u_decoder/fir_filter/I_data_mult_3_buff [9]), .B(
        \u_decoder/fir_filter/I_data_add_4_buff [9]), .CI(
        \u_decoder/fir_filter/add_297/carry [9]), .CO(
        \u_decoder/fir_filter/add_297/carry [10]), .S(
        \u_decoder/fir_filter/I_data_add_3 [9]) );
  ADD32 \u_decoder/fir_filter/add_297/U1_10  ( .A(
        \u_decoder/fir_filter/I_data_mult_3_buff [10]), .B(
        \u_decoder/fir_filter/I_data_add_4_buff [10]), .CI(
        \u_decoder/fir_filter/add_297/carry [10]), .CO(
        \u_decoder/fir_filter/add_297/carry [11]), .S(
        \u_decoder/fir_filter/I_data_add_3 [10]) );
  ADD32 \u_decoder/fir_filter/add_297/U1_11  ( .A(
        \u_decoder/fir_filter/I_data_mult_3_buff [11]), .B(
        \u_decoder/fir_filter/I_data_add_4_buff [11]), .CI(
        \u_decoder/fir_filter/add_297/carry [11]), .CO(
        \u_decoder/fir_filter/add_297/carry [12]), .S(
        \u_decoder/fir_filter/I_data_add_3 [11]) );
  ADD32 \u_decoder/fir_filter/add_297/U1_12  ( .A(
        \u_decoder/fir_filter/I_data_mult_3_buff [12]), .B(
        \u_decoder/fir_filter/I_data_add_4_buff [12]), .CI(
        \u_decoder/fir_filter/add_297/carry [12]), .CO(
        \u_decoder/fir_filter/add_297/carry [13]), .S(
        \u_decoder/fir_filter/I_data_add_3 [12]) );
  ADD32 \u_decoder/fir_filter/add_297/U1_13  ( .A(
        \u_decoder/fir_filter/I_data_mult_3_buff [13]), .B(
        \u_decoder/fir_filter/I_data_add_4_buff [13]), .CI(
        \u_decoder/fir_filter/add_297/carry [13]), .CO(
        \u_decoder/fir_filter/add_297/carry [14]), .S(
        \u_decoder/fir_filter/I_data_add_3 [13]) );
  ADD32 \u_decoder/fir_filter/add_298/U1_1  ( .A(
        \u_decoder/fir_filter/I_data_mult_4_buff [1]), .B(
        \u_decoder/fir_filter/I_data_add_5_buff [1]), .CI(
        \u_decoder/fir_filter/add_298/carry [1]), .CO(
        \u_decoder/fir_filter/add_298/carry [2]), .S(
        \u_decoder/fir_filter/I_data_add_4 [1]) );
  ADD32 \u_decoder/fir_filter/add_298/U1_2  ( .A(
        \u_decoder/fir_filter/I_data_mult_4_buff [2]), .B(
        \u_decoder/fir_filter/I_data_add_5_buff [2]), .CI(
        \u_decoder/fir_filter/add_298/carry [2]), .CO(
        \u_decoder/fir_filter/add_298/carry [3]), .S(
        \u_decoder/fir_filter/I_data_add_4 [2]) );
  ADD32 \u_decoder/fir_filter/add_298/U1_3  ( .A(
        \u_decoder/fir_filter/I_data_mult_4_buff [3]), .B(
        \u_decoder/fir_filter/I_data_add_5_buff [3]), .CI(
        \u_decoder/fir_filter/add_298/carry [3]), .CO(
        \u_decoder/fir_filter/add_298/carry [4]), .S(
        \u_decoder/fir_filter/I_data_add_4 [3]) );
  ADD32 \u_decoder/fir_filter/add_298/U1_4  ( .A(
        \u_decoder/fir_filter/I_data_mult_4_buff [4]), .B(
        \u_decoder/fir_filter/I_data_add_5_buff [4]), .CI(
        \u_decoder/fir_filter/add_298/carry [4]), .CO(
        \u_decoder/fir_filter/add_298/carry [5]), .S(
        \u_decoder/fir_filter/I_data_add_4 [4]) );
  ADD32 \u_decoder/fir_filter/add_298/U1_5  ( .A(
        \u_decoder/fir_filter/I_data_mult_4_buff [5]), .B(
        \u_decoder/fir_filter/I_data_add_5_buff [5]), .CI(
        \u_decoder/fir_filter/add_298/carry [5]), .CO(
        \u_decoder/fir_filter/add_298/carry [6]), .S(
        \u_decoder/fir_filter/I_data_add_4 [5]) );
  ADD32 \u_decoder/fir_filter/add_298/U1_6  ( .A(
        \u_decoder/fir_filter/I_data_mult_4_buff [6]), .B(
        \u_decoder/fir_filter/I_data_add_5_buff [6]), .CI(
        \u_decoder/fir_filter/add_298/carry [6]), .CO(
        \u_decoder/fir_filter/add_298/carry [7]), .S(
        \u_decoder/fir_filter/I_data_add_4 [6]) );
  ADD32 \u_decoder/fir_filter/add_298/U1_7  ( .A(
        \u_decoder/fir_filter/I_data_mult_4_buff [7]), .B(
        \u_decoder/fir_filter/I_data_add_5_buff [7]), .CI(
        \u_decoder/fir_filter/add_298/carry [7]), .CO(
        \u_decoder/fir_filter/add_298/carry [8]), .S(
        \u_decoder/fir_filter/I_data_add_4 [7]) );
  ADD32 \u_decoder/fir_filter/add_298/U1_8  ( .A(
        \u_decoder/fir_filter/I_data_mult_4_buff [8]), .B(
        \u_decoder/fir_filter/I_data_add_5_buff [8]), .CI(
        \u_decoder/fir_filter/add_298/carry [8]), .CO(
        \u_decoder/fir_filter/add_298/carry [9]), .S(
        \u_decoder/fir_filter/I_data_add_4 [8]) );
  ADD32 \u_decoder/fir_filter/add_298/U1_9  ( .A(
        \u_decoder/fir_filter/I_data_mult_4_buff [9]), .B(
        \u_decoder/fir_filter/I_data_add_5_buff [9]), .CI(
        \u_decoder/fir_filter/add_298/carry [9]), .CO(
        \u_decoder/fir_filter/add_298/carry [10]), .S(
        \u_decoder/fir_filter/I_data_add_4 [9]) );
  ADD32 \u_decoder/fir_filter/add_298/U1_10  ( .A(
        \u_decoder/fir_filter/I_data_mult_4_buff [10]), .B(
        \u_decoder/fir_filter/I_data_add_5_buff [10]), .CI(
        \u_decoder/fir_filter/add_298/carry [10]), .CO(
        \u_decoder/fir_filter/add_298/carry [11]), .S(
        \u_decoder/fir_filter/I_data_add_4 [10]) );
  ADD32 \u_decoder/fir_filter/add_298/U1_11  ( .A(
        \u_decoder/fir_filter/I_data_mult_4_buff [11]), .B(
        \u_decoder/fir_filter/I_data_add_5_buff [11]), .CI(
        \u_decoder/fir_filter/add_298/carry [11]), .CO(
        \u_decoder/fir_filter/add_298/carry [12]), .S(
        \u_decoder/fir_filter/I_data_add_4 [11]) );
  ADD32 \u_decoder/fir_filter/add_298/U1_12  ( .A(
        \u_decoder/fir_filter/I_data_mult_4_buff [12]), .B(
        \u_decoder/fir_filter/I_data_add_5_buff [12]), .CI(
        \u_decoder/fir_filter/add_298/carry [12]), .CO(
        \u_decoder/fir_filter/add_298/carry [13]), .S(
        \u_decoder/fir_filter/I_data_add_4 [12]) );
  ADD32 \u_decoder/fir_filter/add_298/U1_13  ( .A(
        \u_decoder/fir_filter/I_data_mult_4_buff [13]), .B(
        \u_decoder/fir_filter/I_data_add_5_buff [13]), .CI(
        \u_decoder/fir_filter/add_298/carry [13]), .CO(
        \u_decoder/fir_filter/add_298/carry [14]), .S(
        \u_decoder/fir_filter/I_data_add_4 [13]) );
  ADD32 \u_decoder/fir_filter/add_299/U1_1  ( .A(
        \u_decoder/fir_filter/I_data_mult_5_buff [1]), .B(
        \u_decoder/fir_filter/I_data_add_6_buff [1]), .CI(
        \u_decoder/fir_filter/add_299/carry [1]), .CO(
        \u_decoder/fir_filter/add_299/carry [2]), .S(
        \u_decoder/fir_filter/I_data_add_5 [1]) );
  ADD32 \u_decoder/fir_filter/add_299/U1_2  ( .A(
        \u_decoder/fir_filter/I_data_mult_5_buff [2]), .B(
        \u_decoder/fir_filter/I_data_add_6_buff [2]), .CI(
        \u_decoder/fir_filter/add_299/carry [2]), .CO(
        \u_decoder/fir_filter/add_299/carry [3]), .S(
        \u_decoder/fir_filter/I_data_add_5 [2]) );
  ADD32 \u_decoder/fir_filter/add_299/U1_3  ( .A(
        \u_decoder/fir_filter/I_data_mult_5_buff [3]), .B(
        \u_decoder/fir_filter/I_data_add_6_buff [3]), .CI(
        \u_decoder/fir_filter/add_299/carry [3]), .CO(
        \u_decoder/fir_filter/add_299/carry [4]), .S(
        \u_decoder/fir_filter/I_data_add_5 [3]) );
  ADD32 \u_decoder/fir_filter/add_299/U1_4  ( .A(
        \u_decoder/fir_filter/I_data_mult_5_buff [4]), .B(
        \u_decoder/fir_filter/I_data_add_6_buff [4]), .CI(
        \u_decoder/fir_filter/add_299/carry [4]), .CO(
        \u_decoder/fir_filter/add_299/carry [5]), .S(
        \u_decoder/fir_filter/I_data_add_5 [4]) );
  ADD32 \u_decoder/fir_filter/add_299/U1_5  ( .A(
        \u_decoder/fir_filter/I_data_mult_5_buff [5]), .B(
        \u_decoder/fir_filter/I_data_add_6_buff [5]), .CI(
        \u_decoder/fir_filter/add_299/carry [5]), .CO(
        \u_decoder/fir_filter/add_299/carry [6]), .S(
        \u_decoder/fir_filter/I_data_add_5 [5]) );
  ADD32 \u_decoder/fir_filter/add_299/U1_6  ( .A(
        \u_decoder/fir_filter/I_data_mult_5_buff [6]), .B(
        \u_decoder/fir_filter/I_data_add_6_buff [6]), .CI(
        \u_decoder/fir_filter/add_299/carry [6]), .CO(
        \u_decoder/fir_filter/add_299/carry [7]), .S(
        \u_decoder/fir_filter/I_data_add_5 [6]) );
  ADD32 \u_decoder/fir_filter/add_299/U1_7  ( .A(
        \u_decoder/fir_filter/I_data_mult_5_buff [7]), .B(
        \u_decoder/fir_filter/I_data_add_6_buff [7]), .CI(
        \u_decoder/fir_filter/add_299/carry [7]), .CO(
        \u_decoder/fir_filter/add_299/carry [8]), .S(
        \u_decoder/fir_filter/I_data_add_5 [7]) );
  ADD32 \u_decoder/fir_filter/add_299/U1_8  ( .A(
        \u_decoder/fir_filter/I_data_mult_5_buff [8]), .B(
        \u_decoder/fir_filter/I_data_add_6_buff [8]), .CI(
        \u_decoder/fir_filter/add_299/carry [8]), .CO(
        \u_decoder/fir_filter/add_299/carry [9]), .S(
        \u_decoder/fir_filter/I_data_add_5 [8]) );
  ADD32 \u_decoder/fir_filter/add_299/U1_9  ( .A(
        \u_decoder/fir_filter/I_data_mult_5_buff [9]), .B(
        \u_decoder/fir_filter/I_data_add_6_buff [9]), .CI(
        \u_decoder/fir_filter/add_299/carry [9]), .CO(
        \u_decoder/fir_filter/add_299/carry [10]), .S(
        \u_decoder/fir_filter/I_data_add_5 [9]) );
  ADD32 \u_decoder/fir_filter/add_299/U1_10  ( .A(
        \u_decoder/fir_filter/I_data_mult_5_buff [10]), .B(
        \u_decoder/fir_filter/I_data_add_6_buff [10]), .CI(
        \u_decoder/fir_filter/add_299/carry [10]), .CO(
        \u_decoder/fir_filter/add_299/carry [11]), .S(
        \u_decoder/fir_filter/I_data_add_5 [10]) );
  ADD32 \u_decoder/fir_filter/add_299/U1_11  ( .A(
        \u_decoder/fir_filter/I_data_mult_5_buff [11]), .B(
        \u_decoder/fir_filter/I_data_add_6_buff [11]), .CI(
        \u_decoder/fir_filter/add_299/carry [11]), .CO(
        \u_decoder/fir_filter/add_299/carry [12]), .S(
        \u_decoder/fir_filter/I_data_add_5 [11]) );
  ADD32 \u_decoder/fir_filter/add_299/U1_12  ( .A(
        \u_decoder/fir_filter/I_data_mult_5_buff [12]), .B(
        \u_decoder/fir_filter/I_data_add_6_buff [12]), .CI(
        \u_decoder/fir_filter/add_299/carry [12]), .CO(
        \u_decoder/fir_filter/add_299/carry [13]), .S(
        \u_decoder/fir_filter/I_data_add_5 [12]) );
  ADD32 \u_decoder/fir_filter/add_299/U1_13  ( .A(
        \u_decoder/fir_filter/I_data_mult_5_buff [13]), .B(
        \u_decoder/fir_filter/I_data_add_6_buff [13]), .CI(
        \u_decoder/fir_filter/add_299/carry [13]), .CO(
        \u_decoder/fir_filter/add_299/carry [14]), .S(
        \u_decoder/fir_filter/I_data_add_5 [13]) );
  ADD32 \u_decoder/fir_filter/add_300/U1_1  ( .A(
        \u_decoder/fir_filter/I_data_mult_6_buff [1]), .B(
        \u_decoder/fir_filter/I_data_add_7_buff [1]), .CI(
        \u_decoder/fir_filter/add_300/carry [1]), .CO(
        \u_decoder/fir_filter/add_300/carry [2]), .S(
        \u_decoder/fir_filter/I_data_add_6 [1]) );
  ADD32 \u_decoder/fir_filter/add_300/U1_2  ( .A(
        \u_decoder/fir_filter/I_data_mult_6_buff [2]), .B(
        \u_decoder/fir_filter/I_data_add_7_buff [2]), .CI(
        \u_decoder/fir_filter/add_300/carry [2]), .CO(
        \u_decoder/fir_filter/add_300/carry [3]), .S(
        \u_decoder/fir_filter/I_data_add_6 [2]) );
  ADD32 \u_decoder/fir_filter/add_300/U1_3  ( .A(
        \u_decoder/fir_filter/I_data_mult_6_buff [3]), .B(
        \u_decoder/fir_filter/I_data_add_7_buff [3]), .CI(
        \u_decoder/fir_filter/add_300/carry [3]), .CO(
        \u_decoder/fir_filter/add_300/carry [4]), .S(
        \u_decoder/fir_filter/I_data_add_6 [3]) );
  ADD32 \u_decoder/fir_filter/add_300/U1_4  ( .A(
        \u_decoder/fir_filter/I_data_mult_6_buff [4]), .B(
        \u_decoder/fir_filter/I_data_add_7_buff [4]), .CI(
        \u_decoder/fir_filter/add_300/carry [4]), .CO(
        \u_decoder/fir_filter/add_300/carry [5]), .S(
        \u_decoder/fir_filter/I_data_add_6 [4]) );
  ADD32 \u_decoder/fir_filter/add_300/U1_5  ( .A(
        \u_decoder/fir_filter/I_data_mult_6_buff [5]), .B(
        \u_decoder/fir_filter/I_data_add_7_buff [5]), .CI(
        \u_decoder/fir_filter/add_300/carry [5]), .CO(
        \u_decoder/fir_filter/add_300/carry [6]), .S(
        \u_decoder/fir_filter/I_data_add_6 [5]) );
  ADD32 \u_decoder/fir_filter/add_300/U1_6  ( .A(
        \u_decoder/fir_filter/I_data_mult_6_buff [6]), .B(
        \u_decoder/fir_filter/I_data_add_7_buff [6]), .CI(
        \u_decoder/fir_filter/add_300/carry [6]), .CO(
        \u_decoder/fir_filter/add_300/carry [7]), .S(
        \u_decoder/fir_filter/I_data_add_6 [6]) );
  ADD32 \u_decoder/fir_filter/add_300/U1_7  ( .A(
        \u_decoder/fir_filter/I_data_mult_6_buff [7]), .B(
        \u_decoder/fir_filter/I_data_add_7_buff [7]), .CI(
        \u_decoder/fir_filter/add_300/carry [7]), .CO(
        \u_decoder/fir_filter/add_300/carry [8]), .S(
        \u_decoder/fir_filter/I_data_add_6 [7]) );
  ADD32 \u_decoder/fir_filter/add_300/U1_8  ( .A(
        \u_decoder/fir_filter/I_data_mult_6_buff [8]), .B(
        \u_decoder/fir_filter/I_data_add_7_buff [8]), .CI(
        \u_decoder/fir_filter/add_300/carry [8]), .CO(
        \u_decoder/fir_filter/add_300/carry [9]), .S(
        \u_decoder/fir_filter/I_data_add_6 [8]) );
  ADD32 \u_decoder/fir_filter/add_300/U1_9  ( .A(
        \u_decoder/fir_filter/I_data_mult_6_buff [9]), .B(
        \u_decoder/fir_filter/I_data_add_7_buff [9]), .CI(
        \u_decoder/fir_filter/add_300/carry [9]), .CO(
        \u_decoder/fir_filter/add_300/carry [10]), .S(
        \u_decoder/fir_filter/I_data_add_6 [9]) );
  ADD32 \u_decoder/fir_filter/add_300/U1_10  ( .A(
        \u_decoder/fir_filter/I_data_mult_6_buff [10]), .B(
        \u_decoder/fir_filter/I_data_add_7_buff [10]), .CI(
        \u_decoder/fir_filter/add_300/carry [10]), .CO(
        \u_decoder/fir_filter/add_300/carry [11]), .S(
        \u_decoder/fir_filter/I_data_add_6 [10]) );
  ADD32 \u_decoder/fir_filter/add_300/U1_11  ( .A(
        \u_decoder/fir_filter/I_data_mult_6_buff [11]), .B(
        \u_decoder/fir_filter/I_data_add_7_buff [11]), .CI(
        \u_decoder/fir_filter/add_300/carry [11]), .CO(
        \u_decoder/fir_filter/add_300/carry [12]), .S(
        \u_decoder/fir_filter/I_data_add_6 [11]) );
  ADD32 \u_decoder/fir_filter/add_300/U1_12  ( .A(
        \u_decoder/fir_filter/I_data_mult_6_buff [12]), .B(
        \u_decoder/fir_filter/I_data_add_7_buff [12]), .CI(
        \u_decoder/fir_filter/add_300/carry [12]), .CO(
        \u_decoder/fir_filter/add_300/carry [13]), .S(
        \u_decoder/fir_filter/I_data_add_6 [12]) );
  ADD32 \u_decoder/fir_filter/add_300/U1_13  ( .A(
        \u_decoder/fir_filter/I_data_mult_6_buff [13]), .B(
        \u_decoder/fir_filter/I_data_add_7_buff [13]), .CI(
        \u_decoder/fir_filter/add_300/carry [13]), .CO(
        \u_decoder/fir_filter/add_300/carry [14]), .S(
        \u_decoder/fir_filter/I_data_add_6 [13]) );
  ADD32 \u_decoder/fir_filter/add_301/U1_1  ( .A(
        \u_decoder/fir_filter/I_data_mult_7_buff [1]), .B(
        \u_decoder/fir_filter/I_data_mult_8_buff [1]), .CI(
        \u_decoder/fir_filter/add_301/carry [1]), .CO(
        \u_decoder/fir_filter/add_301/carry [2]), .S(
        \u_decoder/fir_filter/I_data_add_7 [1]) );
  ADD32 \u_decoder/fir_filter/add_301/U1_2  ( .A(
        \u_decoder/fir_filter/I_data_mult_7_buff [2]), .B(
        \u_decoder/fir_filter/I_data_mult_8_buff [2]), .CI(
        \u_decoder/fir_filter/add_301/carry [2]), .CO(
        \u_decoder/fir_filter/add_301/carry [3]), .S(
        \u_decoder/fir_filter/I_data_add_7 [2]) );
  ADD32 \u_decoder/fir_filter/add_301/U1_3  ( .A(
        \u_decoder/fir_filter/I_data_mult_7_buff [3]), .B(
        \u_decoder/fir_filter/I_data_mult_8_buff [3]), .CI(
        \u_decoder/fir_filter/add_301/carry [3]), .CO(
        \u_decoder/fir_filter/add_301/carry [4]), .S(
        \u_decoder/fir_filter/I_data_add_7 [3]) );
  ADD32 \u_decoder/fir_filter/add_301/U1_4  ( .A(
        \u_decoder/fir_filter/I_data_mult_7_buff [4]), .B(
        \u_decoder/fir_filter/I_data_mult_8_buff [4]), .CI(
        \u_decoder/fir_filter/add_301/carry [4]), .CO(
        \u_decoder/fir_filter/add_301/carry [5]), .S(
        \u_decoder/fir_filter/I_data_add_7 [4]) );
  ADD32 \u_decoder/fir_filter/add_301/U1_5  ( .A(
        \u_decoder/fir_filter/I_data_mult_7_buff [5]), .B(
        \u_decoder/fir_filter/I_data_mult_8_buff [5]), .CI(
        \u_decoder/fir_filter/add_301/carry [5]), .CO(
        \u_decoder/fir_filter/add_301/carry [6]), .S(
        \u_decoder/fir_filter/I_data_add_7 [5]) );
  ADD32 \u_decoder/fir_filter/add_301/U1_6  ( .A(
        \u_decoder/fir_filter/I_data_mult_7_buff [6]), .B(
        \u_decoder/fir_filter/I_data_mult_8_buff [6]), .CI(
        \u_decoder/fir_filter/add_301/carry [6]), .CO(
        \u_decoder/fir_filter/add_301/carry [7]), .S(
        \u_decoder/fir_filter/I_data_add_7 [6]) );
  ADD32 \u_decoder/fir_filter/add_301/U1_7  ( .A(
        \u_decoder/fir_filter/I_data_mult_7_buff [7]), .B(
        \u_decoder/fir_filter/I_data_mult_8_buff [7]), .CI(
        \u_decoder/fir_filter/add_301/carry [7]), .CO(
        \u_decoder/fir_filter/add_301/carry [8]), .S(
        \u_decoder/fir_filter/I_data_add_7 [7]) );
  ADD32 \u_decoder/fir_filter/add_301/U1_8  ( .A(
        \u_decoder/fir_filter/I_data_mult_7_buff [8]), .B(
        \u_decoder/fir_filter/I_data_mult_8_buff [8]), .CI(
        \u_decoder/fir_filter/add_301/carry [8]), .CO(
        \u_decoder/fir_filter/add_301/carry [9]), .S(
        \u_decoder/fir_filter/I_data_add_7 [8]) );
  ADD32 \u_decoder/fir_filter/add_301/U1_9  ( .A(
        \u_decoder/fir_filter/I_data_mult_7_buff [9]), .B(
        \u_decoder/fir_filter/I_data_mult_8_buff [9]), .CI(
        \u_decoder/fir_filter/add_301/carry [9]), .CO(
        \u_decoder/fir_filter/add_301/carry [10]), .S(
        \u_decoder/fir_filter/I_data_add_7 [9]) );
  ADD32 \u_decoder/fir_filter/add_301/U1_10  ( .A(
        \u_decoder/fir_filter/I_data_mult_7_buff [10]), .B(
        \u_decoder/fir_filter/I_data_mult_8_buff [10]), .CI(
        \u_decoder/fir_filter/add_301/carry [10]), .CO(
        \u_decoder/fir_filter/add_301/carry [11]), .S(
        \u_decoder/fir_filter/I_data_add_7 [10]) );
  ADD32 \u_decoder/fir_filter/add_301/U1_11  ( .A(
        \u_decoder/fir_filter/I_data_mult_7_buff [11]), .B(
        \u_decoder/fir_filter/I_data_mult_8_buff [11]), .CI(
        \u_decoder/fir_filter/add_301/carry [11]), .CO(
        \u_decoder/fir_filter/add_301/carry [12]), .S(
        \u_decoder/fir_filter/I_data_add_7 [11]) );
  ADD32 \u_decoder/fir_filter/add_301/U1_12  ( .A(
        \u_decoder/fir_filter/I_data_mult_7_buff [12]), .B(
        \u_decoder/fir_filter/I_data_mult_8_buff [12]), .CI(
        \u_decoder/fir_filter/add_301/carry [12]), .CO(
        \u_decoder/fir_filter/add_301/carry [13]), .S(
        \u_decoder/fir_filter/I_data_add_7 [12]) );
  ADD32 \u_decoder/fir_filter/add_301/U1_13  ( .A(
        \u_decoder/fir_filter/I_data_mult_7_buff [13]), .B(
        \u_decoder/fir_filter/I_data_mult_8_buff [13]), .CI(
        \u_decoder/fir_filter/add_301/carry [13]), .CO(
        \u_decoder/fir_filter/add_301/carry [14]), .S(
        \u_decoder/fir_filter/I_data_add_7 [13]) );
  ADD32 \u_decoder/fir_filter/add_326/U1_11  ( .A(
        \u_decoder/fir_filter/Q_data_mult_0_buff [11]), .B(
        \u_decoder/fir_filter/Q_data_add_1_buff [11]), .CI(
        \u_decoder/fir_filter/add_326/carry [11]), .CO(
        \u_decoder/fir_filter/add_326/carry [12]), .S(
        \u_decoder/fir_filter/Q_data_add_0 [11]) );
  ADD32 \u_decoder/fir_filter/add_326/U1_12  ( .A(
        \u_decoder/fir_filter/Q_data_mult_0_buff [12]), .B(
        \u_decoder/fir_filter/Q_data_add_1_buff [12]), .CI(
        \u_decoder/fir_filter/add_326/carry [12]), .CO(
        \u_decoder/fir_filter/add_326/carry [13]), .S(
        \u_decoder/fir_filter/Q_data_add_0 [12]) );
  ADD32 \u_decoder/fir_filter/add_326/U1_13  ( .A(
        \u_decoder/fir_filter/Q_data_mult_0_buff [13]), .B(
        \u_decoder/fir_filter/Q_data_add_1_buff [13]), .CI(
        \u_decoder/fir_filter/add_326/carry [13]), .CO(
        \u_decoder/fir_filter/add_326/carry [14]), .S(
        \u_decoder/fir_filter/Q_data_add_0 [13]) );
  ADD32 \u_decoder/fir_filter/add_327/U1_1  ( .A(
        \u_decoder/fir_filter/Q_data_mult_1_buff [1]), .B(
        \u_decoder/fir_filter/Q_data_add_2_buff [1]), .CI(
        \u_decoder/fir_filter/add_327/carry [1]), .CO(
        \u_decoder/fir_filter/add_327/carry [2]), .S(
        \u_decoder/fir_filter/Q_data_add_1 [1]) );
  ADD32 \u_decoder/fir_filter/add_327/U1_2  ( .A(
        \u_decoder/fir_filter/Q_data_mult_1_buff [2]), .B(
        \u_decoder/fir_filter/Q_data_add_2_buff [2]), .CI(
        \u_decoder/fir_filter/add_327/carry [2]), .CO(
        \u_decoder/fir_filter/add_327/carry [3]), .S(
        \u_decoder/fir_filter/Q_data_add_1 [2]) );
  ADD32 \u_decoder/fir_filter/add_327/U1_3  ( .A(
        \u_decoder/fir_filter/Q_data_mult_1_buff [3]), .B(
        \u_decoder/fir_filter/Q_data_add_2_buff [3]), .CI(
        \u_decoder/fir_filter/add_327/carry [3]), .CO(
        \u_decoder/fir_filter/add_327/carry [4]), .S(
        \u_decoder/fir_filter/Q_data_add_1 [3]) );
  ADD32 \u_decoder/fir_filter/add_327/U1_4  ( .A(
        \u_decoder/fir_filter/Q_data_mult_1_buff [4]), .B(
        \u_decoder/fir_filter/Q_data_add_2_buff [4]), .CI(
        \u_decoder/fir_filter/add_327/carry [4]), .CO(
        \u_decoder/fir_filter/add_327/carry [5]), .S(
        \u_decoder/fir_filter/Q_data_add_1 [4]) );
  ADD32 \u_decoder/fir_filter/add_327/U1_5  ( .A(
        \u_decoder/fir_filter/Q_data_mult_1_buff [5]), .B(
        \u_decoder/fir_filter/Q_data_add_2_buff [5]), .CI(
        \u_decoder/fir_filter/add_327/carry [5]), .CO(
        \u_decoder/fir_filter/add_327/carry [6]), .S(
        \u_decoder/fir_filter/Q_data_add_1 [5]) );
  ADD32 \u_decoder/fir_filter/add_327/U1_6  ( .A(
        \u_decoder/fir_filter/Q_data_mult_1_buff [6]), .B(
        \u_decoder/fir_filter/Q_data_add_2_buff [6]), .CI(
        \u_decoder/fir_filter/add_327/carry [6]), .CO(
        \u_decoder/fir_filter/add_327/carry [7]), .S(
        \u_decoder/fir_filter/Q_data_add_1 [6]) );
  ADD32 \u_decoder/fir_filter/add_327/U1_7  ( .A(
        \u_decoder/fir_filter/Q_data_mult_1_buff [7]), .B(
        \u_decoder/fir_filter/Q_data_add_2_buff [7]), .CI(
        \u_decoder/fir_filter/add_327/carry [7]), .CO(
        \u_decoder/fir_filter/add_327/carry [8]), .S(
        \u_decoder/fir_filter/Q_data_add_1 [7]) );
  ADD32 \u_decoder/fir_filter/add_327/U1_8  ( .A(
        \u_decoder/fir_filter/Q_data_mult_1_buff [8]), .B(
        \u_decoder/fir_filter/Q_data_add_2_buff [8]), .CI(
        \u_decoder/fir_filter/add_327/carry [8]), .CO(
        \u_decoder/fir_filter/add_327/carry [9]), .S(
        \u_decoder/fir_filter/Q_data_add_1 [8]) );
  ADD32 \u_decoder/fir_filter/add_327/U1_9  ( .A(
        \u_decoder/fir_filter/Q_data_mult_1_buff [9]), .B(
        \u_decoder/fir_filter/Q_data_add_2_buff [9]), .CI(
        \u_decoder/fir_filter/add_327/carry [9]), .CO(
        \u_decoder/fir_filter/add_327/carry [10]), .S(
        \u_decoder/fir_filter/Q_data_add_1 [9]) );
  ADD32 \u_decoder/fir_filter/add_327/U1_10  ( .A(
        \u_decoder/fir_filter/Q_data_mult_1_buff [10]), .B(
        \u_decoder/fir_filter/Q_data_add_2_buff [10]), .CI(
        \u_decoder/fir_filter/add_327/carry [10]), .CO(
        \u_decoder/fir_filter/add_327/carry [11]), .S(
        \u_decoder/fir_filter/Q_data_add_1 [10]) );
  ADD32 \u_decoder/fir_filter/add_327/U1_11  ( .A(
        \u_decoder/fir_filter/Q_data_mult_1_buff [11]), .B(
        \u_decoder/fir_filter/Q_data_add_2_buff [11]), .CI(
        \u_decoder/fir_filter/add_327/carry [11]), .CO(
        \u_decoder/fir_filter/add_327/carry [12]), .S(
        \u_decoder/fir_filter/Q_data_add_1 [11]) );
  ADD32 \u_decoder/fir_filter/add_327/U1_12  ( .A(
        \u_decoder/fir_filter/Q_data_mult_1_buff [12]), .B(
        \u_decoder/fir_filter/Q_data_add_2_buff [12]), .CI(
        \u_decoder/fir_filter/add_327/carry [12]), .CO(
        \u_decoder/fir_filter/add_327/carry [13]), .S(
        \u_decoder/fir_filter/Q_data_add_1 [12]) );
  ADD32 \u_decoder/fir_filter/add_327/U1_13  ( .A(
        \u_decoder/fir_filter/Q_data_mult_1_buff [13]), .B(
        \u_decoder/fir_filter/Q_data_add_2_buff [13]), .CI(
        \u_decoder/fir_filter/add_327/carry [13]), .CO(
        \u_decoder/fir_filter/add_327/carry [14]), .S(
        \u_decoder/fir_filter/Q_data_add_1 [13]) );
  ADD32 \u_decoder/fir_filter/add_328/U1_1  ( .A(
        \u_decoder/fir_filter/Q_data_mult_2_buff [1]), .B(
        \u_decoder/fir_filter/Q_data_add_3_buff [1]), .CI(
        \u_decoder/fir_filter/add_328/carry [1]), .CO(
        \u_decoder/fir_filter/add_328/carry [2]), .S(
        \u_decoder/fir_filter/Q_data_add_2 [1]) );
  ADD32 \u_decoder/fir_filter/add_328/U1_2  ( .A(
        \u_decoder/fir_filter/Q_data_mult_2_buff [2]), .B(
        \u_decoder/fir_filter/Q_data_add_3_buff [2]), .CI(
        \u_decoder/fir_filter/add_328/carry [2]), .CO(
        \u_decoder/fir_filter/add_328/carry [3]), .S(
        \u_decoder/fir_filter/Q_data_add_2 [2]) );
  ADD32 \u_decoder/fir_filter/add_328/U1_3  ( .A(
        \u_decoder/fir_filter/Q_data_mult_2_buff [3]), .B(
        \u_decoder/fir_filter/Q_data_add_3_buff [3]), .CI(
        \u_decoder/fir_filter/add_328/carry [3]), .CO(
        \u_decoder/fir_filter/add_328/carry [4]), .S(
        \u_decoder/fir_filter/Q_data_add_2 [3]) );
  ADD32 \u_decoder/fir_filter/add_328/U1_4  ( .A(
        \u_decoder/fir_filter/Q_data_mult_2_buff [4]), .B(
        \u_decoder/fir_filter/Q_data_add_3_buff [4]), .CI(
        \u_decoder/fir_filter/add_328/carry [4]), .CO(
        \u_decoder/fir_filter/add_328/carry [5]), .S(
        \u_decoder/fir_filter/Q_data_add_2 [4]) );
  ADD32 \u_decoder/fir_filter/add_328/U1_5  ( .A(
        \u_decoder/fir_filter/Q_data_mult_2_buff [5]), .B(
        \u_decoder/fir_filter/Q_data_add_3_buff [5]), .CI(
        \u_decoder/fir_filter/add_328/carry [5]), .CO(
        \u_decoder/fir_filter/add_328/carry [6]), .S(
        \u_decoder/fir_filter/Q_data_add_2 [5]) );
  ADD32 \u_decoder/fir_filter/add_328/U1_6  ( .A(
        \u_decoder/fir_filter/Q_data_mult_2_buff [6]), .B(
        \u_decoder/fir_filter/Q_data_add_3_buff [6]), .CI(
        \u_decoder/fir_filter/add_328/carry [6]), .CO(
        \u_decoder/fir_filter/add_328/carry [7]), .S(
        \u_decoder/fir_filter/Q_data_add_2 [6]) );
  ADD32 \u_decoder/fir_filter/add_328/U1_7  ( .A(
        \u_decoder/fir_filter/Q_data_mult_2_buff [7]), .B(
        \u_decoder/fir_filter/Q_data_add_3_buff [7]), .CI(
        \u_decoder/fir_filter/add_328/carry [7]), .CO(
        \u_decoder/fir_filter/add_328/carry [8]), .S(
        \u_decoder/fir_filter/Q_data_add_2 [7]) );
  ADD32 \u_decoder/fir_filter/add_328/U1_8  ( .A(
        \u_decoder/fir_filter/Q_data_mult_2_buff [8]), .B(
        \u_decoder/fir_filter/Q_data_add_3_buff [8]), .CI(
        \u_decoder/fir_filter/add_328/carry [8]), .CO(
        \u_decoder/fir_filter/add_328/carry [9]), .S(
        \u_decoder/fir_filter/Q_data_add_2 [8]) );
  ADD32 \u_decoder/fir_filter/add_328/U1_9  ( .A(
        \u_decoder/fir_filter/Q_data_mult_2_buff [9]), .B(
        \u_decoder/fir_filter/Q_data_add_3_buff [9]), .CI(
        \u_decoder/fir_filter/add_328/carry [9]), .CO(
        \u_decoder/fir_filter/add_328/carry [10]), .S(
        \u_decoder/fir_filter/Q_data_add_2 [9]) );
  ADD32 \u_decoder/fir_filter/add_328/U1_10  ( .A(
        \u_decoder/fir_filter/Q_data_mult_2_buff [10]), .B(
        \u_decoder/fir_filter/Q_data_add_3_buff [10]), .CI(
        \u_decoder/fir_filter/add_328/carry [10]), .CO(
        \u_decoder/fir_filter/add_328/carry [11]), .S(
        \u_decoder/fir_filter/Q_data_add_2 [10]) );
  ADD32 \u_decoder/fir_filter/add_328/U1_11  ( .A(
        \u_decoder/fir_filter/Q_data_mult_2_buff [11]), .B(
        \u_decoder/fir_filter/Q_data_add_3_buff [11]), .CI(
        \u_decoder/fir_filter/add_328/carry [11]), .CO(
        \u_decoder/fir_filter/add_328/carry [12]), .S(
        \u_decoder/fir_filter/Q_data_add_2 [11]) );
  ADD32 \u_decoder/fir_filter/add_328/U1_12  ( .A(
        \u_decoder/fir_filter/Q_data_mult_2_buff [12]), .B(
        \u_decoder/fir_filter/Q_data_add_3_buff [12]), .CI(
        \u_decoder/fir_filter/add_328/carry [12]), .CO(
        \u_decoder/fir_filter/add_328/carry [13]), .S(
        \u_decoder/fir_filter/Q_data_add_2 [12]) );
  ADD32 \u_decoder/fir_filter/add_328/U1_13  ( .A(
        \u_decoder/fir_filter/Q_data_mult_2_buff [13]), .B(
        \u_decoder/fir_filter/Q_data_add_3_buff [13]), .CI(
        \u_decoder/fir_filter/add_328/carry [13]), .CO(
        \u_decoder/fir_filter/add_328/carry [14]), .S(
        \u_decoder/fir_filter/Q_data_add_2 [13]) );
  ADD32 \u_decoder/fir_filter/add_329/U1_1  ( .A(
        \u_decoder/fir_filter/Q_data_mult_3_buff [1]), .B(
        \u_decoder/fir_filter/Q_data_add_4_buff [1]), .CI(
        \u_decoder/fir_filter/add_329/carry [1]), .CO(
        \u_decoder/fir_filter/add_329/carry [2]), .S(
        \u_decoder/fir_filter/Q_data_add_3 [1]) );
  ADD32 \u_decoder/fir_filter/add_329/U1_2  ( .A(
        \u_decoder/fir_filter/Q_data_mult_3_buff [2]), .B(
        \u_decoder/fir_filter/Q_data_add_4_buff [2]), .CI(
        \u_decoder/fir_filter/add_329/carry [2]), .CO(
        \u_decoder/fir_filter/add_329/carry [3]), .S(
        \u_decoder/fir_filter/Q_data_add_3 [2]) );
  ADD32 \u_decoder/fir_filter/add_329/U1_3  ( .A(
        \u_decoder/fir_filter/Q_data_mult_3_buff [3]), .B(
        \u_decoder/fir_filter/Q_data_add_4_buff [3]), .CI(
        \u_decoder/fir_filter/add_329/carry [3]), .CO(
        \u_decoder/fir_filter/add_329/carry [4]), .S(
        \u_decoder/fir_filter/Q_data_add_3 [3]) );
  ADD32 \u_decoder/fir_filter/add_329/U1_4  ( .A(
        \u_decoder/fir_filter/Q_data_mult_3_buff [4]), .B(
        \u_decoder/fir_filter/Q_data_add_4_buff [4]), .CI(
        \u_decoder/fir_filter/add_329/carry [4]), .CO(
        \u_decoder/fir_filter/add_329/carry [5]), .S(
        \u_decoder/fir_filter/Q_data_add_3 [4]) );
  ADD32 \u_decoder/fir_filter/add_329/U1_5  ( .A(
        \u_decoder/fir_filter/Q_data_mult_3_buff [5]), .B(
        \u_decoder/fir_filter/Q_data_add_4_buff [5]), .CI(
        \u_decoder/fir_filter/add_329/carry [5]), .CO(
        \u_decoder/fir_filter/add_329/carry [6]), .S(
        \u_decoder/fir_filter/Q_data_add_3 [5]) );
  ADD32 \u_decoder/fir_filter/add_329/U1_6  ( .A(
        \u_decoder/fir_filter/Q_data_mult_3_buff [6]), .B(
        \u_decoder/fir_filter/Q_data_add_4_buff [6]), .CI(
        \u_decoder/fir_filter/add_329/carry [6]), .CO(
        \u_decoder/fir_filter/add_329/carry [7]), .S(
        \u_decoder/fir_filter/Q_data_add_3 [6]) );
  ADD32 \u_decoder/fir_filter/add_329/U1_7  ( .A(
        \u_decoder/fir_filter/Q_data_mult_3_buff [7]), .B(
        \u_decoder/fir_filter/Q_data_add_4_buff [7]), .CI(
        \u_decoder/fir_filter/add_329/carry [7]), .CO(
        \u_decoder/fir_filter/add_329/carry [8]), .S(
        \u_decoder/fir_filter/Q_data_add_3 [7]) );
  ADD32 \u_decoder/fir_filter/add_329/U1_8  ( .A(
        \u_decoder/fir_filter/Q_data_mult_3_buff [8]), .B(
        \u_decoder/fir_filter/Q_data_add_4_buff [8]), .CI(
        \u_decoder/fir_filter/add_329/carry [8]), .CO(
        \u_decoder/fir_filter/add_329/carry [9]), .S(
        \u_decoder/fir_filter/Q_data_add_3 [8]) );
  ADD32 \u_decoder/fir_filter/add_329/U1_9  ( .A(
        \u_decoder/fir_filter/Q_data_mult_3_buff [9]), .B(
        \u_decoder/fir_filter/Q_data_add_4_buff [9]), .CI(
        \u_decoder/fir_filter/add_329/carry [9]), .CO(
        \u_decoder/fir_filter/add_329/carry [10]), .S(
        \u_decoder/fir_filter/Q_data_add_3 [9]) );
  ADD32 \u_decoder/fir_filter/add_329/U1_10  ( .A(
        \u_decoder/fir_filter/Q_data_mult_3_buff [10]), .B(
        \u_decoder/fir_filter/Q_data_add_4_buff [10]), .CI(
        \u_decoder/fir_filter/add_329/carry [10]), .CO(
        \u_decoder/fir_filter/add_329/carry [11]), .S(
        \u_decoder/fir_filter/Q_data_add_3 [10]) );
  ADD32 \u_decoder/fir_filter/add_329/U1_11  ( .A(
        \u_decoder/fir_filter/Q_data_mult_3_buff [11]), .B(
        \u_decoder/fir_filter/Q_data_add_4_buff [11]), .CI(
        \u_decoder/fir_filter/add_329/carry [11]), .CO(
        \u_decoder/fir_filter/add_329/carry [12]), .S(
        \u_decoder/fir_filter/Q_data_add_3 [11]) );
  ADD32 \u_decoder/fir_filter/add_329/U1_12  ( .A(
        \u_decoder/fir_filter/Q_data_mult_3_buff [12]), .B(
        \u_decoder/fir_filter/Q_data_add_4_buff [12]), .CI(
        \u_decoder/fir_filter/add_329/carry [12]), .CO(
        \u_decoder/fir_filter/add_329/carry [13]), .S(
        \u_decoder/fir_filter/Q_data_add_3 [12]) );
  ADD32 \u_decoder/fir_filter/add_329/U1_13  ( .A(
        \u_decoder/fir_filter/Q_data_mult_3_buff [13]), .B(
        \u_decoder/fir_filter/Q_data_add_4_buff [13]), .CI(
        \u_decoder/fir_filter/add_329/carry [13]), .CO(
        \u_decoder/fir_filter/add_329/carry [14]), .S(
        \u_decoder/fir_filter/Q_data_add_3 [13]) );
  ADD32 \u_decoder/fir_filter/add_330/U1_1  ( .A(
        \u_decoder/fir_filter/Q_data_mult_4_buff [1]), .B(
        \u_decoder/fir_filter/Q_data_add_5_buff [1]), .CI(
        \u_decoder/fir_filter/add_330/carry [1]), .CO(
        \u_decoder/fir_filter/add_330/carry [2]), .S(
        \u_decoder/fir_filter/Q_data_add_4 [1]) );
  ADD32 \u_decoder/fir_filter/add_330/U1_2  ( .A(
        \u_decoder/fir_filter/Q_data_mult_4_buff [2]), .B(
        \u_decoder/fir_filter/Q_data_add_5_buff [2]), .CI(
        \u_decoder/fir_filter/add_330/carry [2]), .CO(
        \u_decoder/fir_filter/add_330/carry [3]), .S(
        \u_decoder/fir_filter/Q_data_add_4 [2]) );
  ADD32 \u_decoder/fir_filter/add_330/U1_3  ( .A(
        \u_decoder/fir_filter/Q_data_mult_4_buff [3]), .B(
        \u_decoder/fir_filter/Q_data_add_5_buff [3]), .CI(
        \u_decoder/fir_filter/add_330/carry [3]), .CO(
        \u_decoder/fir_filter/add_330/carry [4]), .S(
        \u_decoder/fir_filter/Q_data_add_4 [3]) );
  ADD32 \u_decoder/fir_filter/add_330/U1_4  ( .A(
        \u_decoder/fir_filter/Q_data_mult_4_buff [4]), .B(
        \u_decoder/fir_filter/Q_data_add_5_buff [4]), .CI(
        \u_decoder/fir_filter/add_330/carry [4]), .CO(
        \u_decoder/fir_filter/add_330/carry [5]), .S(
        \u_decoder/fir_filter/Q_data_add_4 [4]) );
  ADD32 \u_decoder/fir_filter/add_330/U1_5  ( .A(
        \u_decoder/fir_filter/Q_data_mult_4_buff [5]), .B(
        \u_decoder/fir_filter/Q_data_add_5_buff [5]), .CI(
        \u_decoder/fir_filter/add_330/carry [5]), .CO(
        \u_decoder/fir_filter/add_330/carry [6]), .S(
        \u_decoder/fir_filter/Q_data_add_4 [5]) );
  ADD32 \u_decoder/fir_filter/add_330/U1_6  ( .A(
        \u_decoder/fir_filter/Q_data_mult_4_buff [6]), .B(
        \u_decoder/fir_filter/Q_data_add_5_buff [6]), .CI(
        \u_decoder/fir_filter/add_330/carry [6]), .CO(
        \u_decoder/fir_filter/add_330/carry [7]), .S(
        \u_decoder/fir_filter/Q_data_add_4 [6]) );
  ADD32 \u_decoder/fir_filter/add_330/U1_7  ( .A(
        \u_decoder/fir_filter/Q_data_mult_4_buff [7]), .B(
        \u_decoder/fir_filter/Q_data_add_5_buff [7]), .CI(
        \u_decoder/fir_filter/add_330/carry [7]), .CO(
        \u_decoder/fir_filter/add_330/carry [8]), .S(
        \u_decoder/fir_filter/Q_data_add_4 [7]) );
  ADD32 \u_decoder/fir_filter/add_330/U1_8  ( .A(
        \u_decoder/fir_filter/Q_data_mult_4_buff [8]), .B(
        \u_decoder/fir_filter/Q_data_add_5_buff [8]), .CI(
        \u_decoder/fir_filter/add_330/carry [8]), .CO(
        \u_decoder/fir_filter/add_330/carry [9]), .S(
        \u_decoder/fir_filter/Q_data_add_4 [8]) );
  ADD32 \u_decoder/fir_filter/add_330/U1_9  ( .A(
        \u_decoder/fir_filter/Q_data_mult_4_buff [9]), .B(
        \u_decoder/fir_filter/Q_data_add_5_buff [9]), .CI(
        \u_decoder/fir_filter/add_330/carry [9]), .CO(
        \u_decoder/fir_filter/add_330/carry [10]), .S(
        \u_decoder/fir_filter/Q_data_add_4 [9]) );
  ADD32 \u_decoder/fir_filter/add_330/U1_10  ( .A(
        \u_decoder/fir_filter/Q_data_mult_4_buff [10]), .B(
        \u_decoder/fir_filter/Q_data_add_5_buff [10]), .CI(
        \u_decoder/fir_filter/add_330/carry [10]), .CO(
        \u_decoder/fir_filter/add_330/carry [11]), .S(
        \u_decoder/fir_filter/Q_data_add_4 [10]) );
  ADD32 \u_decoder/fir_filter/add_330/U1_11  ( .A(
        \u_decoder/fir_filter/Q_data_mult_4_buff [11]), .B(
        \u_decoder/fir_filter/Q_data_add_5_buff [11]), .CI(
        \u_decoder/fir_filter/add_330/carry [11]), .CO(
        \u_decoder/fir_filter/add_330/carry [12]), .S(
        \u_decoder/fir_filter/Q_data_add_4 [11]) );
  ADD32 \u_decoder/fir_filter/add_330/U1_12  ( .A(
        \u_decoder/fir_filter/Q_data_mult_4_buff [12]), .B(
        \u_decoder/fir_filter/Q_data_add_5_buff [12]), .CI(
        \u_decoder/fir_filter/add_330/carry [12]), .CO(
        \u_decoder/fir_filter/add_330/carry [13]), .S(
        \u_decoder/fir_filter/Q_data_add_4 [12]) );
  ADD32 \u_decoder/fir_filter/add_330/U1_13  ( .A(
        \u_decoder/fir_filter/Q_data_mult_4_buff [13]), .B(
        \u_decoder/fir_filter/Q_data_add_5_buff [13]), .CI(
        \u_decoder/fir_filter/add_330/carry [13]), .CO(
        \u_decoder/fir_filter/add_330/carry [14]), .S(
        \u_decoder/fir_filter/Q_data_add_4 [13]) );
  ADD32 \u_decoder/fir_filter/add_331/U1_1  ( .A(
        \u_decoder/fir_filter/Q_data_mult_5_buff [1]), .B(
        \u_decoder/fir_filter/Q_data_add_6_buff [1]), .CI(
        \u_decoder/fir_filter/add_331/carry [1]), .CO(
        \u_decoder/fir_filter/add_331/carry [2]), .S(
        \u_decoder/fir_filter/Q_data_add_5 [1]) );
  ADD32 \u_decoder/fir_filter/add_331/U1_2  ( .A(
        \u_decoder/fir_filter/Q_data_mult_5_buff [2]), .B(
        \u_decoder/fir_filter/Q_data_add_6_buff [2]), .CI(
        \u_decoder/fir_filter/add_331/carry [2]), .CO(
        \u_decoder/fir_filter/add_331/carry [3]), .S(
        \u_decoder/fir_filter/Q_data_add_5 [2]) );
  ADD32 \u_decoder/fir_filter/add_331/U1_3  ( .A(
        \u_decoder/fir_filter/Q_data_mult_5_buff [3]), .B(
        \u_decoder/fir_filter/Q_data_add_6_buff [3]), .CI(
        \u_decoder/fir_filter/add_331/carry [3]), .CO(
        \u_decoder/fir_filter/add_331/carry [4]), .S(
        \u_decoder/fir_filter/Q_data_add_5 [3]) );
  ADD32 \u_decoder/fir_filter/add_331/U1_4  ( .A(
        \u_decoder/fir_filter/Q_data_mult_5_buff [4]), .B(
        \u_decoder/fir_filter/Q_data_add_6_buff [4]), .CI(
        \u_decoder/fir_filter/add_331/carry [4]), .CO(
        \u_decoder/fir_filter/add_331/carry [5]), .S(
        \u_decoder/fir_filter/Q_data_add_5 [4]) );
  ADD32 \u_decoder/fir_filter/add_331/U1_5  ( .A(
        \u_decoder/fir_filter/Q_data_mult_5_buff [5]), .B(
        \u_decoder/fir_filter/Q_data_add_6_buff [5]), .CI(
        \u_decoder/fir_filter/add_331/carry [5]), .CO(
        \u_decoder/fir_filter/add_331/carry [6]), .S(
        \u_decoder/fir_filter/Q_data_add_5 [5]) );
  ADD32 \u_decoder/fir_filter/add_331/U1_6  ( .A(
        \u_decoder/fir_filter/Q_data_mult_5_buff [6]), .B(
        \u_decoder/fir_filter/Q_data_add_6_buff [6]), .CI(
        \u_decoder/fir_filter/add_331/carry [6]), .CO(
        \u_decoder/fir_filter/add_331/carry [7]), .S(
        \u_decoder/fir_filter/Q_data_add_5 [6]) );
  ADD32 \u_decoder/fir_filter/add_331/U1_7  ( .A(
        \u_decoder/fir_filter/Q_data_mult_5_buff [7]), .B(
        \u_decoder/fir_filter/Q_data_add_6_buff [7]), .CI(
        \u_decoder/fir_filter/add_331/carry [7]), .CO(
        \u_decoder/fir_filter/add_331/carry [8]), .S(
        \u_decoder/fir_filter/Q_data_add_5 [7]) );
  ADD32 \u_decoder/fir_filter/add_331/U1_8  ( .A(
        \u_decoder/fir_filter/Q_data_mult_5_buff [8]), .B(
        \u_decoder/fir_filter/Q_data_add_6_buff [8]), .CI(
        \u_decoder/fir_filter/add_331/carry [8]), .CO(
        \u_decoder/fir_filter/add_331/carry [9]), .S(
        \u_decoder/fir_filter/Q_data_add_5 [8]) );
  ADD32 \u_decoder/fir_filter/add_331/U1_9  ( .A(
        \u_decoder/fir_filter/Q_data_mult_5_buff [9]), .B(
        \u_decoder/fir_filter/Q_data_add_6_buff [9]), .CI(
        \u_decoder/fir_filter/add_331/carry [9]), .CO(
        \u_decoder/fir_filter/add_331/carry [10]), .S(
        \u_decoder/fir_filter/Q_data_add_5 [9]) );
  ADD32 \u_decoder/fir_filter/add_331/U1_10  ( .A(
        \u_decoder/fir_filter/Q_data_mult_5_buff [10]), .B(
        \u_decoder/fir_filter/Q_data_add_6_buff [10]), .CI(
        \u_decoder/fir_filter/add_331/carry [10]), .CO(
        \u_decoder/fir_filter/add_331/carry [11]), .S(
        \u_decoder/fir_filter/Q_data_add_5 [10]) );
  ADD32 \u_decoder/fir_filter/add_331/U1_11  ( .A(
        \u_decoder/fir_filter/Q_data_mult_5_buff [11]), .B(
        \u_decoder/fir_filter/Q_data_add_6_buff [11]), .CI(
        \u_decoder/fir_filter/add_331/carry [11]), .CO(
        \u_decoder/fir_filter/add_331/carry [12]), .S(
        \u_decoder/fir_filter/Q_data_add_5 [11]) );
  ADD32 \u_decoder/fir_filter/add_331/U1_12  ( .A(
        \u_decoder/fir_filter/Q_data_mult_5_buff [12]), .B(
        \u_decoder/fir_filter/Q_data_add_6_buff [12]), .CI(
        \u_decoder/fir_filter/add_331/carry [12]), .CO(
        \u_decoder/fir_filter/add_331/carry [13]), .S(
        \u_decoder/fir_filter/Q_data_add_5 [12]) );
  ADD32 \u_decoder/fir_filter/add_331/U1_13  ( .A(
        \u_decoder/fir_filter/Q_data_mult_5_buff [13]), .B(
        \u_decoder/fir_filter/Q_data_add_6_buff [13]), .CI(
        \u_decoder/fir_filter/add_331/carry [13]), .CO(
        \u_decoder/fir_filter/add_331/carry [14]), .S(
        \u_decoder/fir_filter/Q_data_add_5 [13]) );
  ADD32 \u_decoder/fir_filter/add_332/U1_1  ( .A(
        \u_decoder/fir_filter/Q_data_mult_6_buff [1]), .B(
        \u_decoder/fir_filter/Q_data_add_7_buff [1]), .CI(
        \u_decoder/fir_filter/add_332/carry [1]), .CO(
        \u_decoder/fir_filter/add_332/carry [2]), .S(
        \u_decoder/fir_filter/Q_data_add_6 [1]) );
  ADD32 \u_decoder/fir_filter/add_332/U1_2  ( .A(
        \u_decoder/fir_filter/Q_data_mult_6_buff [2]), .B(
        \u_decoder/fir_filter/Q_data_add_7_buff [2]), .CI(
        \u_decoder/fir_filter/add_332/carry [2]), .CO(
        \u_decoder/fir_filter/add_332/carry [3]), .S(
        \u_decoder/fir_filter/Q_data_add_6 [2]) );
  ADD32 \u_decoder/fir_filter/add_332/U1_3  ( .A(
        \u_decoder/fir_filter/Q_data_mult_6_buff [3]), .B(
        \u_decoder/fir_filter/Q_data_add_7_buff [3]), .CI(
        \u_decoder/fir_filter/add_332/carry [3]), .CO(
        \u_decoder/fir_filter/add_332/carry [4]), .S(
        \u_decoder/fir_filter/Q_data_add_6 [3]) );
  ADD32 \u_decoder/fir_filter/add_332/U1_4  ( .A(
        \u_decoder/fir_filter/Q_data_mult_6_buff [4]), .B(
        \u_decoder/fir_filter/Q_data_add_7_buff [4]), .CI(
        \u_decoder/fir_filter/add_332/carry [4]), .CO(
        \u_decoder/fir_filter/add_332/carry [5]), .S(
        \u_decoder/fir_filter/Q_data_add_6 [4]) );
  ADD32 \u_decoder/fir_filter/add_332/U1_5  ( .A(
        \u_decoder/fir_filter/Q_data_mult_6_buff [5]), .B(
        \u_decoder/fir_filter/Q_data_add_7_buff [5]), .CI(
        \u_decoder/fir_filter/add_332/carry [5]), .CO(
        \u_decoder/fir_filter/add_332/carry [6]), .S(
        \u_decoder/fir_filter/Q_data_add_6 [5]) );
  ADD32 \u_decoder/fir_filter/add_332/U1_6  ( .A(
        \u_decoder/fir_filter/Q_data_mult_6_buff [6]), .B(
        \u_decoder/fir_filter/Q_data_add_7_buff [6]), .CI(
        \u_decoder/fir_filter/add_332/carry [6]), .CO(
        \u_decoder/fir_filter/add_332/carry [7]), .S(
        \u_decoder/fir_filter/Q_data_add_6 [6]) );
  ADD32 \u_decoder/fir_filter/add_332/U1_7  ( .A(
        \u_decoder/fir_filter/Q_data_mult_6_buff [7]), .B(
        \u_decoder/fir_filter/Q_data_add_7_buff [7]), .CI(
        \u_decoder/fir_filter/add_332/carry [7]), .CO(
        \u_decoder/fir_filter/add_332/carry [8]), .S(
        \u_decoder/fir_filter/Q_data_add_6 [7]) );
  ADD32 \u_decoder/fir_filter/add_332/U1_8  ( .A(
        \u_decoder/fir_filter/Q_data_mult_6_buff [8]), .B(
        \u_decoder/fir_filter/Q_data_add_7_buff [8]), .CI(
        \u_decoder/fir_filter/add_332/carry [8]), .CO(
        \u_decoder/fir_filter/add_332/carry [9]), .S(
        \u_decoder/fir_filter/Q_data_add_6 [8]) );
  ADD32 \u_decoder/fir_filter/add_332/U1_9  ( .A(
        \u_decoder/fir_filter/Q_data_mult_6_buff [9]), .B(
        \u_decoder/fir_filter/Q_data_add_7_buff [9]), .CI(
        \u_decoder/fir_filter/add_332/carry [9]), .CO(
        \u_decoder/fir_filter/add_332/carry [10]), .S(
        \u_decoder/fir_filter/Q_data_add_6 [9]) );
  ADD32 \u_decoder/fir_filter/add_332/U1_10  ( .A(
        \u_decoder/fir_filter/Q_data_mult_6_buff [10]), .B(
        \u_decoder/fir_filter/Q_data_add_7_buff [10]), .CI(
        \u_decoder/fir_filter/add_332/carry [10]), .CO(
        \u_decoder/fir_filter/add_332/carry [11]), .S(
        \u_decoder/fir_filter/Q_data_add_6 [10]) );
  ADD32 \u_decoder/fir_filter/add_332/U1_11  ( .A(
        \u_decoder/fir_filter/Q_data_mult_6_buff [11]), .B(
        \u_decoder/fir_filter/Q_data_add_7_buff [11]), .CI(
        \u_decoder/fir_filter/add_332/carry [11]), .CO(
        \u_decoder/fir_filter/add_332/carry [12]), .S(
        \u_decoder/fir_filter/Q_data_add_6 [11]) );
  ADD32 \u_decoder/fir_filter/add_332/U1_12  ( .A(
        \u_decoder/fir_filter/Q_data_mult_6_buff [12]), .B(
        \u_decoder/fir_filter/Q_data_add_7_buff [12]), .CI(
        \u_decoder/fir_filter/add_332/carry [12]), .CO(
        \u_decoder/fir_filter/add_332/carry [13]), .S(
        \u_decoder/fir_filter/Q_data_add_6 [12]) );
  ADD32 \u_decoder/fir_filter/add_332/U1_13  ( .A(
        \u_decoder/fir_filter/Q_data_mult_6_buff [13]), .B(
        \u_decoder/fir_filter/Q_data_add_7_buff [13]), .CI(
        \u_decoder/fir_filter/add_332/carry [13]), .CO(
        \u_decoder/fir_filter/add_332/carry [14]), .S(
        \u_decoder/fir_filter/Q_data_add_6 [13]) );
  ADD32 \u_decoder/fir_filter/add_333/U1_1  ( .A(
        \u_decoder/fir_filter/Q_data_mult_7_buff [1]), .B(
        \u_decoder/fir_filter/Q_data_mult_8_buff [1]), .CI(
        \u_decoder/fir_filter/add_333/carry [1]), .CO(
        \u_decoder/fir_filter/add_333/carry [2]), .S(
        \u_decoder/fir_filter/Q_data_add_7 [1]) );
  ADD32 \u_decoder/fir_filter/add_333/U1_2  ( .A(
        \u_decoder/fir_filter/Q_data_mult_7_buff [2]), .B(
        \u_decoder/fir_filter/Q_data_mult_8_buff [2]), .CI(
        \u_decoder/fir_filter/add_333/carry [2]), .CO(
        \u_decoder/fir_filter/add_333/carry [3]), .S(
        \u_decoder/fir_filter/Q_data_add_7 [2]) );
  ADD32 \u_decoder/fir_filter/add_333/U1_3  ( .A(
        \u_decoder/fir_filter/Q_data_mult_7_buff [3]), .B(
        \u_decoder/fir_filter/Q_data_mult_8_buff [3]), .CI(
        \u_decoder/fir_filter/add_333/carry [3]), .CO(
        \u_decoder/fir_filter/add_333/carry [4]), .S(
        \u_decoder/fir_filter/Q_data_add_7 [3]) );
  ADD32 \u_decoder/fir_filter/add_333/U1_4  ( .A(
        \u_decoder/fir_filter/Q_data_mult_7_buff [4]), .B(
        \u_decoder/fir_filter/Q_data_mult_8_buff [4]), .CI(
        \u_decoder/fir_filter/add_333/carry [4]), .CO(
        \u_decoder/fir_filter/add_333/carry [5]), .S(
        \u_decoder/fir_filter/Q_data_add_7 [4]) );
  ADD32 \u_decoder/fir_filter/add_333/U1_5  ( .A(
        \u_decoder/fir_filter/Q_data_mult_7_buff [5]), .B(
        \u_decoder/fir_filter/Q_data_mult_8_buff [5]), .CI(
        \u_decoder/fir_filter/add_333/carry [5]), .CO(
        \u_decoder/fir_filter/add_333/carry [6]), .S(
        \u_decoder/fir_filter/Q_data_add_7 [5]) );
  ADD32 \u_decoder/fir_filter/add_333/U1_6  ( .A(
        \u_decoder/fir_filter/Q_data_mult_7_buff [6]), .B(
        \u_decoder/fir_filter/Q_data_mult_8_buff [6]), .CI(
        \u_decoder/fir_filter/add_333/carry [6]), .CO(
        \u_decoder/fir_filter/add_333/carry [7]), .S(
        \u_decoder/fir_filter/Q_data_add_7 [6]) );
  ADD32 \u_decoder/fir_filter/add_333/U1_7  ( .A(
        \u_decoder/fir_filter/Q_data_mult_7_buff [7]), .B(
        \u_decoder/fir_filter/Q_data_mult_8_buff [7]), .CI(
        \u_decoder/fir_filter/add_333/carry [7]), .CO(
        \u_decoder/fir_filter/add_333/carry [8]), .S(
        \u_decoder/fir_filter/Q_data_add_7 [7]) );
  ADD32 \u_decoder/fir_filter/add_333/U1_8  ( .A(
        \u_decoder/fir_filter/Q_data_mult_7_buff [8]), .B(
        \u_decoder/fir_filter/Q_data_mult_8_buff [8]), .CI(
        \u_decoder/fir_filter/add_333/carry [8]), .CO(
        \u_decoder/fir_filter/add_333/carry [9]), .S(
        \u_decoder/fir_filter/Q_data_add_7 [8]) );
  ADD32 \u_decoder/fir_filter/add_333/U1_9  ( .A(
        \u_decoder/fir_filter/Q_data_mult_7_buff [9]), .B(
        \u_decoder/fir_filter/Q_data_mult_8_buff [9]), .CI(
        \u_decoder/fir_filter/add_333/carry [9]), .CO(
        \u_decoder/fir_filter/add_333/carry [10]), .S(
        \u_decoder/fir_filter/Q_data_add_7 [9]) );
  ADD32 \u_decoder/fir_filter/add_333/U1_10  ( .A(
        \u_decoder/fir_filter/Q_data_mult_7_buff [10]), .B(
        \u_decoder/fir_filter/Q_data_mult_8_buff [10]), .CI(
        \u_decoder/fir_filter/add_333/carry [10]), .CO(
        \u_decoder/fir_filter/add_333/carry [11]), .S(
        \u_decoder/fir_filter/Q_data_add_7 [10]) );
  ADD32 \u_decoder/fir_filter/add_333/U1_11  ( .A(
        \u_decoder/fir_filter/Q_data_mult_7_buff [11]), .B(
        \u_decoder/fir_filter/Q_data_mult_8_buff [11]), .CI(
        \u_decoder/fir_filter/add_333/carry [11]), .CO(
        \u_decoder/fir_filter/add_333/carry [12]), .S(
        \u_decoder/fir_filter/Q_data_add_7 [11]) );
  ADD32 \u_decoder/fir_filter/add_333/U1_12  ( .A(
        \u_decoder/fir_filter/Q_data_mult_7_buff [12]), .B(
        \u_decoder/fir_filter/Q_data_mult_8_buff [12]), .CI(
        \u_decoder/fir_filter/add_333/carry [12]), .CO(
        \u_decoder/fir_filter/add_333/carry [13]), .S(
        \u_decoder/fir_filter/Q_data_add_7 [12]) );
  ADD32 \u_decoder/fir_filter/add_333/U1_13  ( .A(
        \u_decoder/fir_filter/Q_data_mult_7_buff [13]), .B(
        \u_decoder/fir_filter/Q_data_mult_8_buff [13]), .CI(
        \u_decoder/fir_filter/add_333/carry [13]), .CO(
        \u_decoder/fir_filter/add_333/carry [14]), .S(
        \u_decoder/fir_filter/Q_data_add_7 [13]) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/mult_276/S2_2_5  ( .A(n770), .B(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[1][5] ), .CI(
        \u_decoder/I_prefilter [1]), .CO(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[2][5] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/SUMB[2][5] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/mult_276/S2_3_5  ( .A(n769), .B(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[2][5] ), .CI(n770), 
        .CO(\u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[3][5] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/SUMB[3][5] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/mult_276/S2_3_3  ( .A(n769), .B(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[2][3] ), .CI(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/SUMB[1][5] ), .CO(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[3][3] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/SUMB[3][3] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/mult_276/S2_4_5  ( .A(n767), .B(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[3][5] ), .CI(n768), 
        .CO(\u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[4][5] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/SUMB[4][5] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/mult_276/S2_4_3  ( .A(n767), .B(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[3][3] ), .CI(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/SUMB[2][5] ), .CO(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[4][3] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/SUMB[4][3] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/mult_276/S1_4_0  ( .A(n766), .B(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[3][0] ), .CI(
        \u_decoder/I_prefilter [1]), .CO(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[4][0] ), .S(
        \u_decoder/fir_filter/I_data_mult_4 [4]) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/mult_276/S2_5_5  ( .A(n765), .B(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[4][5] ), .CI(n766), 
        .CO(\u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[5][5] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/SUMB[5][5] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/mult_276/S2_5_3  ( .A(n765), .B(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[4][3] ), .CI(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/SUMB[3][5] ), .CO(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[5][3] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/SUMB[5][3] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/mult_276/S1_5_0  ( .A(
        \u_decoder/I_prefilter [5]), .B(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[4][0] ), .CI(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/SUMB[2][3] ), .CO(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[5][0] ), .S(
        \u_decoder/fir_filter/I_data_mult_4 [5]) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/mult_276/S2_6_5  ( .A(n764), .B(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[5][5] ), .CI(
        \u_decoder/I_prefilter [5]), .CO(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[6][5] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/SUMB[6][5] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/mult_276/S2_6_3  ( .A(n764), .B(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[5][3] ), .CI(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/SUMB[4][5] ), .CO(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[6][3] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/SUMB[6][3] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/mult_276/S1_6_0  ( .A(
        \u_decoder/I_prefilter [6]), .B(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[5][0] ), .CI(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/SUMB[3][3] ), .CO(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[6][0] ), .S(
        \u_decoder/fir_filter/I_data_mult_4 [6]) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r167/S1_2_0  ( .A(n770), .B(
        \u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[1][0] ), .CI(
        \u_decoder/I_prefilter [1]), .CO(
        \u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[2][0] ), .S(
        \u_decoder/fir_filter/I_data_mult_3 [2]) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r167/S2_3_1  ( .A(n768), .B(
        \u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[2][1] ), .CI(
        \u_decoder/I_prefilter [1]), .CO(
        \u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[3][1] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/r167/SUMB[3][1] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r167/S1_3_0  ( .A(n769), .B(
        \u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[2][0] ), .CI(
        \u_decoder/fir_filter/dp_cluster_0/r167/SUMB[2][1] ), .CO(
        \u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[3][0] ), .S(
        \u_decoder/fir_filter/I_data_mult_3 [3]) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r167/S2_4_3  ( .A(n766), .B(
        \u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[3][3] ), .CI(
        \u_decoder/I_prefilter [1]), .CO(
        \u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[4][3] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/r167/SUMB[4][3] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r167/S2_4_1  ( .A(n766), .B(
        \u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[3][1] ), .CI(n771), 
        .CO(\u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[4][1] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/r167/SUMB[4][1] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r167/S1_4_0  ( .A(n767), .B(
        \u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[3][0] ), .CI(
        \u_decoder/fir_filter/dp_cluster_0/r167/SUMB[3][1] ), .CO(
        \u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[4][0] ), .S(
        \u_decoder/fir_filter/I_data_mult_3 [4]) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r167/S2_5_3  ( .A(
        \u_decoder/I_prefilter [5]), .B(
        \u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[4][3] ), .CI(n770), 
        .CO(\u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[5][3] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/r167/SUMB[5][3] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r167/S2_5_1  ( .A(
        \u_decoder/I_prefilter [5]), .B(
        \u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[4][1] ), .CI(
        \u_decoder/fir_filter/dp_cluster_0/r167/SUMB[3][3] ), .CO(
        \u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[5][1] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/r167/SUMB[5][1] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r167/S1_5_0  ( .A(n765), .B(
        \u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[4][0] ), .CI(
        \u_decoder/fir_filter/dp_cluster_0/r167/SUMB[4][1] ), .CO(
        \u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[5][0] ), .S(
        \u_decoder/fir_filter/I_data_mult_3 [5]) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r167/S2_6_3  ( .A(
        \u_decoder/I_prefilter [6]), .B(
        \u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[5][3] ), .CI(n769), 
        .CO(\u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[6][3] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/r167/SUMB[6][3] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r167/S2_6_1  ( .A(
        \u_decoder/I_prefilter [6]), .B(
        \u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[5][1] ), .CI(
        \u_decoder/fir_filter/dp_cluster_0/r167/SUMB[4][3] ), .CO(
        \u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[6][1] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/r167/SUMB[6][1] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r167/S1_6_0  ( .A(n764), .B(
        \u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[5][0] ), .CI(
        \u_decoder/fir_filter/dp_cluster_0/r167/SUMB[5][1] ), .CO(
        \u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[6][0] ), .S(
        \u_decoder/fir_filter/I_data_mult_3 [6]) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r166/S2_2_3  ( .A(n770), .B(
        \u_decoder/fir_filter/dp_cluster_0/r166/CARRYB[1][3] ), .CI(
        \u_decoder/I_prefilter [1]), .CO(
        \u_decoder/fir_filter/dp_cluster_0/r166/CARRYB[2][3] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/r166/SUMB[2][3] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r166/S2_3_3  ( .A(n769), .B(
        \u_decoder/fir_filter/dp_cluster_0/r166/CARRYB[2][3] ), .CI(n771), 
        .CO(\u_decoder/fir_filter/dp_cluster_0/r166/CARRYB[3][3] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/r166/SUMB[3][3] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r166/S2_3_1  ( .A(n768), .B(
        \u_decoder/fir_filter/dp_cluster_0/r166/CARRYB[2][1] ), .CI(
        \u_decoder/fir_filter/dp_cluster_0/r166/SUMB[1][3] ), .CO(
        \u_decoder/fir_filter/dp_cluster_0/r166/CARRYB[3][1] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/r166/SUMB[3][1] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r166/S2_4_3  ( .A(n767), .B(
        \u_decoder/fir_filter/dp_cluster_0/r166/CARRYB[3][3] ), .CI(n768), 
        .CO(\u_decoder/fir_filter/dp_cluster_0/r166/CARRYB[4][3] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/r166/SUMB[4][3] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r166/S2_4_1  ( .A(n766), .B(
        \u_decoder/fir_filter/dp_cluster_0/r166/CARRYB[3][1] ), .CI(
        \u_decoder/fir_filter/dp_cluster_0/r166/SUMB[2][3] ), .CO(
        \u_decoder/fir_filter/dp_cluster_0/r166/CARRYB[4][1] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/r166/SUMB[4][1] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r166/S2_5_3  ( .A(n765), .B(
        \u_decoder/fir_filter/dp_cluster_0/r166/CARRYB[4][3] ), .CI(n766), 
        .CO(\u_decoder/fir_filter/dp_cluster_0/r166/CARRYB[5][3] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/r166/SUMB[5][3] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r166/S2_5_1  ( .A(
        \u_decoder/I_prefilter [5]), .B(
        \u_decoder/fir_filter/dp_cluster_0/r166/CARRYB[4][1] ), .CI(
        \u_decoder/fir_filter/dp_cluster_0/r166/SUMB[3][3] ), .CO(
        \u_decoder/fir_filter/dp_cluster_0/r166/CARRYB[5][1] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/r166/SUMB[5][1] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r166/S2_6_3  ( .A(n764), .B(
        \u_decoder/fir_filter/dp_cluster_0/r166/CARRYB[5][3] ), .CI(
        \u_decoder/I_prefilter [5]), .CO(
        \u_decoder/fir_filter/dp_cluster_0/r166/CARRYB[6][3] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/r166/SUMB[6][3] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r166/S2_6_1  ( .A(
        \u_decoder/I_prefilter [6]), .B(
        \u_decoder/fir_filter/dp_cluster_0/r166/CARRYB[5][1] ), .CI(
        \u_decoder/fir_filter/dp_cluster_0/r166/SUMB[4][3] ), .CO(
        \u_decoder/fir_filter/dp_cluster_0/r166/CARRYB[6][1] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/r166/SUMB[6][1] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r165/S2_3_3  ( .A(n768), .B(
        \u_decoder/fir_filter/dp_cluster_0/r165/CARRYB[2][3] ), .CI(n59), .CO(
        \u_decoder/fir_filter/dp_cluster_0/r165/CARRYB[3][3] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/r165/SUMB[3][3] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r165/S2_4_3  ( .A(n766), .B(
        \u_decoder/fir_filter/dp_cluster_0/r165/CARRYB[3][3] ), .CI(n53), .CO(
        \u_decoder/fir_filter/dp_cluster_0/r165/CARRYB[4][3] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/r165/SUMB[4][3] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r165/S1_4_0  ( .A(n767), .B(
        \u_decoder/fir_filter/dp_cluster_0/r165/CARRYB[3][0] ), .CI(
        \u_decoder/I_prefilter [1]), .CO(
        \u_decoder/fir_filter/dp_cluster_0/r165/CARRYB[4][0] ), .S(
        \u_decoder/fir_filter/I_data_mult_1[4] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r165/S2_5_3  ( .A(
        \u_decoder/I_prefilter [5]), .B(
        \u_decoder/fir_filter/dp_cluster_0/r165/CARRYB[4][3] ), .CI(n69), .CO(
        \u_decoder/fir_filter/dp_cluster_0/r165/CARRYB[5][3] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/r165/SUMB[5][3] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r165/S1_5_0  ( .A(n765), .B(
        \u_decoder/fir_filter/dp_cluster_0/r165/CARRYB[4][0] ), .CI(
        \u_decoder/fir_filter/dp_cluster_0/r165/SUMB[2][3] ), .CO(
        \u_decoder/fir_filter/dp_cluster_0/r165/CARRYB[5][0] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/r165/PROD1[5] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r165/S2_6_3  ( .A(
        \u_decoder/I_prefilter [6]), .B(
        \u_decoder/fir_filter/dp_cluster_0/r165/CARRYB[5][3] ), .CI(n164), 
        .CO(\u_decoder/fir_filter/dp_cluster_0/r165/CARRYB[6][3] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/r165/SUMB[6][3] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r165/S1_6_0  ( .A(n764), .B(
        \u_decoder/fir_filter/dp_cluster_0/r165/CARRYB[5][0] ), .CI(
        \u_decoder/fir_filter/dp_cluster_0/r165/SUMB[3][3] ), .CO(
        \u_decoder/fir_filter/dp_cluster_0/r165/CARRYB[6][0] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/r165/A1[4] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r164/S2_3_2  ( .A(n768), .B(
        \u_decoder/fir_filter/dp_cluster_0/r164/CARRYB[2][2] ), .CI(n59), .CO(
        \u_decoder/fir_filter/dp_cluster_0/r164/CARRYB[3][2] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/r164/SUMB[3][2] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r164/S1_3_0  ( .A(n769), .B(
        \u_decoder/fir_filter/dp_cluster_0/r164/CARRYB[2][0] ), .CI(
        \u_decoder/I_prefilter [1]), .CO(
        \u_decoder/fir_filter/dp_cluster_0/r164/CARRYB[3][0] ), .S(
        \u_decoder/fir_filter/I_data_mult_0 [3]) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r164/S2_4_2  ( .A(n766), .B(
        \u_decoder/fir_filter/dp_cluster_0/r164/CARRYB[3][2] ), .CI(n53), .CO(
        \u_decoder/fir_filter/dp_cluster_0/r164/CARRYB[4][2] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/r164/SUMB[4][2] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r164/S1_4_0  ( .A(n767), .B(
        \u_decoder/fir_filter/dp_cluster_0/r164/CARRYB[3][0] ), .CI(
        \u_decoder/fir_filter/dp_cluster_0/r164/SUMB[2][2] ), .CO(
        \u_decoder/fir_filter/dp_cluster_0/r164/CARRYB[4][0] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/r164/PROD1[4] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r164/S2_5_2  ( .A(
        \u_decoder/I_prefilter [5]), .B(
        \u_decoder/fir_filter/dp_cluster_0/r164/CARRYB[4][2] ), .CI(n69), .CO(
        \u_decoder/fir_filter/dp_cluster_0/r164/CARRYB[5][2] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/r164/SUMB[5][2] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r164/S1_5_0  ( .A(n765), .B(
        \u_decoder/fir_filter/dp_cluster_0/r164/CARRYB[4][0] ), .CI(
        \u_decoder/fir_filter/dp_cluster_0/r164/SUMB[3][2] ), .CO(
        \u_decoder/fir_filter/dp_cluster_0/r164/CARRYB[5][0] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/r164/A1[3] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r164/S2_6_2  ( .A(
        \u_decoder/I_prefilter [6]), .B(
        \u_decoder/fir_filter/dp_cluster_0/r164/CARRYB[5][2] ), .CI(n164), 
        .CO(\u_decoder/fir_filter/dp_cluster_0/r164/CARRYB[6][2] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/r164/SUMB[6][2] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r164/S1_6_0  ( .A(n764), .B(
        \u_decoder/fir_filter/dp_cluster_0/r164/CARRYB[5][0] ), .CI(
        \u_decoder/fir_filter/dp_cluster_0/r164/SUMB[4][2] ), .CO(
        \u_decoder/fir_filter/dp_cluster_0/r164/CARRYB[6][0] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/r164/A1[4] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/mult_308/S2_2_5  ( .A(n760), .B(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[1][5] ), .CI(
        \u_decoder/Q_prefilter [1]), .CO(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[2][5] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/SUMB[2][5] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/mult_308/S2_3_5  ( .A(n759), .B(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[2][5] ), .CI(n760), 
        .CO(\u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[3][5] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/SUMB[3][5] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/mult_308/S2_3_3  ( .A(n759), .B(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[2][3] ), .CI(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/SUMB[1][5] ), .CO(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[3][3] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/SUMB[3][3] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/mult_308/S2_4_5  ( .A(n757), .B(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[3][5] ), .CI(n758), 
        .CO(\u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[4][5] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/SUMB[4][5] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/mult_308/S2_4_3  ( .A(n757), .B(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[3][3] ), .CI(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/SUMB[2][5] ), .CO(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[4][3] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/SUMB[4][3] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/mult_308/S1_4_0  ( .A(n756), .B(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[3][0] ), .CI(
        \u_decoder/Q_prefilter [1]), .CO(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[4][0] ), .S(
        \u_decoder/fir_filter/Q_data_mult_4 [4]) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/mult_308/S2_5_5  ( .A(n755), .B(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[4][5] ), .CI(n756), 
        .CO(\u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[5][5] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/SUMB[5][5] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/mult_308/S2_5_3  ( .A(n755), .B(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[4][3] ), .CI(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/SUMB[3][5] ), .CO(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[5][3] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/SUMB[5][3] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/mult_308/S1_5_0  ( .A(
        \u_decoder/Q_prefilter [5]), .B(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[4][0] ), .CI(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/SUMB[2][3] ), .CO(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[5][0] ), .S(
        \u_decoder/fir_filter/Q_data_mult_4 [5]) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/mult_308/S2_6_5  ( .A(n754), .B(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[5][5] ), .CI(
        \u_decoder/Q_prefilter [5]), .CO(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[6][5] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/SUMB[6][5] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/mult_308/S2_6_3  ( .A(n754), .B(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[5][3] ), .CI(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/SUMB[4][5] ), .CO(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[6][3] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/SUMB[6][3] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/mult_308/S1_6_0  ( .A(
        \u_decoder/Q_prefilter [6]), .B(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[5][0] ), .CI(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/SUMB[3][3] ), .CO(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[6][0] ), .S(
        \u_decoder/fir_filter/Q_data_mult_4 [6]) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r180/S1_2_0  ( .A(n760), .B(
        \u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[1][0] ), .CI(
        \u_decoder/Q_prefilter [1]), .CO(
        \u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[2][0] ), .S(
        \u_decoder/fir_filter/Q_data_mult_3 [2]) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r180/S2_3_1  ( .A(n758), .B(
        \u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[2][1] ), .CI(
        \u_decoder/Q_prefilter [1]), .CO(
        \u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[3][1] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/r180/SUMB[3][1] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r180/S1_3_0  ( .A(n759), .B(
        \u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[2][0] ), .CI(
        \u_decoder/fir_filter/dp_cluster_0/r180/SUMB[2][1] ), .CO(
        \u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[3][0] ), .S(
        \u_decoder/fir_filter/Q_data_mult_3 [3]) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r180/S2_4_3  ( .A(n756), .B(
        \u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[3][3] ), .CI(
        \u_decoder/Q_prefilter [1]), .CO(
        \u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[4][3] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/r180/SUMB[4][3] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r180/S2_4_1  ( .A(n756), .B(
        \u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[3][1] ), .CI(n761), 
        .CO(\u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[4][1] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/r180/SUMB[4][1] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r180/S1_4_0  ( .A(n757), .B(
        \u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[3][0] ), .CI(
        \u_decoder/fir_filter/dp_cluster_0/r180/SUMB[3][1] ), .CO(
        \u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[4][0] ), .S(
        \u_decoder/fir_filter/Q_data_mult_3 [4]) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r180/S2_5_3  ( .A(
        \u_decoder/Q_prefilter [5]), .B(
        \u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[4][3] ), .CI(n760), 
        .CO(\u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[5][3] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/r180/SUMB[5][3] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r180/S2_5_1  ( .A(
        \u_decoder/Q_prefilter [5]), .B(
        \u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[4][1] ), .CI(
        \u_decoder/fir_filter/dp_cluster_0/r180/SUMB[3][3] ), .CO(
        \u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[5][1] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/r180/SUMB[5][1] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r180/S1_5_0  ( .A(n755), .B(
        \u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[4][0] ), .CI(
        \u_decoder/fir_filter/dp_cluster_0/r180/SUMB[4][1] ), .CO(
        \u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[5][0] ), .S(
        \u_decoder/fir_filter/Q_data_mult_3 [5]) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r180/S2_6_3  ( .A(
        \u_decoder/Q_prefilter [6]), .B(
        \u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[5][3] ), .CI(n759), 
        .CO(\u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[6][3] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/r180/SUMB[6][3] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r180/S2_6_1  ( .A(
        \u_decoder/Q_prefilter [6]), .B(
        \u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[5][1] ), .CI(
        \u_decoder/fir_filter/dp_cluster_0/r180/SUMB[4][3] ), .CO(
        \u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[6][1] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/r180/SUMB[6][1] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r180/S1_6_0  ( .A(n754), .B(
        \u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[5][0] ), .CI(
        \u_decoder/fir_filter/dp_cluster_0/r180/SUMB[5][1] ), .CO(
        \u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[6][0] ), .S(
        \u_decoder/fir_filter/Q_data_mult_3 [6]) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r179/S2_2_3  ( .A(n760), .B(
        \u_decoder/fir_filter/dp_cluster_0/r179/CARRYB[1][3] ), .CI(
        \u_decoder/Q_prefilter [1]), .CO(
        \u_decoder/fir_filter/dp_cluster_0/r179/CARRYB[2][3] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/r179/SUMB[2][3] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r179/S2_3_3  ( .A(n759), .B(
        \u_decoder/fir_filter/dp_cluster_0/r179/CARRYB[2][3] ), .CI(n761), 
        .CO(\u_decoder/fir_filter/dp_cluster_0/r179/CARRYB[3][3] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/r179/SUMB[3][3] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r179/S2_3_1  ( .A(n758), .B(
        \u_decoder/fir_filter/dp_cluster_0/r179/CARRYB[2][1] ), .CI(
        \u_decoder/fir_filter/dp_cluster_0/r179/SUMB[1][3] ), .CO(
        \u_decoder/fir_filter/dp_cluster_0/r179/CARRYB[3][1] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/r179/SUMB[3][1] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r179/S2_4_3  ( .A(n757), .B(
        \u_decoder/fir_filter/dp_cluster_0/r179/CARRYB[3][3] ), .CI(n758), 
        .CO(\u_decoder/fir_filter/dp_cluster_0/r179/CARRYB[4][3] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/r179/SUMB[4][3] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r179/S2_4_1  ( .A(n756), .B(
        \u_decoder/fir_filter/dp_cluster_0/r179/CARRYB[3][1] ), .CI(
        \u_decoder/fir_filter/dp_cluster_0/r179/SUMB[2][3] ), .CO(
        \u_decoder/fir_filter/dp_cluster_0/r179/CARRYB[4][1] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/r179/SUMB[4][1] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r179/S2_5_3  ( .A(n755), .B(
        \u_decoder/fir_filter/dp_cluster_0/r179/CARRYB[4][3] ), .CI(n756), 
        .CO(\u_decoder/fir_filter/dp_cluster_0/r179/CARRYB[5][3] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/r179/SUMB[5][3] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r179/S2_5_1  ( .A(
        \u_decoder/Q_prefilter [5]), .B(
        \u_decoder/fir_filter/dp_cluster_0/r179/CARRYB[4][1] ), .CI(
        \u_decoder/fir_filter/dp_cluster_0/r179/SUMB[3][3] ), .CO(
        \u_decoder/fir_filter/dp_cluster_0/r179/CARRYB[5][1] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/r179/SUMB[5][1] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r179/S2_6_3  ( .A(n754), .B(
        \u_decoder/fir_filter/dp_cluster_0/r179/CARRYB[5][3] ), .CI(
        \u_decoder/Q_prefilter [5]), .CO(
        \u_decoder/fir_filter/dp_cluster_0/r179/CARRYB[6][3] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/r179/SUMB[6][3] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r179/S2_6_1  ( .A(
        \u_decoder/Q_prefilter [6]), .B(
        \u_decoder/fir_filter/dp_cluster_0/r179/CARRYB[5][1] ), .CI(
        \u_decoder/fir_filter/dp_cluster_0/r179/SUMB[4][3] ), .CO(
        \u_decoder/fir_filter/dp_cluster_0/r179/CARRYB[6][1] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/r179/SUMB[6][1] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r178/S2_3_3  ( .A(n758), .B(
        \u_decoder/fir_filter/dp_cluster_0/r178/CARRYB[2][3] ), .CI(n60), .CO(
        \u_decoder/fir_filter/dp_cluster_0/r178/CARRYB[3][3] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/r178/SUMB[3][3] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r178/S2_4_3  ( .A(n756), .B(
        \u_decoder/fir_filter/dp_cluster_0/r178/CARRYB[3][3] ), .CI(n54), .CO(
        \u_decoder/fir_filter/dp_cluster_0/r178/CARRYB[4][3] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/r178/SUMB[4][3] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r178/S1_4_0  ( .A(n757), .B(
        \u_decoder/fir_filter/dp_cluster_0/r178/CARRYB[3][0] ), .CI(
        \u_decoder/Q_prefilter [1]), .CO(
        \u_decoder/fir_filter/dp_cluster_0/r178/CARRYB[4][0] ), .S(
        \u_decoder/fir_filter/Q_data_mult_1[4] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r178/S2_5_3  ( .A(
        \u_decoder/Q_prefilter [5]), .B(
        \u_decoder/fir_filter/dp_cluster_0/r178/CARRYB[4][3] ), .CI(n70), .CO(
        \u_decoder/fir_filter/dp_cluster_0/r178/CARRYB[5][3] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/r178/SUMB[5][3] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r178/S1_5_0  ( .A(n755), .B(
        \u_decoder/fir_filter/dp_cluster_0/r178/CARRYB[4][0] ), .CI(
        \u_decoder/fir_filter/dp_cluster_0/r178/SUMB[2][3] ), .CO(
        \u_decoder/fir_filter/dp_cluster_0/r178/CARRYB[5][0] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/r178/PROD1[5] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r178/S2_6_3  ( .A(
        \u_decoder/Q_prefilter [6]), .B(
        \u_decoder/fir_filter/dp_cluster_0/r178/CARRYB[5][3] ), .CI(n165), 
        .CO(\u_decoder/fir_filter/dp_cluster_0/r178/CARRYB[6][3] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/r178/SUMB[6][3] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r178/S1_6_0  ( .A(n754), .B(
        \u_decoder/fir_filter/dp_cluster_0/r178/CARRYB[5][0] ), .CI(
        \u_decoder/fir_filter/dp_cluster_0/r178/SUMB[3][3] ), .CO(
        \u_decoder/fir_filter/dp_cluster_0/r178/CARRYB[6][0] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/r178/A1[4] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r177/S2_3_2  ( .A(n758), .B(
        \u_decoder/fir_filter/dp_cluster_0/r177/CARRYB[2][2] ), .CI(n60), .CO(
        \u_decoder/fir_filter/dp_cluster_0/r177/CARRYB[3][2] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/r177/SUMB[3][2] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r177/S1_3_0  ( .A(n759), .B(
        \u_decoder/fir_filter/dp_cluster_0/r177/CARRYB[2][0] ), .CI(
        \u_decoder/Q_prefilter [1]), .CO(
        \u_decoder/fir_filter/dp_cluster_0/r177/CARRYB[3][0] ), .S(
        \u_decoder/fir_filter/Q_data_mult_0 [3]) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r177/S2_4_2  ( .A(n756), .B(
        \u_decoder/fir_filter/dp_cluster_0/r177/CARRYB[3][2] ), .CI(n54), .CO(
        \u_decoder/fir_filter/dp_cluster_0/r177/CARRYB[4][2] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/r177/SUMB[4][2] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r177/S1_4_0  ( .A(n757), .B(
        \u_decoder/fir_filter/dp_cluster_0/r177/CARRYB[3][0] ), .CI(
        \u_decoder/fir_filter/dp_cluster_0/r177/SUMB[2][2] ), .CO(
        \u_decoder/fir_filter/dp_cluster_0/r177/CARRYB[4][0] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/r177/PROD1[4] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r177/S2_5_2  ( .A(
        \u_decoder/Q_prefilter [5]), .B(
        \u_decoder/fir_filter/dp_cluster_0/r177/CARRYB[4][2] ), .CI(n70), .CO(
        \u_decoder/fir_filter/dp_cluster_0/r177/CARRYB[5][2] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/r177/SUMB[5][2] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r177/S1_5_0  ( .A(n755), .B(
        \u_decoder/fir_filter/dp_cluster_0/r177/CARRYB[4][0] ), .CI(
        \u_decoder/fir_filter/dp_cluster_0/r177/SUMB[3][2] ), .CO(
        \u_decoder/fir_filter/dp_cluster_0/r177/CARRYB[5][0] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/r177/A1[3] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r177/S2_6_2  ( .A(
        \u_decoder/Q_prefilter [6]), .B(
        \u_decoder/fir_filter/dp_cluster_0/r177/CARRYB[5][2] ), .CI(n165), 
        .CO(\u_decoder/fir_filter/dp_cluster_0/r177/CARRYB[6][2] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/r177/SUMB[6][2] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r177/S1_6_0  ( .A(n754), .B(
        \u_decoder/fir_filter/dp_cluster_0/r177/CARRYB[5][0] ), .CI(
        \u_decoder/fir_filter/dp_cluster_0/r177/SUMB[4][2] ), .CO(
        \u_decoder/fir_filter/dp_cluster_0/r177/CARRYB[6][0] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/r177/A1[4] ) );
  ADD32 \u_decoder/iq_demod/dp_cluster_0/mult_151/S3_2_2  ( .A(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/ab[2][2] ), .B(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/CARRYB[1][2] ), .CI(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/ab[1][3] ), .CO(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/CARRYB[2][2] ), .S(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/SUMB[2][2] ) );
  ADD32 \u_decoder/iq_demod/dp_cluster_0/mult_151/S2_2_1  ( .A(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/ab[2][1] ), .B(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/CARRYB[1][1] ), .CI(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/SUMB[1][2] ), .CO(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/CARRYB[2][1] ), .S(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/SUMB[2][1] ) );
  ADD32 \u_decoder/iq_demod/dp_cluster_0/mult_151/S1_2_0  ( .A(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/ab[2][0] ), .B(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/CARRYB[1][0] ), .CI(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/SUMB[1][1] ), .CO(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/CARRYB[2][0] ), .S(
        \u_decoder/iq_demod/dp_cluster_0/mult_Q_sin_out [2]) );
  ADD32 \u_decoder/iq_demod/dp_cluster_0/mult_151/S14_3  ( .A(
        \u_decoder/iq_demod/Q_if_buff[3] ), .B(n6), .CI(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/ab[3][3] ), .CO(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/CARRYB[3][3] ), .S(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/SUMB[3][3] ) );
  ADD32 \u_decoder/iq_demod/dp_cluster_0/mult_151/S5_2  ( .A(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/ab[3][2] ), .B(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/CARRYB[2][2] ), .CI(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/ab[2][3] ), .CO(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/CARRYB[3][2] ), .S(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/SUMB[3][2] ) );
  ADD32 \u_decoder/iq_demod/dp_cluster_0/mult_151/S4_1  ( .A(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/ab[3][1] ), .B(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/CARRYB[2][1] ), .CI(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/SUMB[2][2] ), .CO(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/CARRYB[3][1] ), .S(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/SUMB[3][1] ) );
  ADD32 \u_decoder/iq_demod/dp_cluster_0/mult_151/S4_0  ( .A(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/ab[3][0] ), .B(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/CARRYB[2][0] ), .CI(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/SUMB[2][1] ), .CO(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/CARRYB[3][0] ), .S(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/SUMB[3][0] ) );
  ADD32 \u_decoder/iq_demod/dp_cluster_0/mult_151/S14_3_0  ( .A(
        \u_decoder/iq_demod/Q_if_signed [3]), .B(
        \u_decoder/iq_demod/sin_out [3]), .CI(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/SUMB[3][0] ), .CO(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/A2[2] ), .S(
        \u_decoder/iq_demod/dp_cluster_0/mult_Q_sin_out [3]) );
  ADD32 \u_decoder/iq_demod/dp_cluster_0/mult_148/S3_2_2  ( .A(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/ab[2][2] ), .B(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/CARRYB[1][2] ), .CI(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/ab[1][3] ), .CO(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/CARRYB[2][2] ), .S(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/SUMB[2][2] ) );
  ADD32 \u_decoder/iq_demod/dp_cluster_0/mult_148/S2_2_1  ( .A(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/ab[2][1] ), .B(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/CARRYB[1][1] ), .CI(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/SUMB[1][2] ), .CO(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/CARRYB[2][1] ), .S(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/SUMB[2][1] ) );
  ADD32 \u_decoder/iq_demod/dp_cluster_0/mult_148/S1_2_0  ( .A(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/ab[2][0] ), .B(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/CARRYB[1][0] ), .CI(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/SUMB[1][1] ), .CO(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/CARRYB[2][0] ), .S(
        \u_decoder/iq_demod/dp_cluster_0/mult_I_cos_out [2]) );
  ADD32 \u_decoder/iq_demod/dp_cluster_0/mult_148/S14_3  ( .A(
        \u_decoder/iq_demod/I_if_buff[3] ), .B(n5), .CI(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/ab[3][3] ), .CO(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/CARRYB[3][3] ), .S(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/SUMB[3][3] ) );
  ADD32 \u_decoder/iq_demod/dp_cluster_0/mult_148/S5_2  ( .A(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/ab[3][2] ), .B(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/CARRYB[2][2] ), .CI(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/ab[2][3] ), .CO(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/CARRYB[3][2] ), .S(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/SUMB[3][2] ) );
  ADD32 \u_decoder/iq_demod/dp_cluster_0/mult_148/S4_1  ( .A(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/ab[3][1] ), .B(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/CARRYB[2][1] ), .CI(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/SUMB[2][2] ), .CO(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/CARRYB[3][1] ), .S(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/SUMB[3][1] ) );
  ADD32 \u_decoder/iq_demod/dp_cluster_0/mult_148/S4_0  ( .A(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/ab[3][0] ), .B(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/CARRYB[2][0] ), .CI(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/SUMB[2][1] ), .CO(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/CARRYB[3][0] ), .S(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/SUMB[3][0] ) );
  ADD32 \u_decoder/iq_demod/dp_cluster_0/mult_148/S14_3_0  ( .A(
        \u_decoder/iq_demod/I_if_signed [3]), .B(
        \u_decoder/iq_demod/cos_out [3]), .CI(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/SUMB[3][0] ), .CO(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/A2[2] ), .S(
        \u_decoder/iq_demod/dp_cluster_0/mult_I_cos_out [3]) );
  ADD32 \u_decoder/iq_demod/dp_cluster_0/sub_153/U2_1  ( .A(
        \u_decoder/iq_demod/dp_cluster_0/mult_I_cos_out [1]), .B(n139), .CI(
        \u_decoder/iq_demod/dp_cluster_0/sub_153/carry [1]), .CO(
        \u_decoder/iq_demod/dp_cluster_0/sub_153/carry [2]), .S(
        \u_decoder/iq_demod/add_I_out [1]) );
  ADD32 \u_decoder/iq_demod/dp_cluster_0/sub_153/U2_2  ( .A(
        \u_decoder/iq_demod/dp_cluster_0/mult_I_cos_out [2]), .B(n1951), .CI(
        \u_decoder/iq_demod/dp_cluster_0/sub_153/carry [2]), .CO(
        \u_decoder/iq_demod/dp_cluster_0/sub_153/carry [3]), .S(
        \u_decoder/iq_demod/add_I_out [2]) );
  ADD32 \u_decoder/iq_demod/dp_cluster_0/sub_153/U2_3  ( .A(
        \u_decoder/iq_demod/dp_cluster_0/mult_I_cos_out [3]), .B(n1950), .CI(
        \u_decoder/iq_demod/dp_cluster_0/sub_153/carry [3]), .CO(
        \u_decoder/iq_demod/dp_cluster_0/sub_153/carry [4]), .S(
        \u_decoder/iq_demod/add_I_out [3]) );
  ADD32 \u_decoder/iq_demod/dp_cluster_0/sub_153/U2_4  ( .A(
        \u_decoder/iq_demod/dp_cluster_0/mult_I_cos_out [4]), .B(n67), .CI(
        \u_decoder/iq_demod/dp_cluster_0/sub_153/carry [4]), .CO(
        \u_decoder/iq_demod/dp_cluster_0/sub_153/carry [5]), .S(
        \u_decoder/iq_demod/add_I_out [4]) );
  ADD32 \u_decoder/iq_demod/dp_cluster_0/sub_153/U2_5  ( .A(
        \u_decoder/iq_demod/dp_cluster_0/mult_I_cos_out [5]), .B(n109), .CI(
        \u_decoder/iq_demod/dp_cluster_0/sub_153/carry [5]), .CO(
        \u_decoder/iq_demod/dp_cluster_0/sub_153/carry [6]), .S(
        \u_decoder/iq_demod/add_I_out [5]) );
  ADD32 \u_decoder/iq_demod/dp_cluster_0/sub_153/U2_6  ( .A(
        \u_decoder/iq_demod/dp_cluster_0/mult_I_cos_out [6]), .B(n343), .CI(
        \u_decoder/iq_demod/dp_cluster_0/sub_153/carry [6]), .CO(
        \u_decoder/iq_demod/dp_cluster_0/sub_153/carry [7]), .S(
        \u_decoder/iq_demod/add_I_out [6]) );
  ADD32 \u_decoder/iq_demod/dp_cluster_1/mult_150/S3_2_2  ( .A(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/ab[2][2] ), .B(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/CARRYB[1][2] ), .CI(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/ab[1][3] ), .CO(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/CARRYB[2][2] ), .S(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/SUMB[2][2] ) );
  ADD32 \u_decoder/iq_demod/dp_cluster_1/mult_150/S2_2_1  ( .A(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/ab[2][1] ), .B(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/CARRYB[1][1] ), .CI(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/SUMB[1][2] ), .CO(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/CARRYB[2][1] ), .S(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/SUMB[2][1] ) );
  ADD32 \u_decoder/iq_demod/dp_cluster_1/mult_150/S1_2_0  ( .A(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/ab[2][0] ), .B(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/CARRYB[1][0] ), .CI(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/SUMB[1][1] ), .CO(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/CARRYB[2][0] ), .S(
        \u_decoder/iq_demod/dp_cluster_1/mult_Q_cos_out [2]) );
  ADD32 \u_decoder/iq_demod/dp_cluster_1/mult_150/S14_3  ( .A(
        \u_decoder/iq_demod/Q_if_buff[3] ), .B(n5), .CI(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/ab[3][3] ), .CO(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/CARRYB[3][3] ), .S(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/SUMB[3][3] ) );
  ADD32 \u_decoder/iq_demod/dp_cluster_1/mult_150/S5_2  ( .A(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/ab[3][2] ), .B(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/CARRYB[2][2] ), .CI(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/ab[2][3] ), .CO(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/CARRYB[3][2] ), .S(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/SUMB[3][2] ) );
  ADD32 \u_decoder/iq_demod/dp_cluster_1/mult_150/S4_1  ( .A(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/ab[3][1] ), .B(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/CARRYB[2][1] ), .CI(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/SUMB[2][2] ), .CO(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/CARRYB[3][1] ), .S(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/SUMB[3][1] ) );
  ADD32 \u_decoder/iq_demod/dp_cluster_1/mult_150/S4_0  ( .A(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/ab[3][0] ), .B(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/CARRYB[2][0] ), .CI(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/SUMB[2][1] ), .CO(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/CARRYB[3][0] ), .S(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/SUMB[3][0] ) );
  ADD32 \u_decoder/iq_demod/dp_cluster_1/mult_150/S14_3_0  ( .A(
        \u_decoder/iq_demod/Q_if_signed [3]), .B(
        \u_decoder/iq_demod/cos_out [3]), .CI(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/SUMB[3][0] ), .CO(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/A2[2] ), .S(
        \u_decoder/iq_demod/dp_cluster_1/mult_Q_cos_out [3]) );
  ADD32 \u_decoder/iq_demod/dp_cluster_1/mult_149/S3_2_2  ( .A(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/ab[2][2] ), .B(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/CARRYB[1][2] ), .CI(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/ab[1][3] ), .CO(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/CARRYB[2][2] ), .S(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/SUMB[2][2] ) );
  ADD32 \u_decoder/iq_demod/dp_cluster_1/mult_149/S2_2_1  ( .A(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/ab[2][1] ), .B(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/CARRYB[1][1] ), .CI(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/SUMB[1][2] ), .CO(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/CARRYB[2][1] ), .S(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/SUMB[2][1] ) );
  ADD32 \u_decoder/iq_demod/dp_cluster_1/mult_149/S1_2_0  ( .A(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/ab[2][0] ), .B(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/CARRYB[1][0] ), .CI(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/SUMB[1][1] ), .CO(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/CARRYB[2][0] ), .S(
        \u_decoder/iq_demod/dp_cluster_1/mult_I_sin_out [2]) );
  ADD32 \u_decoder/iq_demod/dp_cluster_1/mult_149/S14_3  ( .A(
        \u_decoder/iq_demod/I_if_buff[3] ), .B(n6), .CI(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/ab[3][3] ), .CO(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/CARRYB[3][3] ), .S(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/SUMB[3][3] ) );
  ADD32 \u_decoder/iq_demod/dp_cluster_1/mult_149/S5_2  ( .A(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/ab[3][2] ), .B(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/CARRYB[2][2] ), .CI(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/ab[2][3] ), .CO(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/CARRYB[3][2] ), .S(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/SUMB[3][2] ) );
  ADD32 \u_decoder/iq_demod/dp_cluster_1/mult_149/S4_1  ( .A(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/ab[3][1] ), .B(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/CARRYB[2][1] ), .CI(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/SUMB[2][2] ), .CO(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/CARRYB[3][1] ), .S(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/SUMB[3][1] ) );
  ADD32 \u_decoder/iq_demod/dp_cluster_1/mult_149/S4_0  ( .A(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/ab[3][0] ), .B(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/CARRYB[2][0] ), .CI(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/SUMB[2][1] ), .CO(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/CARRYB[3][0] ), .S(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/SUMB[3][0] ) );
  ADD32 \u_decoder/iq_demod/dp_cluster_1/mult_149/S14_3_0  ( .A(
        \u_decoder/iq_demod/I_if_signed [3]), .B(
        \u_decoder/iq_demod/sin_out [3]), .CI(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/SUMB[3][0] ), .CO(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/A2[2] ), .S(
        \u_decoder/iq_demod/dp_cluster_1/mult_I_sin_out [3]) );
  ADD32 \u_decoder/iq_demod/dp_cluster_1/add_154/U1_1  ( .A(
        \u_decoder/iq_demod/dp_cluster_1/mult_I_sin_out [1]), .B(
        \u_decoder/iq_demod/dp_cluster_1/mult_Q_cos_out [1]), .CI(
        \u_decoder/iq_demod/dp_cluster_1/add_154/carry [1]), .CO(
        \u_decoder/iq_demod/dp_cluster_1/add_154/carry [2]), .S(
        \u_decoder/iq_demod/add_Q_out [1]) );
  ADD32 \u_decoder/iq_demod/dp_cluster_1/add_154/U1_2  ( .A(
        \u_decoder/iq_demod/dp_cluster_1/mult_I_sin_out [2]), .B(
        \u_decoder/iq_demod/dp_cluster_1/mult_Q_cos_out [2]), .CI(
        \u_decoder/iq_demod/dp_cluster_1/add_154/carry [2]), .CO(
        \u_decoder/iq_demod/dp_cluster_1/add_154/carry [3]), .S(
        \u_decoder/iq_demod/add_Q_out [2]) );
  ADD32 \u_decoder/iq_demod/dp_cluster_1/add_154/U1_3  ( .A(
        \u_decoder/iq_demod/dp_cluster_1/mult_I_sin_out [3]), .B(
        \u_decoder/iq_demod/dp_cluster_1/mult_Q_cos_out [3]), .CI(
        \u_decoder/iq_demod/dp_cluster_1/add_154/carry [3]), .CO(
        \u_decoder/iq_demod/dp_cluster_1/add_154/carry [4]), .S(
        \u_decoder/iq_demod/add_Q_out [3]) );
  ADD32 \u_decoder/iq_demod/dp_cluster_1/add_154/U1_4  ( .A(
        \u_decoder/iq_demod/dp_cluster_1/mult_I_sin_out [4]), .B(
        \u_decoder/iq_demod/dp_cluster_1/mult_Q_cos_out [4]), .CI(
        \u_decoder/iq_demod/dp_cluster_1/add_154/carry [4]), .CO(
        \u_decoder/iq_demod/dp_cluster_1/add_154/carry [5]), .S(
        \u_decoder/iq_demod/add_Q_out [4]) );
  ADD32 \u_decoder/iq_demod/dp_cluster_1/add_154/U1_5  ( .A(
        \u_decoder/iq_demod/dp_cluster_1/mult_I_sin_out [5]), .B(
        \u_decoder/iq_demod/dp_cluster_1/mult_Q_cos_out [5]), .CI(
        \u_decoder/iq_demod/dp_cluster_1/add_154/carry [5]), .CO(
        \u_decoder/iq_demod/dp_cluster_1/add_154/carry [6]), .S(
        \u_decoder/iq_demod/add_Q_out [5]) );
  ADD32 \u_decoder/iq_demod/dp_cluster_1/add_154/U1_6  ( .A(
        \u_decoder/iq_demod/dp_cluster_1/mult_I_sin_out [6]), .B(
        \u_decoder/iq_demod/dp_cluster_1/mult_Q_cos_out [6]), .CI(
        \u_decoder/iq_demod/dp_cluster_1/add_154/carry [6]), .CO(
        \u_decoder/iq_demod/dp_cluster_1/add_154/carry [7]), .S(
        \u_decoder/iq_demod/add_Q_out [6]) );
  ADD32 \u_outFIFO/r98/U2_1  ( .A(\u_outFIFO/outWriteCount[1] ), .B(n162), 
        .CI(\u_outFIFO/r98/carry [1]), .CO(\u_outFIFO/r98/carry [2]), .S(
        \u_outFIFO/N132 ) );
  ADD32 \u_outFIFO/r98/U2_2  ( .A(\u_outFIFO/outWriteCount[2] ), .B(n181), 
        .CI(\u_outFIFO/r98/carry [2]), .CO(\u_outFIFO/r98/carry [3]), .S(
        \u_outFIFO/N133 ) );
  ADD32 \u_outFIFO/r98/U2_3  ( .A(\u_outFIFO/outWriteCount[3] ), .B(n227), 
        .CI(\u_outFIFO/r98/carry [3]), .CO(\u_outFIFO/r98/carry [4]), .S(
        \u_outFIFO/N134 ) );
  ADD32 \u_outFIFO/r98/U2_4  ( .A(\u_outFIFO/outWriteCount[4] ), .B(n226), 
        .CI(\u_outFIFO/r98/carry [4]), .CO(\u_outFIFO/r98/carry [5]), .S(
        \u_outFIFO/N135 ) );
  ADD22 \u_outFIFO/add_255/U1_1_1  ( .A(\u_outFIFO/outWriteCount[1] ), .B(
        \u_outFIFO/outWriteCount[0] ), .CO(\u_outFIFO/add_255/carry [2]), .S(
        \u_outFIFO/N114 ) );
  ADD22 \u_outFIFO/add_255/U1_1_2  ( .A(\u_outFIFO/outWriteCount[2] ), .B(
        \u_outFIFO/add_255/carry [2]), .CO(\u_outFIFO/add_255/carry [3]), .S(
        \u_outFIFO/N115 ) );
  ADD22 \u_outFIFO/add_255/U1_1_3  ( .A(\u_outFIFO/outWriteCount[3] ), .B(
        \u_outFIFO/add_255/carry [3]), .CO(\u_outFIFO/add_255/carry [4]), .S(
        \u_outFIFO/N116 ) );
  ADD22 \u_outFIFO/add_255/U1_1_4  ( .A(\u_outFIFO/outWriteCount[4] ), .B(
        \u_outFIFO/add_255/carry [4]), .CO(\u_outFIFO/add_255/carry [5]), .S(
        \u_outFIFO/N117 ) );
  ADD22 \u_outFIFO/add_256/U1_1_1  ( .A(\u_outFIFO/i_FIFO [1]), .B(
        \u_outFIFO/i_FIFO [0]), .CO(\u_outFIFO/add_256/carry [2]), .S(
        \u_outFIFO/N120 ) );
  ADD22 \u_outFIFO/add_256/U1_1_2  ( .A(\u_outFIFO/i_FIFO [2]), .B(
        \u_outFIFO/add_256/carry [2]), .CO(\u_outFIFO/add_256/carry [3]), .S(
        \u_outFIFO/N121 ) );
  ADD22 \u_outFIFO/add_256/U1_1_3  ( .A(\u_outFIFO/i_FIFO [3]), .B(
        \u_outFIFO/add_256/carry [3]), .CO(\u_outFIFO/add_256/carry [4]), .S(
        \u_outFIFO/N122 ) );
  ADD22 \u_outFIFO/add_260/U1_1_1  ( .A(\u_outFIFO/outReadCount[1] ), .B(
        \u_outFIFO/outReadCount[0] ), .CO(\u_outFIFO/add_260/carry [2]), .S(
        \u_outFIFO/N126 ) );
  ADD22 \u_outFIFO/add_260/U1_1_2  ( .A(\u_outFIFO/outReadCount[2] ), .B(
        \u_outFIFO/add_260/carry [2]), .CO(\u_outFIFO/add_260/carry [3]), .S(
        \u_outFIFO/N127 ) );
  ADD22 \u_outFIFO/add_260/U1_1_3  ( .A(\u_outFIFO/outReadCount[3] ), .B(
        \u_outFIFO/add_260/carry [3]), .CO(\u_outFIFO/add_260/carry [4]), .S(
        \u_outFIFO/N128 ) );
  ADD22 \u_outFIFO/add_360/U1_1_1  ( .A(n943), .B(n35), .CO(
        \u_outFIFO/add_360/carry [2]), .S(\u_outFIFO/N196 ) );
  ADD22 \u_outFIFO/add_360/U1_1_2  ( .A(n774), .B(\u_outFIFO/add_360/carry [2]), .CO(\u_outFIFO/add_360/carry [3]), .S(\u_outFIFO/N197 ) );
  ADD22 \u_outFIFO/add_360/U1_1_3  ( .A(n775), .B(\u_outFIFO/add_360/carry [3]), .CO(\u_outFIFO/add_360/carry [4]), .S(\u_outFIFO/N198 ) );
  ADD22 \u_coder/add_93/U1_1_1  ( .A(\u_coder/c [1]), .B(\u_coder/c [0]), .CO(
        \u_coder/add_93/carry [2]), .S(\u_coder/N459 ) );
  ADD22 \u_coder/add_93/U1_1_2  ( .A(\u_coder/c [2]), .B(
        \u_coder/add_93/carry [2]), .CO(\u_coder/add_93/carry [3]), .S(
        \u_coder/N460 ) );
  ADD22 \u_coder/add_93/U1_1_3  ( .A(\u_coder/c [3]), .B(
        \u_coder/add_93/carry [3]), .CO(\u_coder/add_93/carry [4]), .S(
        \u_coder/N461 ) );
  ADD22 \u_coder/add_93/U1_1_4  ( .A(\u_coder/c [4]), .B(
        \u_coder/add_93/carry [4]), .CO(\u_coder/add_93/carry [5]), .S(
        \u_coder/N462 ) );
  ADD22 \u_coder/add_93/U1_1_5  ( .A(\u_coder/c [5]), .B(
        \u_coder/add_93/carry [5]), .CO(\u_coder/add_93/carry [6]), .S(
        \u_coder/N463 ) );
  ADD22 \u_coder/add_93/U1_1_6  ( .A(\u_coder/c [6]), .B(
        \u_coder/add_93/carry [6]), .CO(\u_coder/add_93/carry [7]), .S(
        \u_coder/N464 ) );
  ADD22 \u_coder/add_93/U1_1_7  ( .A(\u_coder/c [7]), .B(
        \u_coder/add_93/carry [7]), .CO(\u_coder/add_93/carry [8]), .S(
        \u_coder/N465 ) );
  ADD22 \u_coder/add_93/U1_1_8  ( .A(\u_coder/c [8]), .B(
        \u_coder/add_93/carry [8]), .CO(\u_coder/add_93/carry [9]), .S(
        \u_coder/N466 ) );
  ADD22 \u_coder/add_93/U1_1_9  ( .A(\u_coder/c [9]), .B(
        \u_coder/add_93/carry [9]), .CO(\u_coder/add_93/carry [10]), .S(
        \u_coder/N467 ) );
  ADD22 \u_coder/add_93/U1_1_10  ( .A(\u_coder/c [10]), .B(
        \u_coder/add_93/carry [10]), .CO(\u_coder/add_93/carry [11]), .S(
        \u_coder/N468 ) );
  ADD22 \u_coder/add_93/U1_1_11  ( .A(\u_coder/c [11]), .B(
        \u_coder/add_93/carry [11]), .CO(\u_coder/add_93/carry [12]), .S(
        \u_coder/N469 ) );
  ADD22 \u_coder/add_93/U1_1_12  ( .A(\u_coder/c [12]), .B(
        \u_coder/add_93/carry [12]), .CO(\u_coder/add_93/carry [13]), .S(
        \u_coder/N470 ) );
  ADD22 \u_coder/add_93/U1_1_13  ( .A(\u_coder/c [13]), .B(
        \u_coder/add_93/carry [13]), .CO(\u_coder/add_93/carry [14]), .S(
        \u_coder/N471 ) );
  ADD22 \u_coder/add_93/U1_1_14  ( .A(\u_coder/c [14]), .B(
        \u_coder/add_93/carry [14]), .CO(\u_coder/add_93/carry [15]), .S(
        \u_coder/N472 ) );
  ADD22 \u_coder/add_93/U1_1_15  ( .A(\u_coder/c [15]), .B(
        \u_coder/add_93/carry [15]), .CO(\u_coder/add_93/carry [16]), .S(
        \u_coder/N473 ) );
  ADD22 \u_coder/add_93/U1_1_16  ( .A(\u_coder/c [16]), .B(
        \u_coder/add_93/carry [16]), .CO(\u_coder/add_93/carry [17]), .S(
        \u_coder/N474 ) );
  ADD22 \u_coder/add_93/U1_1_17  ( .A(\u_coder/c [17]), .B(
        \u_coder/add_93/carry [17]), .CO(\u_coder/add_93/carry [18]), .S(
        \u_coder/N475 ) );
  ADD22 \u_coder/add_93/U1_1_18  ( .A(\u_coder/c [18]), .B(
        \u_coder/add_93/carry [18]), .CO(\u_coder/add_93/carry [19]), .S(
        \u_coder/N476 ) );
  ADD22 \u_coder/add_206/U1_1_1  ( .A(\u_coder/i [1]), .B(n778), .CO(
        \u_coder/add_206/carry [2]), .S(\u_coder/N708 ) );
  ADD22 \u_coder/add_206/U1_1_2  ( .A(\u_coder/i [2]), .B(
        \u_coder/add_206/carry [2]), .CO(\u_coder/add_206/carry [3]), .S(
        \u_coder/N709 ) );
  ADD22 \u_coder/add_206/U1_1_3  ( .A(\u_coder/i [3]), .B(
        \u_coder/add_206/carry [3]), .CO(\u_coder/add_206/carry [4]), .S(
        \u_coder/N710 ) );
  ADD22 \u_coder/add_206/U1_1_4  ( .A(\u_coder/i [4]), .B(
        \u_coder/add_206/carry [4]), .CO(\u_coder/add_206/carry [5]), .S(
        \u_coder/N711 ) );
  ADD22 \u_coder/add_206/U1_1_5  ( .A(\u_coder/i [5]), .B(
        \u_coder/add_206/carry [5]), .CO(\u_coder/add_206/carry [6]), .S(
        \u_coder/N712 ) );
  ADD22 \u_coder/add_206/U1_1_6  ( .A(\u_coder/i [6]), .B(
        \u_coder/add_206/carry [6]), .CO(\u_coder/add_206/carry [7]), .S(
        \u_coder/N713 ) );
  ADD22 \u_coder/add_206/U1_1_7  ( .A(\u_coder/i [7]), .B(
        \u_coder/add_206/carry [7]), .CO(\u_coder/add_206/carry [8]), .S(
        \u_coder/N714 ) );
  ADD22 \u_coder/add_206/U1_1_8  ( .A(\u_coder/i [8]), .B(
        \u_coder/add_206/carry [8]), .CO(\u_coder/add_206/carry [9]), .S(
        \u_coder/N715 ) );
  ADD22 \u_coder/add_206/U1_1_9  ( .A(\u_coder/i [9]), .B(
        \u_coder/add_206/carry [9]), .CO(\u_coder/add_206/carry [10]), .S(
        \u_coder/N716 ) );
  ADD22 \u_coder/add_206/U1_1_10  ( .A(\u_coder/i [10]), .B(
        \u_coder/add_206/carry [10]), .CO(\u_coder/add_206/carry [11]), .S(
        \u_coder/N717 ) );
  ADD22 \u_coder/add_206/U1_1_11  ( .A(\u_coder/i [11]), .B(
        \u_coder/add_206/carry [11]), .CO(\u_coder/add_206/carry [12]), .S(
        \u_coder/N718 ) );
  ADD22 \u_coder/add_206/U1_1_12  ( .A(\u_coder/i [12]), .B(
        \u_coder/add_206/carry [12]), .CO(\u_coder/add_206/carry [13]), .S(
        \u_coder/N719 ) );
  ADD22 \u_coder/add_206/U1_1_13  ( .A(\u_coder/i [13]), .B(
        \u_coder/add_206/carry [13]), .CO(\u_coder/add_206/carry [14]), .S(
        \u_coder/N720 ) );
  ADD22 \u_coder/add_206/U1_1_14  ( .A(\u_coder/i [14]), .B(
        \u_coder/add_206/carry [14]), .CO(\u_coder/add_206/carry [15]), .S(
        \u_coder/N721 ) );
  ADD22 \u_coder/add_206/U1_1_15  ( .A(\u_coder/i [15]), .B(
        \u_coder/add_206/carry [15]), .CO(\u_coder/add_206/carry [16]), .S(
        \u_coder/N722 ) );
  ADD22 \u_coder/add_206/U1_1_16  ( .A(\u_coder/i [16]), .B(
        \u_coder/add_206/carry [16]), .CO(\u_coder/add_206/carry [17]), .S(
        \u_coder/N723 ) );
  ADD22 \u_coder/add_206/U1_1_17  ( .A(\u_coder/i [17]), .B(
        \u_coder/add_206/carry [17]), .CO(\u_coder/add_206/carry [18]), .S(
        \u_coder/N724 ) );
  ADD22 \u_coder/add_206/U1_1_18  ( .A(\u_coder/i [18]), .B(
        \u_coder/add_206/carry [18]), .CO(\u_coder/add_206/carry [19]), .S(
        \u_coder/N725 ) );
  ADD22 \u_coder/add_282/U1_1_1  ( .A(\u_coder/j [1]), .B(n777), .CO(
        \u_coder/add_282/carry [2]), .S(\u_coder/N1014 ) );
  ADD22 \u_coder/add_282/U1_1_2  ( .A(\u_coder/j [2]), .B(
        \u_coder/add_282/carry [2]), .CO(\u_coder/add_282/carry [3]), .S(
        \u_coder/N1015 ) );
  ADD22 \u_coder/add_282/U1_1_3  ( .A(n776), .B(\u_coder/add_282/carry [3]), 
        .CO(\u_coder/add_282/carry [4]), .S(\u_coder/N1016 ) );
  ADD22 \u_coder/add_282/U1_1_4  ( .A(\u_coder/j [4]), .B(
        \u_coder/add_282/carry [4]), .CO(\u_coder/add_282/carry [5]), .S(
        \u_coder/N1017 ) );
  ADD22 \u_coder/add_282/U1_1_5  ( .A(\u_coder/j [5]), .B(
        \u_coder/add_282/carry [5]), .CO(\u_coder/add_282/carry [6]), .S(
        \u_coder/N1018 ) );
  ADD22 \u_coder/add_282/U1_1_6  ( .A(\u_coder/j [6]), .B(
        \u_coder/add_282/carry [6]), .CO(\u_coder/add_282/carry [7]), .S(
        \u_coder/N1019 ) );
  ADD22 \u_coder/add_282/U1_1_7  ( .A(\u_coder/j [7]), .B(
        \u_coder/add_282/carry [7]), .CO(\u_coder/add_282/carry [8]), .S(
        \u_coder/N1020 ) );
  ADD22 \u_coder/add_282/U1_1_8  ( .A(\u_coder/j [8]), .B(
        \u_coder/add_282/carry [8]), .CO(\u_coder/add_282/carry [9]), .S(
        \u_coder/N1021 ) );
  ADD22 \u_coder/add_282/U1_1_9  ( .A(\u_coder/j [9]), .B(
        \u_coder/add_282/carry [9]), .CO(\u_coder/add_282/carry [10]), .S(
        \u_coder/N1022 ) );
  ADD22 \u_coder/add_282/U1_1_10  ( .A(\u_coder/j [10]), .B(
        \u_coder/add_282/carry [10]), .CO(\u_coder/add_282/carry [11]), .S(
        \u_coder/N1023 ) );
  ADD22 \u_coder/add_282/U1_1_11  ( .A(\u_coder/j [11]), .B(
        \u_coder/add_282/carry [11]), .CO(\u_coder/add_282/carry [12]), .S(
        \u_coder/N1024 ) );
  ADD22 \u_coder/add_282/U1_1_12  ( .A(\u_coder/j [12]), .B(
        \u_coder/add_282/carry [12]), .CO(\u_coder/add_282/carry [13]), .S(
        \u_coder/N1025 ) );
  ADD22 \u_coder/add_282/U1_1_13  ( .A(\u_coder/j [13]), .B(
        \u_coder/add_282/carry [13]), .CO(\u_coder/add_282/carry [14]), .S(
        \u_coder/N1026 ) );
  ADD22 \u_coder/add_282/U1_1_14  ( .A(\u_coder/j [14]), .B(
        \u_coder/add_282/carry [14]), .CO(\u_coder/add_282/carry [15]), .S(
        \u_coder/N1027 ) );
  ADD22 \u_coder/add_282/U1_1_15  ( .A(\u_coder/j [15]), .B(
        \u_coder/add_282/carry [15]), .CO(\u_coder/add_282/carry [16]), .S(
        \u_coder/N1028 ) );
  ADD22 \u_coder/add_282/U1_1_16  ( .A(\u_coder/j [16]), .B(
        \u_coder/add_282/carry [16]), .CO(\u_coder/add_282/carry [17]), .S(
        \u_coder/N1029 ) );
  ADD22 \u_coder/add_282/U1_1_17  ( .A(\u_coder/j [17]), .B(
        \u_coder/add_282/carry [17]), .CO(\u_coder/add_282/carry [18]), .S(
        \u_coder/N1030 ) );
  ADD22 \u_coder/add_282/U1_1_18  ( .A(\u_coder/j [18]), .B(
        \u_coder/add_282/carry [18]), .CO(\u_coder/add_282/carry [19]), .S(
        \u_coder/N1031 ) );
  ADD32 \u_inFIFO/r96/U2_1  ( .A(\u_inFIFO/outWriteCount[1] ), .B(n161), .CI(
        \u_inFIFO/r96/carry [1]), .CO(\u_inFIFO/r96/carry [2]), .S(
        \u_inFIFO/N124 ) );
  ADD32 \u_inFIFO/r96/U2_2  ( .A(\u_inFIFO/outWriteCount[2] ), .B(n106), .CI(
        \u_inFIFO/r96/carry [2]), .CO(\u_inFIFO/r96/carry [3]), .S(
        \u_inFIFO/N125 ) );
  ADD32 \u_inFIFO/r96/U2_3  ( .A(\u_inFIFO/outWriteCount[3] ), .B(n193), .CI(
        \u_inFIFO/r96/carry [3]), .CO(\u_inFIFO/r96/carry [4]), .S(
        \u_inFIFO/N126 ) );
  ADD32 \u_inFIFO/r96/U2_4  ( .A(\u_inFIFO/outWriteCount[4] ), .B(n225), .CI(
        \u_inFIFO/r96/carry [4]), .CO(\u_inFIFO/r96/carry [5]), .S(
        \u_inFIFO/N127 ) );
  ADD22 \u_inFIFO/add_252/U1_1_1  ( .A(\u_inFIFO/outReadCount[1] ), .B(
        \u_inFIFO/outReadCount[0] ), .CO(\u_inFIFO/add_252/carry [2]), .S(
        \u_inFIFO/N113 ) );
  ADD22 \u_inFIFO/add_252/U1_1_2  ( .A(\u_inFIFO/outReadCount[2] ), .B(
        \u_inFIFO/add_252/carry [2]), .CO(\u_inFIFO/add_252/carry [3]), .S(
        \u_inFIFO/N114 ) );
  ADD22 \u_inFIFO/add_252/U1_1_3  ( .A(\u_inFIFO/outReadCount[3] ), .B(
        \u_inFIFO/add_252/carry [3]), .CO(\u_inFIFO/add_252/carry [4]), .S(
        \u_inFIFO/N115 ) );
  ADD22 \u_inFIFO/add_253/U1_1_1  ( .A(n965), .B(n34), .CO(
        \u_inFIFO/add_253/carry [2]), .S(\u_inFIFO/N118 ) );
  ADD22 \u_inFIFO/add_253/U1_1_2  ( .A(n779), .B(\u_inFIFO/add_253/carry [2]), 
        .CO(\u_inFIFO/add_253/carry [3]), .S(\u_inFIFO/N119 ) );
  ADD22 \u_inFIFO/add_253/U1_1_3  ( .A(n780), .B(\u_inFIFO/add_253/carry [3]), 
        .CO(\u_inFIFO/add_253/carry [4]), .S(\u_inFIFO/N120 ) );
  ADD22 \u_inFIFO/add_263/U1_1_1  ( .A(\u_inFIFO/outWriteCount[1] ), .B(
        \u_inFIFO/outWriteCount[0] ), .CO(\u_inFIFO/add_263/carry [2]), .S(
        \u_inFIFO/N131 ) );
  ADD22 \u_inFIFO/add_263/U1_1_2  ( .A(\u_inFIFO/outWriteCount[2] ), .B(
        \u_inFIFO/add_263/carry [2]), .CO(\u_inFIFO/add_263/carry [3]), .S(
        \u_inFIFO/N132 ) );
  ADD22 \u_inFIFO/add_263/U1_1_3  ( .A(\u_inFIFO/outWriteCount[3] ), .B(
        \u_inFIFO/add_263/carry [3]), .CO(\u_inFIFO/add_263/carry [4]), .S(
        \u_inFIFO/N133 ) );
  ADD22 \u_inFIFO/add_263/U1_1_4  ( .A(\u_inFIFO/outWriteCount[4] ), .B(
        \u_inFIFO/add_263/carry [4]), .CO(\u_inFIFO/add_263/carry [5]), .S(
        \u_inFIFO/N134 ) );
  ADD22 \u_inFIFO/add_357/U1_1_1  ( .A(\u_inFIFO/j_FIFO [1]), .B(
        \u_inFIFO/j_FIFO [0]), .CO(\u_inFIFO/add_357/carry [2]), .S(
        \u_inFIFO/N192 ) );
  ADD22 \u_inFIFO/add_357/U1_1_2  ( .A(\u_inFIFO/j_FIFO [2]), .B(
        \u_inFIFO/add_357/carry [2]), .CO(\u_inFIFO/add_357/carry [3]), .S(
        \u_inFIFO/N193 ) );
  ADD22 \u_inFIFO/add_357/U1_1_3  ( .A(\u_inFIFO/j_FIFO [3]), .B(
        \u_inFIFO/add_357/carry [3]), .CO(\u_inFIFO/add_357/carry [4]), .S(
        \u_inFIFO/N194 ) );
  DF3 \u_inFIFO/sigOutData_reg  ( .D(\u_inFIFO/n245 ), .C(inClock), .Q(
        \sig_MUX_inMUX4[0] ), .QN(\u_inFIFO/n96 ) );
  DF3 \u_inFIFO/j_FIFO_reg[4]  ( .D(n1619), .C(inClock), .Q(
        \u_inFIFO/j_FIFO [4]), .QN(\u_inFIFO/n97 ) );
  DF3 \u_inFIFO/j_FIFO_reg[3]  ( .D(n1618), .C(inClock), .Q(
        \u_inFIFO/j_FIFO [3]), .QN(\u_inFIFO/n98 ) );
  DF3 \u_inFIFO/j_FIFO_reg[2]  ( .D(n1617), .C(inClock), .Q(
        \u_inFIFO/j_FIFO [2]), .QN(\u_inFIFO/n99 ) );
  DF3 \u_inFIFO/j_FIFO_reg[1]  ( .D(n1616), .C(inClock), .Q(
        \u_inFIFO/j_FIFO [1]), .QN(\u_inFIFO/n100 ) );
  DF3 \u_inFIFO/j_FIFO_reg[0]  ( .D(n1615), .C(inClock), .Q(
        \u_inFIFO/j_FIFO [0]), .QN(\u_inFIFO/n101 ) );
  DF3 \u_inFIFO/currentState_reg[1]  ( .D(\u_inFIFO/N42 ), .C(inClock), .Q(
        \u_inFIFO/currentState [1]), .QN(\u_inFIFO/n76 ) );
  DF3 \u_inFIFO/currentState_reg[2]  ( .D(\u_inFIFO/N43 ), .C(inClock), .QN(
        \u_inFIFO/n73 ) );
  DF3 \u_inFIFO/currentState_reg[0]  ( .D(\u_inFIFO/N41 ), .C(inClock), .Q(
        \u_inFIFO/currentState [0]), .QN(\u_inFIFO/n77 ) );
  DF3 \u_inFIFO/k_FIFO_reg[1]  ( .D(\u_inFIFO/n246 ), .C(inClock), .Q(
        \u_inFIFO/N39 ), .QN(\u_inFIFO/n93 ) );
  DF3 \u_inFIFO/k_FIFO_reg[0]  ( .D(\u_inFIFO/n247 ), .C(inClock), .Q(
        \u_inFIFO/N38 ), .QN(\u_inFIFO/n94 ) );
  DF3 \u_inFIFO/currentState_reg[3]  ( .D(\u_inFIFO/N44 ), .C(inClock), .Q(
        \u_inFIFO/currentState [3]), .QN(\u_inFIFO/n26 ) );
  DF3 \u_inFIFO/sigWRCOUNT_reg[3]  ( .D(\u_inFIFO/n250 ), .C(inClock), .Q(
        \u_inFIFO/outWriteCount[3] ), .QN(\u_inFIFO/n83 ) );
  DF3 \u_inFIFO/sigWRCOUNT_reg[2]  ( .D(\u_inFIFO/n249 ), .C(inClock), .Q(
        \u_inFIFO/outWriteCount[2] ), .QN(\u_inFIFO/n84 ) );
  DF3 \u_inFIFO/sigWRCOUNT_reg[1]  ( .D(\u_inFIFO/n248 ), .C(inClock), .Q(
        \u_inFIFO/outWriteCount[1] ), .QN(\u_inFIFO/n85 ) );
  DF3 \u_inFIFO/sigWRCOUNT_reg[0]  ( .D(\u_inFIFO/n252 ), .C(inClock), .Q(
        \u_inFIFO/outWriteCount[0] ), .QN(\u_inFIFO/n86 ) );
  DF3 \u_inFIFO/sigWRCOUNT_reg[4]  ( .D(\u_inFIFO/n251 ), .C(inClock), .Q(
        \u_inFIFO/outWriteCount[4] ), .QN(\u_inFIFO/n82 ) );
  DF3 \u_inFIFO/sigRDCOUNT_reg[3]  ( .D(n1484), .C(inClock), .Q(
        \u_inFIFO/outReadCount[3] ), .QN(n193) );
  DF3 \u_inFIFO/sigRDCOUNT_reg[2]  ( .D(n1483), .C(inClock), .Q(
        \u_inFIFO/outReadCount[2] ), .QN(n106) );
  DF3 \u_inFIFO/sigRDCOUNT_reg[1]  ( .D(n1482), .C(inClock), .Q(
        \u_inFIFO/outReadCount[1] ), .QN(n161) );
  DF3 \u_inFIFO/sigRDCOUNT_reg[0]  ( .D(n1481), .C(inClock), .Q(
        \u_inFIFO/outReadCount[0] ), .QN(n105) );
  DF3 \u_inFIFO/sigRDCOUNT_reg[4]  ( .D(n1480), .C(inClock), .Q(
        \u_inFIFO/outReadCount[4] ), .QN(n225) );
  DF3 \u_inFIFO/sigWRCOUNT_reg[5]  ( .D(\u_inFIFO/n253 ), .C(inClock), .Q(
        \u_inFIFO/outWriteCount[5] ), .QN(\u_inFIFO/n78 ) );
  DF3 \u_inFIFO/i_FIFO_reg[4]  ( .D(n1479), .C(inClock), .Q(\u_inFIFO/N37 ) );
  DF3 \u_inFIFO/i_FIFO_reg[3]  ( .D(n1478), .C(inClock), .Q(\u_inFIFO/N36 ) );
  DF3 \u_inFIFO/i_FIFO_reg[2]  ( .D(n1477), .C(inClock), .Q(\u_inFIFO/N35 ) );
  DF3 \u_inFIFO/i_FIFO_reg[1]  ( .D(n1476), .C(inClock), .Q(\u_inFIFO/N34 ) );
  DF3 \u_inFIFO/i_FIFO_reg[0]  ( .D(n1475), .C(inClock), .Q(n34), .QN(n216) );
  DF3 \u_inFIFO/sigEnableCounter_reg  ( .D(\u_inFIFO/N176 ), .C(inClock), .Q(
        \u_inFIFO/sigEnableCounter ) );
  DF3 \u_coder/o_sinQ_four_reg[0]  ( .D(\u_coder/n342 ), .C(inClock), .Q(
        sig_coder_outSinQMasked[0]) );
  DF3 \u_coder/o_sinQ_four_reg[1]  ( .D(\u_coder/n341 ), .C(inClock), .Q(
        sig_coder_outSinQMasked[1]) );
  DF3 \u_coder/o_sinQ_four_reg[2]  ( .D(\u_coder/n340 ), .C(inClock), .Q(
        sig_coder_outSinQMasked[2]) );
  DF3 \u_coder/o_sinQ_four_reg[3]  ( .D(\u_coder/n339 ), .C(inClock), .Q(
        sig_coder_outSinQMasked[3]) );
  DF3 \u_coder/o_sinQ_reg[0]  ( .D(\u_coder/n337 ), .C(inClock), .Q(
        sig_coder_outSinQ[0]) );
  DF3 \u_coder/o_sinQ_reg[1]  ( .D(\u_coder/n336 ), .C(inClock), .Q(
        sig_coder_outSinQ[1]) );
  DF3 \u_coder/o_sinQ_reg[2]  ( .D(\u_coder/n335 ), .C(inClock), .Q(
        sig_coder_outSinQ[2]) );
  DF3 \u_coder/o_sinQ_reg[3]  ( .D(n1471), .C(inClock), .Q(
        sig_coder_outSinQ[3]) );
  DF3 \u_coder/o_sinI_reg[0]  ( .D(\u_coder/n334 ), .C(inClock), .Q(
        sig_coder_outSinI[0]) );
  DF3 \u_coder/o_sinI_reg[3]  ( .D(\u_coder/n333 ), .C(inClock), .Q(
        sig_coder_outSinI[3]), .QN(\u_coder/n146 ) );
  DF3 \u_coder/o_sinI_reg[1]  ( .D(n1588), .C(inClock), .Q(
        sig_coder_outSinI[1]) );
  DF3 \u_coder/o_sinI_reg[2]  ( .D(n1587), .C(inClock), .Q(
        sig_coder_outSinI[2]) );
  DF3 \u_coder/is9_reg  ( .D(\u_coder/n338 ), .C(inClock), .Q(\u_coder/is9 ), 
        .QN(\u_coder/n145 ) );
  DF3 \u_coder/o_ready_reg  ( .D(\u_coder/n344 ), .C(inClock), .Q(
        \sig_MUX_inMUX3[0] ) );
  DF3 \u_coder/o_sinI_four_reg[1]  ( .D(\u_coder/n347 ), .C(inClock), .Q(
        sig_coder_outSinIMasked[1]) );
  DF3 \u_coder/o_sinI_four_reg[2]  ( .D(\u_coder/n346 ), .C(inClock), .Q(
        sig_coder_outSinIMasked[2]) );
  DF3 \u_coder/sin_was_positiveI_reg  ( .D(\u_coder/n349 ), .C(inClock), .Q(
        \u_coder/sin_was_positiveI ), .QN(\u_coder/n140 ) );
  DF3 \u_coder/o_sinI_four_reg[3]  ( .D(\u_coder/n345 ), .C(inClock), .Q(
        sig_coder_outSinIMasked[3]) );
  DF3 \u_coder/isPositiveI_reg  ( .D(\u_coder/n350 ), .C(inClock), .Q(
        \u_coder/isPositiveI ), .QN(\u_coder/n141 ) );
  DF3 \u_coder/sin_was_positiveQ_reg  ( .D(n1474), .C(inClock), .Q(
        \u_coder/sin_was_positiveQ ) );
  DF3 \u_coder/isPositiveQ_reg  ( .D(\u_coder/n343 ), .C(inClock), .Q(
        \u_coder/isPositiveQ ), .QN(\u_coder/n144 ) );
  DF3 \u_coder/old_i_data_reg  ( .D(\u_coder/n351 ), .C(inClock), .Q(
        \u_coder/old_i_data ), .QN(n375) );
  DF3 \u_coder/o_sinI_four_reg[0]  ( .D(\u_coder/n348 ), .C(inClock), .Q(
        sig_coder_outSinIMasked[0]) );
  DF3 \u_coder/i_reg[0]  ( .D(n1592), .C(inClock), .Q(\u_coder/i [0]), .QN(
        \u_coder/n89 ) );
  DF3 \u_coder/i_reg[1]  ( .D(n1593), .C(inClock), .Q(\u_coder/i [1]), .QN(
        \u_coder/n88 ) );
  DF3 \u_coder/i_reg[2]  ( .D(n1594), .C(inClock), .Q(\u_coder/i [2]), .QN(
        \u_coder/n86 ) );
  DF3 \u_coder/i_reg[3]  ( .D(n1595), .C(inClock), .Q(\u_coder/i [3]), .QN(
        \u_coder/n85 ) );
  DF3 \u_coder/i_reg[4]  ( .D(n1596), .C(inClock), .Q(\u_coder/i [4]) );
  DF3 \u_coder/i_reg[5]  ( .D(n1597), .C(inClock), .Q(\u_coder/i [5]) );
  DF3 \u_coder/i_reg[6]  ( .D(n1598), .C(inClock), .Q(\u_coder/i [6]) );
  DF3 \u_coder/i_reg[7]  ( .D(n1599), .C(inClock), .Q(\u_coder/i [7]) );
  DF3 \u_coder/i_reg[8]  ( .D(n1600), .C(inClock), .Q(\u_coder/i [8]) );
  DF3 \u_coder/i_reg[9]  ( .D(n1601), .C(inClock), .Q(\u_coder/i [9]) );
  DF3 \u_coder/i_reg[10]  ( .D(n1602), .C(inClock), .Q(\u_coder/i [10]) );
  DF3 \u_coder/i_reg[11]  ( .D(n1603), .C(inClock), .Q(\u_coder/i [11]) );
  DF3 \u_coder/i_reg[12]  ( .D(n1604), .C(inClock), .Q(\u_coder/i [12]) );
  DF3 \u_coder/i_reg[13]  ( .D(n1605), .C(inClock), .Q(\u_coder/i [13]) );
  DF3 \u_coder/i_reg[14]  ( .D(n1606), .C(inClock), .Q(\u_coder/i [14]) );
  DF3 \u_coder/i_reg[15]  ( .D(n1607), .C(inClock), .Q(\u_coder/i [15]) );
  DF3 \u_coder/i_reg[16]  ( .D(n1608), .C(inClock), .Q(\u_coder/i [16]) );
  DF3 \u_coder/i_reg[17]  ( .D(n1609), .C(inClock), .Q(\u_coder/i [17]) );
  DF3 \u_coder/i_reg[18]  ( .D(n1610), .C(inClock), .Q(\u_coder/i [18]) );
  DF3 \u_coder/i_reg[19]  ( .D(n1591), .C(inClock), .Q(\u_coder/i [19]) );
  DF3 \u_coder/stateI_reg[0]  ( .D(\u_coder/N499 ), .C(inClock), .Q(
        \u_coder/stateI[0] ), .QN(\u_coder/n72 ) );
  DF3 \u_coder/next_stateI_reg[0]  ( .D(\u_coder/n372 ), .C(inClock), .QN(
        \u_coder/n147 ) );
  DF3 \u_coder/IorQ_reg  ( .D(\u_coder/n373 ), .C(inClock), .Q(\u_coder/IorQ ), 
        .QN(\u_coder/n139 ) );
  DF3 \u_coder/j_reg[0]  ( .D(\u_coder/n370 ), .C(inClock), .Q(\u_coder/j [0]), 
        .QN(\u_coder/n138 ) );
  DF3 \u_coder/j_reg[1]  ( .D(\u_coder/n369 ), .C(inClock), .Q(\u_coder/j [1]), 
        .QN(\u_coder/n137 ) );
  DF3 \u_coder/j_reg[2]  ( .D(\u_coder/n368 ), .C(inClock), .Q(\u_coder/j [2]), 
        .QN(\u_coder/n135 ) );
  DF3 \u_coder/j_reg[3]  ( .D(\u_coder/n367 ), .C(inClock), .Q(\u_coder/j [3]), 
        .QN(\u_coder/n134 ) );
  DF3 \u_coder/j_reg[4]  ( .D(\u_coder/n366 ), .C(inClock), .Q(\u_coder/j [4]), 
        .QN(\u_coder/n131 ) );
  DF3 \u_coder/j_reg[5]  ( .D(\u_coder/n365 ), .C(inClock), .Q(\u_coder/j [5]), 
        .QN(\u_coder/n130 ) );
  DF3 \u_coder/j_reg[6]  ( .D(\u_coder/n364 ), .C(inClock), .Q(\u_coder/j [6]), 
        .QN(\u_coder/n129 ) );
  DF3 \u_coder/j_reg[7]  ( .D(\u_coder/n363 ), .C(inClock), .Q(\u_coder/j [7]), 
        .QN(\u_coder/n128 ) );
  DF3 \u_coder/j_reg[8]  ( .D(\u_coder/n362 ), .C(inClock), .Q(\u_coder/j [8]), 
        .QN(\u_coder/n127 ) );
  DF3 \u_coder/j_reg[9]  ( .D(\u_coder/n361 ), .C(inClock), .Q(\u_coder/j [9]), 
        .QN(\u_coder/n126 ) );
  DF3 \u_coder/j_reg[10]  ( .D(\u_coder/n360 ), .C(inClock), .Q(
        \u_coder/j [10]), .QN(\u_coder/n125 ) );
  DF3 \u_coder/j_reg[11]  ( .D(\u_coder/n359 ), .C(inClock), .Q(
        \u_coder/j [11]), .QN(\u_coder/n124 ) );
  DF3 \u_coder/j_reg[12]  ( .D(\u_coder/n358 ), .C(inClock), .Q(
        \u_coder/j [12]), .QN(\u_coder/n123 ) );
  DF3 \u_coder/j_reg[13]  ( .D(\u_coder/n357 ), .C(inClock), .Q(
        \u_coder/j [13]), .QN(\u_coder/n122 ) );
  DF3 \u_coder/j_reg[14]  ( .D(\u_coder/n356 ), .C(inClock), .Q(
        \u_coder/j [14]), .QN(\u_coder/n121 ) );
  DF3 \u_coder/j_reg[15]  ( .D(\u_coder/n355 ), .C(inClock), .Q(
        \u_coder/j [15]), .QN(\u_coder/n120 ) );
  DF3 \u_coder/j_reg[16]  ( .D(\u_coder/n354 ), .C(inClock), .Q(
        \u_coder/j [16]), .QN(\u_coder/n119 ) );
  DF3 \u_coder/j_reg[17]  ( .D(\u_coder/n353 ), .C(inClock), .Q(
        \u_coder/j [17]), .QN(\u_coder/n118 ) );
  DF3 \u_coder/j_reg[18]  ( .D(\u_coder/n352 ), .C(inClock), .Q(
        \u_coder/j [18]), .QN(\u_coder/n117 ) );
  DF3 \u_coder/j_reg[19]  ( .D(\u_coder/n371 ), .C(inClock), .Q(
        \u_coder/j [19]), .QN(\u_coder/n90 ) );
  DF3 \u_coder/stateQ_reg[0]  ( .D(\u_coder/N501 ), .C(inClock), .Q(
        \u_coder/stateQ[0] ), .QN(\u_coder/n76 ) );
  DF3 \u_coder/next_stateQ_reg[0]  ( .D(\u_coder/n374 ), .C(inClock), .QN(
        \u_coder/n148 ) );
  DF3 \u_coder/clk_10M_reg  ( .D(n1757), .C(inClock), .Q(\u_coder/clk_10M ) );
  DF3 \u_coder/c_reg[19]  ( .D(\u_coder/N522 ), .C(inClock), .Q(
        \u_coder/c [19]) );
  DF3 \u_coder/c_reg[18]  ( .D(\u_coder/N521 ), .C(inClock), .Q(
        \u_coder/c [18]) );
  DF3 \u_coder/c_reg[17]  ( .D(\u_coder/N520 ), .C(inClock), .Q(
        \u_coder/c [17]) );
  DF3 \u_coder/c_reg[16]  ( .D(\u_coder/N519 ), .C(inClock), .Q(
        \u_coder/c [16]) );
  DF3 \u_coder/c_reg[15]  ( .D(\u_coder/N518 ), .C(inClock), .Q(
        \u_coder/c [15]) );
  DF3 \u_coder/c_reg[14]  ( .D(\u_coder/N517 ), .C(inClock), .Q(
        \u_coder/c [14]) );
  DF3 \u_coder/c_reg[13]  ( .D(\u_coder/N516 ), .C(inClock), .Q(
        \u_coder/c [13]) );
  DF3 \u_coder/c_reg[12]  ( .D(\u_coder/N515 ), .C(inClock), .Q(
        \u_coder/c [12]) );
  DF3 \u_coder/c_reg[11]  ( .D(\u_coder/N514 ), .C(inClock), .Q(
        \u_coder/c [11]) );
  DF3 \u_coder/c_reg[10]  ( .D(\u_coder/N513 ), .C(inClock), .Q(
        \u_coder/c [10]) );
  DF3 \u_coder/c_reg[9]  ( .D(\u_coder/N512 ), .C(inClock), .Q(\u_coder/c [9])
         );
  DF3 \u_coder/c_reg[8]  ( .D(\u_coder/N511 ), .C(inClock), .Q(\u_coder/c [8])
         );
  DF3 \u_coder/c_reg[7]  ( .D(\u_coder/N510 ), .C(inClock), .Q(\u_coder/c [7])
         );
  DF3 \u_coder/c_reg[6]  ( .D(\u_coder/N509 ), .C(inClock), .Q(\u_coder/c [6])
         );
  DF3 \u_coder/c_reg[5]  ( .D(\u_coder/N508 ), .C(inClock), .Q(\u_coder/c [5])
         );
  DF3 \u_coder/c_reg[4]  ( .D(\u_coder/N507 ), .C(inClock), .Q(\u_coder/c [4])
         );
  DF3 \u_coder/c_reg[3]  ( .D(\u_coder/N506 ), .C(inClock), .Q(\u_coder/c [3])
         );
  DF3 \u_coder/c_reg[2]  ( .D(\u_coder/N505 ), .C(inClock), .Q(\u_coder/c [2])
         );
  DF3 \u_coder/c_reg[1]  ( .D(\u_coder/N504 ), .C(inClock), .Q(\u_coder/c [1])
         );
  DF3 \u_coder/c_reg[0]  ( .D(\u_coder/N503 ), .C(inClock), .Q(\u_coder/c [0]), 
        .QN(\u_coder/n33 ) );
  DF3 \u_cordic/o_dir_reg  ( .D(\u_cordic/n37 ), .C(inClock), .Q(
        \sig_MUX_inMUX14[0] ) );
  DF3 \u_cordic/I_reg[0]  ( .D(n1671), .C(inClock), .Q(\u_cordic/I [0]) );
  DF3 \u_cordic/I_reg[1]  ( .D(n1669), .C(inClock), .Q(\u_cordic/I [1]) );
  DF3 \u_cordic/I_reg[2]  ( .D(n1667), .C(inClock), .Q(\u_cordic/I [2]) );
  DF3 \u_cordic/I_reg[3]  ( .D(n1665), .C(inClock), .Q(\u_cordic/I [3]) );
  DF3 \u_cordic/Q_reg[0]  ( .D(n1679), .C(inClock), .Q(\u_cordic/Q [0]) );
  DF3 \u_cordic/Q_reg[1]  ( .D(n1677), .C(inClock), .Q(\u_cordic/Q [1]) );
  DF3 \u_cordic/Q_reg[2]  ( .D(n1675), .C(inClock), .Q(\u_cordic/Q [2]) );
  DF3 \u_cordic/Q_reg[3]  ( .D(n1673), .C(inClock), .Q(\u_cordic/Q [3]) );
  DF3 \u_cordic/present_state_reg[1]  ( .D(\u_cordic/N16 ), .C(inClock), .Q(
        \u_cordic/present_state [1]), .QN(\u_cordic/n12 ) );
  DF3 \u_cordic/present_state_reg[2]  ( .D(\u_cordic/N17 ), .C(inClock), .Q(
        \u_cordic/present_state [2]), .QN(\u_cordic/n11 ) );
  DF3 \u_cordic/present_state_reg[0]  ( .D(\u_cordic/N15 ), .C(inClock), .Q(
        \u_cordic/present_state [0]), .QN(\u_cordic/n13 ) );
  DF3 \u_cdr/dir_reg  ( .D(\u_cdr/n49 ), .C(inClock), .Q(\u_cdr/dir ) );
  DF3 \u_cdr/cnt_reg[2]  ( .D(\u_cdr/n51 ), .C(inClock), .QN(\u_cdr/n16 ) );
  DF3 \u_cdr/cnt_reg[1]  ( .D(\u_cdr/n50 ), .C(inClock), .Q(\u_cdr/cnt [1]), 
        .QN(\u_cdr/n17 ) );
  JK3 \u_cdr/cnt_reg[0]  ( .J(\u_cdr/n32 ), .K(\u_cdr/n34 ), .C(inClock), .Q(
        \u_cdr/cnt [0]) );
  DF3 \u_cdr/flag_reg  ( .D(\u_cdr/n52 ), .C(inClock), .Q(\u_cdr/flag ), .QN(
        n315) );
  DF3 \u_cdr/cnt_d_reg[1]  ( .D(\u_cdr/n53 ), .C(inClock), .Q(\u_cdr/cnt_d [1]), .QN(\u_cdr/n14 ) );
  DF3 \u_cdr/cnt_d_reg[0]  ( .D(\u_cdr/n54 ), .C(inClock), .Q(\u_cdr/cnt_d [0]), .QN(\u_cdr/n15 ) );
  DF3 \u_cdr/cnt_in_reg[3]  ( .D(\u_cdr/n55 ), .C(inClock), .Q(
        \u_cdr/cnt_in [3]), .QN(n36) );
  DF3 \u_cdr/cnt_in_reg[2]  ( .D(\u_cdr/n56 ), .C(inClock), .Q(
        \u_cdr/cnt_in [2]), .QN(n295) );
  DF3 \u_cdr/cnt_in_reg[1]  ( .D(\u_cdr/n57 ), .C(inClock), .Q(
        \u_cdr/cnt_in [1]), .QN(n3) );
  DF3 \u_cdr/cnt_in_reg[0]  ( .D(\u_cdr/n58 ), .C(inClock), .Q(
        \u_cdr/cnt_in [0]), .QN(n294) );
  DF3 \u_outFIFO/sigOutData_reg[0]  ( .D(n1323), .C(inClock), .Q(
        sig_outFIFO_outData[0]) );
  DF3 \u_outFIFO/FIFO_reg[0][0]  ( .D(\u_outFIFO/n551 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[0][0] ) );
  DF3 \u_outFIFO/sigOutData_reg[1]  ( .D(n1324), .C(inClock), .Q(
        sig_outFIFO_outData[1]) );
  DF3 \u_outFIFO/FIFO_reg[0][1]  ( .D(\u_outFIFO/n552 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[0][1] ) );
  DF3 \u_outFIFO/sigOutData_reg[2]  ( .D(n1325), .C(inClock), .Q(
        sig_outFIFO_outData[2]) );
  DF3 \u_outFIFO/FIFO_reg[0][2]  ( .D(\u_outFIFO/n553 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[0][2] ) );
  DF3 \u_outFIFO/sigOutData_reg[3]  ( .D(n1326), .C(inClock), .Q(
        sig_outFIFO_outData[3]) );
  DF3 \u_outFIFO/FIFO_reg[0][3]  ( .D(\u_outFIFO/n554 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[0][3] ) );
  DF3 \u_outFIFO/FIFO_reg[1][0]  ( .D(\u_outFIFO/n555 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[1][0] ) );
  DF3 \u_outFIFO/FIFO_reg[1][1]  ( .D(\u_outFIFO/n556 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[1][1] ) );
  DF3 \u_outFIFO/FIFO_reg[1][2]  ( .D(\u_outFIFO/n557 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[1][2] ) );
  DF3 \u_outFIFO/FIFO_reg[1][3]  ( .D(\u_outFIFO/n558 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[1][3] ) );
  DF3 \u_outFIFO/FIFO_reg[2][0]  ( .D(\u_outFIFO/n559 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[2][0] ) );
  DF3 \u_outFIFO/FIFO_reg[2][1]  ( .D(\u_outFIFO/n560 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[2][1] ) );
  DF3 \u_outFIFO/FIFO_reg[2][2]  ( .D(\u_outFIFO/n561 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[2][2] ) );
  DF3 \u_outFIFO/FIFO_reg[2][3]  ( .D(\u_outFIFO/n562 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[2][3] ) );
  DF3 \u_outFIFO/FIFO_reg[3][0]  ( .D(\u_outFIFO/n563 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[3][0] ) );
  DF3 \u_outFIFO/FIFO_reg[3][1]  ( .D(\u_outFIFO/n564 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[3][1] ) );
  DF3 \u_outFIFO/FIFO_reg[3][2]  ( .D(\u_outFIFO/n565 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[3][2] ) );
  DF3 \u_outFIFO/FIFO_reg[3][3]  ( .D(\u_outFIFO/n566 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[3][3] ) );
  DF3 \u_outFIFO/FIFO_reg[4][0]  ( .D(\u_outFIFO/n567 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[4][0] ) );
  DF3 \u_outFIFO/FIFO_reg[4][1]  ( .D(\u_outFIFO/n568 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[4][1] ) );
  DF3 \u_outFIFO/FIFO_reg[4][2]  ( .D(\u_outFIFO/n569 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[4][2] ) );
  DF3 \u_outFIFO/FIFO_reg[4][3]  ( .D(\u_outFIFO/n570 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[4][3] ) );
  DF3 \u_outFIFO/FIFO_reg[5][0]  ( .D(\u_outFIFO/n571 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[5][0] ) );
  DF3 \u_outFIFO/FIFO_reg[5][1]  ( .D(\u_outFIFO/n572 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[5][1] ) );
  DF3 \u_outFIFO/FIFO_reg[5][2]  ( .D(\u_outFIFO/n573 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[5][2] ) );
  DF3 \u_outFIFO/FIFO_reg[5][3]  ( .D(\u_outFIFO/n574 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[5][3] ) );
  DF3 \u_outFIFO/FIFO_reg[6][0]  ( .D(\u_outFIFO/n575 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[6][0] ) );
  DF3 \u_outFIFO/FIFO_reg[6][1]  ( .D(\u_outFIFO/n576 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[6][1] ) );
  DF3 \u_outFIFO/FIFO_reg[6][2]  ( .D(\u_outFIFO/n577 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[6][2] ) );
  DF3 \u_outFIFO/FIFO_reg[6][3]  ( .D(\u_outFIFO/n578 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[6][3] ) );
  DF3 \u_outFIFO/FIFO_reg[7][0]  ( .D(\u_outFIFO/n579 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[7][0] ) );
  DF3 \u_outFIFO/FIFO_reg[7][1]  ( .D(\u_outFIFO/n580 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[7][1] ) );
  DF3 \u_outFIFO/FIFO_reg[7][2]  ( .D(\u_outFIFO/n581 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[7][2] ) );
  DF3 \u_outFIFO/FIFO_reg[7][3]  ( .D(\u_outFIFO/n582 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[7][3] ) );
  DF3 \u_outFIFO/FIFO_reg[8][0]  ( .D(\u_outFIFO/n583 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[8][0] ) );
  DF3 \u_outFIFO/FIFO_reg[8][1]  ( .D(\u_outFIFO/n584 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[8][1] ) );
  DF3 \u_outFIFO/FIFO_reg[8][2]  ( .D(\u_outFIFO/n585 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[8][2] ) );
  DF3 \u_outFIFO/FIFO_reg[8][3]  ( .D(\u_outFIFO/n586 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[8][3] ) );
  DF3 \u_outFIFO/FIFO_reg[9][0]  ( .D(\u_outFIFO/n587 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[9][0] ) );
  DF3 \u_outFIFO/FIFO_reg[9][1]  ( .D(\u_outFIFO/n588 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[9][1] ) );
  DF3 \u_outFIFO/FIFO_reg[9][2]  ( .D(\u_outFIFO/n589 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[9][2] ) );
  DF3 \u_outFIFO/FIFO_reg[9][3]  ( .D(\u_outFIFO/n590 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[9][3] ) );
  DF3 \u_outFIFO/FIFO_reg[10][0]  ( .D(\u_outFIFO/n591 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[10][0] ) );
  DF3 \u_outFIFO/FIFO_reg[10][1]  ( .D(\u_outFIFO/n592 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[10][1] ) );
  DF3 \u_outFIFO/FIFO_reg[10][2]  ( .D(\u_outFIFO/n593 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[10][2] ) );
  DF3 \u_outFIFO/FIFO_reg[10][3]  ( .D(\u_outFIFO/n594 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[10][3] ) );
  DF3 \u_outFIFO/FIFO_reg[11][0]  ( .D(\u_outFIFO/n595 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[11][0] ) );
  DF3 \u_outFIFO/FIFO_reg[11][1]  ( .D(\u_outFIFO/n596 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[11][1] ) );
  DF3 \u_outFIFO/FIFO_reg[11][2]  ( .D(\u_outFIFO/n597 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[11][2] ) );
  DF3 \u_outFIFO/FIFO_reg[11][3]  ( .D(\u_outFIFO/n598 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[11][3] ) );
  DF3 \u_outFIFO/FIFO_reg[12][0]  ( .D(\u_outFIFO/n599 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[12][0] ) );
  DF3 \u_outFIFO/FIFO_reg[12][1]  ( .D(\u_outFIFO/n600 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[12][1] ) );
  DF3 \u_outFIFO/FIFO_reg[12][2]  ( .D(\u_outFIFO/n601 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[12][2] ) );
  DF3 \u_outFIFO/FIFO_reg[12][3]  ( .D(\u_outFIFO/n602 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[12][3] ) );
  DF3 \u_outFIFO/FIFO_reg[13][0]  ( .D(\u_outFIFO/n603 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[13][0] ) );
  DF3 \u_outFIFO/FIFO_reg[13][1]  ( .D(\u_outFIFO/n604 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[13][1] ) );
  DF3 \u_outFIFO/FIFO_reg[13][2]  ( .D(\u_outFIFO/n605 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[13][2] ) );
  DF3 \u_outFIFO/FIFO_reg[13][3]  ( .D(\u_outFIFO/n606 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[13][3] ) );
  DF3 \u_outFIFO/FIFO_reg[14][0]  ( .D(\u_outFIFO/n607 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[14][0] ) );
  DF3 \u_outFIFO/FIFO_reg[14][1]  ( .D(\u_outFIFO/n608 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[14][1] ) );
  DF3 \u_outFIFO/FIFO_reg[14][2]  ( .D(\u_outFIFO/n609 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[14][2] ) );
  DF3 \u_outFIFO/FIFO_reg[14][3]  ( .D(\u_outFIFO/n610 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[14][3] ) );
  DF3 \u_outFIFO/FIFO_reg[15][0]  ( .D(\u_outFIFO/n611 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[15][0] ) );
  DF3 \u_outFIFO/FIFO_reg[15][1]  ( .D(\u_outFIFO/n612 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[15][1] ) );
  DF3 \u_outFIFO/FIFO_reg[15][2]  ( .D(\u_outFIFO/n613 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[15][2] ) );
  DF3 \u_outFIFO/FIFO_reg[15][3]  ( .D(\u_outFIFO/n614 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[15][3] ) );
  DF3 \u_outFIFO/FIFO_reg[16][0]  ( .D(\u_outFIFO/n615 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[16][0] ) );
  DF3 \u_outFIFO/FIFO_reg[16][1]  ( .D(\u_outFIFO/n616 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[16][1] ) );
  DF3 \u_outFIFO/FIFO_reg[16][2]  ( .D(\u_outFIFO/n617 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[16][2] ) );
  DF3 \u_outFIFO/FIFO_reg[16][3]  ( .D(\u_outFIFO/n618 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[16][3] ) );
  DF3 \u_outFIFO/FIFO_reg[17][0]  ( .D(\u_outFIFO/n619 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[17][0] ) );
  DF3 \u_outFIFO/FIFO_reg[17][1]  ( .D(\u_outFIFO/n620 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[17][1] ) );
  DF3 \u_outFIFO/FIFO_reg[17][2]  ( .D(\u_outFIFO/n621 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[17][2] ) );
  DF3 \u_outFIFO/FIFO_reg[17][3]  ( .D(\u_outFIFO/n622 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[17][3] ) );
  DF3 \u_outFIFO/FIFO_reg[18][0]  ( .D(\u_outFIFO/n623 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[18][0] ) );
  DF3 \u_outFIFO/FIFO_reg[18][1]  ( .D(\u_outFIFO/n624 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[18][1] ) );
  DF3 \u_outFIFO/FIFO_reg[18][2]  ( .D(\u_outFIFO/n625 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[18][2] ) );
  DF3 \u_outFIFO/FIFO_reg[18][3]  ( .D(\u_outFIFO/n626 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[18][3] ) );
  DF3 \u_outFIFO/FIFO_reg[19][0]  ( .D(\u_outFIFO/n627 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[19][0] ) );
  DF3 \u_outFIFO/FIFO_reg[19][1]  ( .D(\u_outFIFO/n628 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[19][1] ) );
  DF3 \u_outFIFO/FIFO_reg[19][2]  ( .D(\u_outFIFO/n629 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[19][2] ) );
  DF3 \u_outFIFO/FIFO_reg[19][3]  ( .D(\u_outFIFO/n630 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[19][3] ) );
  DF3 \u_outFIFO/FIFO_reg[20][0]  ( .D(\u_outFIFO/n631 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[20][0] ) );
  DF3 \u_outFIFO/FIFO_reg[20][1]  ( .D(\u_outFIFO/n632 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[20][1] ) );
  DF3 \u_outFIFO/FIFO_reg[20][2]  ( .D(\u_outFIFO/n633 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[20][2] ) );
  DF3 \u_outFIFO/FIFO_reg[20][3]  ( .D(\u_outFIFO/n634 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[20][3] ) );
  DF3 \u_outFIFO/FIFO_reg[21][0]  ( .D(\u_outFIFO/n635 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[21][0] ) );
  DF3 \u_outFIFO/FIFO_reg[21][1]  ( .D(\u_outFIFO/n636 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[21][1] ) );
  DF3 \u_outFIFO/FIFO_reg[21][2]  ( .D(\u_outFIFO/n637 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[21][2] ) );
  DF3 \u_outFIFO/FIFO_reg[21][3]  ( .D(\u_outFIFO/n638 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[21][3] ) );
  DF3 \u_outFIFO/FIFO_reg[22][0]  ( .D(\u_outFIFO/n639 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[22][0] ) );
  DF3 \u_outFIFO/FIFO_reg[22][1]  ( .D(\u_outFIFO/n640 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[22][1] ) );
  DF3 \u_outFIFO/FIFO_reg[22][2]  ( .D(\u_outFIFO/n641 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[22][2] ) );
  DF3 \u_outFIFO/FIFO_reg[22][3]  ( .D(\u_outFIFO/n642 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[22][3] ) );
  DF3 \u_outFIFO/FIFO_reg[23][0]  ( .D(\u_outFIFO/n643 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[23][0] ) );
  DF3 \u_outFIFO/FIFO_reg[23][1]  ( .D(\u_outFIFO/n644 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[23][1] ) );
  DF3 \u_outFIFO/FIFO_reg[23][2]  ( .D(\u_outFIFO/n645 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[23][2] ) );
  DF3 \u_outFIFO/FIFO_reg[23][3]  ( .D(\u_outFIFO/n646 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[23][3] ) );
  DF3 \u_outFIFO/FIFO_reg[24][0]  ( .D(\u_outFIFO/n647 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[24][0] ) );
  DF3 \u_outFIFO/FIFO_reg[24][1]  ( .D(\u_outFIFO/n648 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[24][1] ) );
  DF3 \u_outFIFO/FIFO_reg[24][2]  ( .D(\u_outFIFO/n649 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[24][2] ) );
  DF3 \u_outFIFO/FIFO_reg[24][3]  ( .D(\u_outFIFO/n650 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[24][3] ) );
  DF3 \u_outFIFO/FIFO_reg[25][0]  ( .D(\u_outFIFO/n651 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[25][0] ) );
  DF3 \u_outFIFO/FIFO_reg[25][1]  ( .D(\u_outFIFO/n652 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[25][1] ) );
  DF3 \u_outFIFO/FIFO_reg[25][2]  ( .D(\u_outFIFO/n653 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[25][2] ) );
  DF3 \u_outFIFO/FIFO_reg[25][3]  ( .D(\u_outFIFO/n654 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[25][3] ) );
  DF3 \u_outFIFO/FIFO_reg[26][0]  ( .D(\u_outFIFO/n655 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[26][0] ) );
  DF3 \u_outFIFO/FIFO_reg[26][1]  ( .D(\u_outFIFO/n656 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[26][1] ) );
  DF3 \u_outFIFO/FIFO_reg[26][2]  ( .D(\u_outFIFO/n657 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[26][2] ) );
  DF3 \u_outFIFO/FIFO_reg[26][3]  ( .D(\u_outFIFO/n658 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[26][3] ) );
  DF3 \u_outFIFO/FIFO_reg[27][0]  ( .D(\u_outFIFO/n659 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[27][0] ) );
  DF3 \u_outFIFO/FIFO_reg[27][1]  ( .D(\u_outFIFO/n660 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[27][1] ) );
  DF3 \u_outFIFO/FIFO_reg[27][2]  ( .D(\u_outFIFO/n661 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[27][2] ) );
  DF3 \u_outFIFO/FIFO_reg[27][3]  ( .D(\u_outFIFO/n662 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[27][3] ) );
  DF3 \u_outFIFO/FIFO_reg[28][0]  ( .D(\u_outFIFO/n663 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[28][0] ) );
  DF3 \u_outFIFO/FIFO_reg[28][1]  ( .D(\u_outFIFO/n664 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[28][1] ) );
  DF3 \u_outFIFO/FIFO_reg[28][2]  ( .D(\u_outFIFO/n665 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[28][2] ) );
  DF3 \u_outFIFO/FIFO_reg[28][3]  ( .D(\u_outFIFO/n666 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[28][3] ) );
  DF3 \u_outFIFO/FIFO_reg[29][0]  ( .D(\u_outFIFO/n667 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[29][0] ) );
  DF3 \u_outFIFO/FIFO_reg[29][1]  ( .D(\u_outFIFO/n668 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[29][1] ) );
  DF3 \u_outFIFO/FIFO_reg[29][2]  ( .D(\u_outFIFO/n669 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[29][2] ) );
  DF3 \u_outFIFO/FIFO_reg[29][3]  ( .D(\u_outFIFO/n670 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[29][3] ) );
  DF3 \u_outFIFO/FIFO_reg[30][0]  ( .D(\u_outFIFO/n671 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[30][0] ) );
  DF3 \u_outFIFO/FIFO_reg[30][1]  ( .D(\u_outFIFO/n672 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[30][1] ) );
  DF3 \u_outFIFO/FIFO_reg[30][2]  ( .D(\u_outFIFO/n673 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[30][2] ) );
  DF3 \u_outFIFO/FIFO_reg[30][3]  ( .D(\u_outFIFO/n674 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[30][3] ) );
  DF3 \u_outFIFO/FIFO_reg[31][0]  ( .D(\u_outFIFO/n675 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[31][0] ) );
  DF3 \u_outFIFO/FIFO_reg[31][1]  ( .D(\u_outFIFO/n676 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[31][1] ) );
  DF3 \u_outFIFO/FIFO_reg[31][2]  ( .D(\u_outFIFO/n677 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[31][2] ) );
  DF3 \u_outFIFO/FIFO_reg[31][3]  ( .D(\u_outFIFO/n678 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[31][3] ) );
  DF3 \u_outFIFO/j_FIFO_reg[4]  ( .D(n1331), .C(inClock), .Q(\u_outFIFO/N39 )
         );
  DF3 \u_outFIFO/j_FIFO_reg[3]  ( .D(n1330), .C(inClock), .Q(\u_outFIFO/N38 )
         );
  DF3 \u_outFIFO/j_FIFO_reg[2]  ( .D(n1329), .C(inClock), .Q(\u_outFIFO/N37 )
         );
  DF3 \u_outFIFO/j_FIFO_reg[1]  ( .D(n1328), .C(inClock), .Q(\u_outFIFO/N36 )
         );
  DF3 \u_outFIFO/j_FIFO_reg[0]  ( .D(n1327), .C(inClock), .Q(n35), .QN(n215)
         );
  DF3 \u_outFIFO/currentState_reg[3]  ( .D(\u_outFIFO/N44 ), .C(inClock), .QN(
        \u_outFIFO/n173 ) );
  DF3 \u_outFIFO/currentState_reg[1]  ( .D(\u_outFIFO/N42 ), .C(inClock), .Q(
        \u_outFIFO/currentState [1]), .QN(\u_outFIFO/n176 ) );
  DF3 \u_outFIFO/currentState_reg[0]  ( .D(\u_outFIFO/N41 ), .C(inClock), .Q(
        \u_outFIFO/currentState [0]), .QN(\u_outFIFO/n177 ) );
  DF3 \u_outFIFO/k_FIFO_reg[1]  ( .D(\u_outFIFO/n679 ), .C(inClock), .Q(
        \u_outFIFO/k_FIFO [1]), .QN(\u_outFIFO/n195 ) );
  JK3 \u_outFIFO/k_FIFO_reg[0]  ( .J(n815), .K(n955), .C(inClock), .Q(
        \u_outFIFO/k_FIFO [0]), .QN(\u_outFIFO/n196 ) );
  DF3 \u_outFIFO/currentState_reg[2]  ( .D(\u_outFIFO/N43 ), .C(inClock), .Q(
        \u_outFIFO/currentState [2]), .QN(\u_outFIFO/n174 ) );
  DF3 \u_outFIFO/sigWRCOUNT_reg[3]  ( .D(\u_outFIFO/n681 ), .C(inClock), .Q(
        \u_outFIFO/outWriteCount[3] ), .QN(\u_outFIFO/n181 ) );
  DF3 \u_outFIFO/sigWRCOUNT_reg[2]  ( .D(\u_outFIFO/n682 ), .C(inClock), .Q(
        \u_outFIFO/outWriteCount[2] ), .QN(\u_outFIFO/n182 ) );
  DF3 \u_outFIFO/sigWRCOUNT_reg[1]  ( .D(\u_outFIFO/n683 ), .C(inClock), .Q(
        \u_outFIFO/outWriteCount[1] ), .QN(\u_outFIFO/n183 ) );
  DF3 \u_outFIFO/sigWRCOUNT_reg[0]  ( .D(\u_outFIFO/n684 ), .C(inClock), .Q(
        \u_outFIFO/outWriteCount[0] ), .QN(\u_outFIFO/n184 ) );
  DF3 \u_outFIFO/sigWRCOUNT_reg[4]  ( .D(\u_outFIFO/n680 ), .C(inClock), .Q(
        \u_outFIFO/outWriteCount[4] ), .QN(\u_outFIFO/n180 ) );
  DF3 \u_outFIFO/sigRDCOUNT_reg[4]  ( .D(n1461), .C(inClock), .Q(
        \u_outFIFO/outReadCount[4] ), .QN(n226) );
  DF3 \u_outFIFO/sigRDCOUNT_reg[3]  ( .D(n1462), .C(inClock), .Q(
        \u_outFIFO/outReadCount[3] ), .QN(n227) );
  DF3 \u_outFIFO/sigRDCOUNT_reg[2]  ( .D(n1463), .C(inClock), .Q(
        \u_outFIFO/outReadCount[2] ), .QN(n181) );
  DF3 \u_outFIFO/sigRDCOUNT_reg[1]  ( .D(n1464), .C(inClock), .Q(
        \u_outFIFO/outReadCount[1] ), .QN(n162) );
  DF3 \u_outFIFO/sigRDCOUNT_reg[0]  ( .D(n1465), .C(inClock), .Q(
        \u_outFIFO/outReadCount[0] ), .QN(n154) );
  DF3 \u_outFIFO/sigWRCOUNT_reg[5]  ( .D(\u_outFIFO/n685 ), .C(inClock), .Q(
        \u_outFIFO/outWriteCount[5] ), .QN(\u_outFIFO/n178 ) );
  DF3 \u_outFIFO/i_FIFO_reg[4]  ( .D(\u_outFIFO/n686 ), .C(inClock), .Q(
        \u_outFIFO/i_FIFO [4]), .QN(\u_outFIFO/n185 ) );
  DF3 \u_outFIFO/i_FIFO_reg[3]  ( .D(\u_outFIFO/n687 ), .C(inClock), .Q(
        \u_outFIFO/i_FIFO [3]), .QN(\u_outFIFO/n191 ) );
  DF3 \u_outFIFO/i_FIFO_reg[2]  ( .D(\u_outFIFO/n688 ), .C(inClock), .Q(
        \u_outFIFO/i_FIFO [2]), .QN(\u_outFIFO/n192 ) );
  DF3 \u_outFIFO/i_FIFO_reg[1]  ( .D(\u_outFIFO/n689 ), .C(inClock), .Q(
        \u_outFIFO/i_FIFO [1]), .QN(\u_outFIFO/n193 ) );
  DF3 \u_outFIFO/i_FIFO_reg[0]  ( .D(\u_outFIFO/n690 ), .C(inClock), .Q(
        \u_outFIFO/i_FIFO [0]), .QN(\u_outFIFO/n194 ) );
  DF3 \u_outFIFO/sigEnableCounter_reg  ( .D(\u_outFIFO/N178 ), .C(inClock), 
        .Q(\u_outFIFO/sigEnableCounter ), .QN(\u_outFIFO/n197 ) );
  DF3 \u_decoder/iq_demod/o_I_prefilter_reg[0]  ( .D(n1837), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_0 [0]), .QN(n51) );
  DF3 \u_decoder/iq_demod/o_I_prefilter_reg[1]  ( .D(n1862), .C(inClock), .Q(
        \u_decoder/I_prefilter [1]), .QN(n59) );
  DF3 \u_decoder/iq_demod/o_I_prefilter_reg[2]  ( .D(n1864), .C(inClock), .Q(
        \u_decoder/I_prefilter [2]), .QN(n53) );
  DF3 \u_decoder/iq_demod/o_I_prefilter_reg[3]  ( .D(n1865), .C(inClock), .Q(
        \u_decoder/I_prefilter [3]), .QN(n69) );
  DF3 \u_decoder/iq_demod/o_I_prefilter_reg[4]  ( .D(n1866), .C(inClock), .Q(
        \u_decoder/I_prefilter [4]), .QN(n164) );
  DF3 \u_decoder/iq_demod/o_I_prefilter_reg[5]  ( .D(n1867), .C(inClock), .Q(
        \u_decoder/I_prefilter [5]), .QN(n30) );
  DF3 \u_decoder/iq_demod/o_I_prefilter_reg[6]  ( .D(n1869), .C(inClock), .Q(
        \u_decoder/I_prefilter [6]), .QN(n37) );
  DF3 \u_decoder/iq_demod/o_I_prefilter_reg[7]  ( .D(n1870), .C(inClock), .Q(
        \u_decoder/I_prefilter [7]), .QN(n229) );
  DF3 \u_decoder/iq_demod/o_Q_prefilter_reg[0]  ( .D(n1908), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_0 [0]), .QN(n52) );
  DF3 \u_decoder/iq_demod/o_Q_prefilter_reg[1]  ( .D(n1933), .C(inClock), .Q(
        \u_decoder/Q_prefilter [1]), .QN(n60) );
  DF3 \u_decoder/iq_demod/o_Q_prefilter_reg[2]  ( .D(n1935), .C(inClock), .Q(
        \u_decoder/Q_prefilter [2]), .QN(n54) );
  DF3 \u_decoder/iq_demod/o_Q_prefilter_reg[3]  ( .D(n1936), .C(inClock), .Q(
        \u_decoder/Q_prefilter [3]), .QN(n70) );
  DF3 \u_decoder/iq_demod/o_Q_prefilter_reg[4]  ( .D(n1937), .C(inClock), .Q(
        \u_decoder/Q_prefilter [4]), .QN(n165) );
  DF3 \u_decoder/iq_demod/o_Q_prefilter_reg[5]  ( .D(n1938), .C(inClock), .Q(
        \u_decoder/Q_prefilter [5]), .QN(n31) );
  DF3 \u_decoder/iq_demod/o_Q_prefilter_reg[6]  ( .D(n1940), .C(inClock), .Q(
        \u_decoder/Q_prefilter [6]), .QN(n38) );
  DF3 \u_decoder/iq_demod/o_Q_prefilter_reg[7]  ( .D(n1941), .C(inClock), .Q(
        \u_decoder/Q_prefilter [7]), .QN(n230) );
  DF3 \u_decoder/iq_demod/o_sample_ready_reg  ( .D(n1942), .C(inClock), .Q(
        \u_decoder/sample_ready ), .QN(n314) );
  DF3 \u_decoder/iq_demod/Q_if_buff_reg[0]  ( .D(n1322), .C(inClock), .Q(
        \u_decoder/iq_demod/Q_if_signed [0]), .QN(n104) );
  DF3 \u_decoder/iq_demod/Q_if_buff_reg[1]  ( .D(n1321), .C(inClock), .Q(
        \u_decoder/iq_demod/Q_if_signed [1]), .QN(n101) );
  DF3 \u_decoder/iq_demod/Q_if_buff_reg[2]  ( .D(n1320), .C(inClock), .Q(
        \u_decoder/iq_demod/Q_if_signed [2]), .QN(n125) );
  DF3 \u_decoder/iq_demod/Q_if_buff_reg[3]  ( .D(n1319), .C(inClock), .Q(
        \u_decoder/iq_demod/Q_if_buff[3] ), .QN(
        \u_decoder/iq_demod/Q_if_signed [3]) );
  DF3 \u_decoder/iq_demod/I_if_buff_reg[0]  ( .D(n1318), .C(inClock), .Q(
        \u_decoder/iq_demod/I_if_signed [0]), .QN(n103) );
  DF3 \u_decoder/iq_demod/I_if_buff_reg[1]  ( .D(n1317), .C(inClock), .Q(
        \u_decoder/iq_demod/I_if_signed [1]), .QN(n102) );
  DF3 \u_decoder/iq_demod/I_if_buff_reg[2]  ( .D(n1316), .C(inClock), .Q(
        \u_decoder/iq_demod/I_if_signed [2]), .QN(n126) );
  DF3 \u_decoder/iq_demod/I_if_buff_reg[3]  ( .D(n1315), .C(inClock), .Q(
        \u_decoder/iq_demod/I_if_buff[3] ), .QN(
        \u_decoder/iq_demod/I_if_signed [3]) );
  DF3 \u_decoder/iq_demod/state_reg[1]  ( .D(n1583), .C(inClock), .Q(
        \u_decoder/iq_demod/state [1]) );
  DF3 \u_decoder/iq_demod/state_reg[0]  ( .D(\u_decoder/iq_demod/N13 ), .C(
        inClock), .Q(\u_decoder/iq_demod/state [0]), .QN(
        \u_decoder/iq_demod/n30 ) );
  DF3 \u_decoder/fir_filter/o_Q_postfilter_reg[3]  ( .D(n1962), .C(inClock), 
        .Q(sig_decod_outQ[3]) );
  DF3 \u_decoder/fir_filter/o_Q_postfilter_reg[2]  ( .D(n1963), .C(inClock), 
        .Q(sig_decod_outQ[2]) );
  DF3 \u_decoder/fir_filter/o_Q_postfilter_reg[1]  ( .D(n1964), .C(inClock), 
        .Q(sig_decod_outQ[1]) );
  DF3 \u_decoder/fir_filter/o_Q_postfilter_reg[0]  ( .D(n1965), .C(inClock), 
        .Q(sig_decod_outQ[0]) );
  DF3 \u_decoder/fir_filter/Q_data_add_1_buff_reg[14]  ( .D(n1966), .C(inClock), .Q(\u_decoder/fir_filter/Q_data_add_1_buff [14]) );
  DF3 \u_decoder/fir_filter/Q_data_add_1_buff_reg[13]  ( .D(n1967), .C(inClock), .Q(\u_decoder/fir_filter/Q_data_add_1_buff [13]) );
  DF3 \u_decoder/fir_filter/Q_data_add_1_buff_reg[12]  ( .D(n1968), .C(inClock), .Q(\u_decoder/fir_filter/Q_data_add_1_buff [12]) );
  DF3 \u_decoder/fir_filter/Q_data_add_1_buff_reg[11]  ( .D(n1969), .C(inClock), .Q(\u_decoder/fir_filter/Q_data_add_1_buff [11]) );
  DF3 \u_decoder/fir_filter/Q_data_add_1_buff_reg[10]  ( .D(n1970), .C(inClock), .Q(\u_decoder/fir_filter/Q_data_add_1_buff [10]) );
  DF3 \u_decoder/fir_filter/Q_data_add_1_buff_reg[9]  ( .D(n1973), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_1_buff [9]) );
  DF3 \u_decoder/fir_filter/Q_data_add_1_buff_reg[8]  ( .D(n1974), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_1_buff [8]) );
  DF3 \u_decoder/fir_filter/Q_data_add_1_buff_reg[7]  ( .D(n1977), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_1_buff [7]) );
  DF3 \u_decoder/fir_filter/Q_data_add_1_buff_reg[6]  ( .D(n1978), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_1_buff [6]) );
  DF3 \u_decoder/fir_filter/Q_data_add_1_buff_reg[5]  ( .D(n1980), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_1_buff [5]) );
  DF3 \u_decoder/fir_filter/Q_data_add_1_buff_reg[4]  ( .D(n1982), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_1_buff [4]) );
  DF3 \u_decoder/fir_filter/Q_data_add_1_buff_reg[3]  ( .D(n1984), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_1_buff [3]) );
  DF3 \u_decoder/fir_filter/Q_data_add_1_buff_reg[2]  ( .D(n1986), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_1_buff [2]) );
  DF3 \u_decoder/fir_filter/Q_data_add_1_buff_reg[1]  ( .D(n1988), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_1_buff [1]), .QN(n7) );
  DF3 \u_decoder/fir_filter/Q_data_add_1_buff_reg[0]  ( .D(n1989), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_1_buff [0]) );
  DF3 \u_decoder/fir_filter/Q_data_add_2_buff_reg[14]  ( .D(n1990), .C(inClock), .Q(\u_decoder/fir_filter/Q_data_add_2_buff [14]) );
  DF3 \u_decoder/fir_filter/Q_data_add_2_buff_reg[13]  ( .D(n1991), .C(inClock), .Q(\u_decoder/fir_filter/Q_data_add_2_buff [13]) );
  DF3 \u_decoder/fir_filter/Q_data_add_2_buff_reg[12]  ( .D(n1992), .C(inClock), .Q(\u_decoder/fir_filter/Q_data_add_2_buff [12]) );
  DF3 \u_decoder/fir_filter/Q_data_add_2_buff_reg[11]  ( .D(n1993), .C(inClock), .Q(\u_decoder/fir_filter/Q_data_add_2_buff [11]) );
  DF3 \u_decoder/fir_filter/Q_data_add_2_buff_reg[10]  ( .D(n1994), .C(inClock), .Q(\u_decoder/fir_filter/Q_data_add_2_buff [10]) );
  DF3 \u_decoder/fir_filter/Q_data_add_2_buff_reg[9]  ( .D(n1995), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_2_buff [9]) );
  DF3 \u_decoder/fir_filter/Q_data_add_2_buff_reg[8]  ( .D(n1996), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_2_buff [8]) );
  DF3 \u_decoder/fir_filter/Q_data_add_2_buff_reg[7]  ( .D(n1997), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_2_buff [7]) );
  DF3 \u_decoder/fir_filter/Q_data_add_2_buff_reg[6]  ( .D(n1998), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_2_buff [6]) );
  DF3 \u_decoder/fir_filter/Q_data_add_2_buff_reg[5]  ( .D(n1999), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_2_buff [5]) );
  DF3 \u_decoder/fir_filter/Q_data_add_2_buff_reg[4]  ( .D(n2000), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_2_buff [4]) );
  DF3 \u_decoder/fir_filter/Q_data_add_2_buff_reg[3]  ( .D(n2001), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_2_buff [3]) );
  DF3 \u_decoder/fir_filter/Q_data_add_2_buff_reg[2]  ( .D(n2002), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_2_buff [2]) );
  DF3 \u_decoder/fir_filter/Q_data_add_2_buff_reg[1]  ( .D(n2003), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_2_buff [1]) );
  DF3 \u_decoder/fir_filter/Q_data_add_2_buff_reg[0]  ( .D(n2004), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_2_buff [0]), .QN(n100) );
  DF3 \u_decoder/fir_filter/Q_data_add_3_buff_reg[14]  ( .D(n2005), .C(inClock), .Q(\u_decoder/fir_filter/Q_data_add_3_buff [14]) );
  DF3 \u_decoder/fir_filter/Q_data_add_3_buff_reg[13]  ( .D(n2006), .C(inClock), .Q(\u_decoder/fir_filter/Q_data_add_3_buff [13]) );
  DF3 \u_decoder/fir_filter/Q_data_add_3_buff_reg[12]  ( .D(n2007), .C(inClock), .Q(\u_decoder/fir_filter/Q_data_add_3_buff [12]) );
  DF3 \u_decoder/fir_filter/Q_data_add_3_buff_reg[11]  ( .D(n2008), .C(inClock), .Q(\u_decoder/fir_filter/Q_data_add_3_buff [11]) );
  DF3 \u_decoder/fir_filter/Q_data_add_3_buff_reg[10]  ( .D(n2009), .C(inClock), .Q(\u_decoder/fir_filter/Q_data_add_3_buff [10]) );
  DF3 \u_decoder/fir_filter/Q_data_add_3_buff_reg[9]  ( .D(n2010), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_3_buff [9]) );
  DF3 \u_decoder/fir_filter/Q_data_add_3_buff_reg[8]  ( .D(n2011), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_3_buff [8]) );
  DF3 \u_decoder/fir_filter/Q_data_add_3_buff_reg[7]  ( .D(n2012), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_3_buff [7]) );
  DF3 \u_decoder/fir_filter/Q_data_add_3_buff_reg[6]  ( .D(n2013), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_3_buff [6]) );
  DF3 \u_decoder/fir_filter/Q_data_add_3_buff_reg[5]  ( .D(n2014), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_3_buff [5]) );
  DF3 \u_decoder/fir_filter/Q_data_add_3_buff_reg[4]  ( .D(n2015), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_3_buff [4]) );
  DF3 \u_decoder/fir_filter/Q_data_add_3_buff_reg[3]  ( .D(n2016), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_3_buff [3]) );
  DF3 \u_decoder/fir_filter/Q_data_add_3_buff_reg[2]  ( .D(n2017), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_3_buff [2]) );
  DF3 \u_decoder/fir_filter/Q_data_add_3_buff_reg[1]  ( .D(n2018), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_3_buff [1]) );
  DF3 \u_decoder/fir_filter/Q_data_add_3_buff_reg[0]  ( .D(n2019), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_3_buff [0]), .QN(n99) );
  DF3 \u_decoder/fir_filter/Q_data_add_4_buff_reg[14]  ( .D(n2020), .C(inClock), .Q(\u_decoder/fir_filter/Q_data_add_4_buff [14]) );
  DF3 \u_decoder/fir_filter/Q_data_add_4_buff_reg[13]  ( .D(n2021), .C(inClock), .Q(\u_decoder/fir_filter/Q_data_add_4_buff [13]) );
  DF3 \u_decoder/fir_filter/Q_data_add_4_buff_reg[12]  ( .D(n2022), .C(inClock), .Q(\u_decoder/fir_filter/Q_data_add_4_buff [12]) );
  DF3 \u_decoder/fir_filter/Q_data_add_4_buff_reg[11]  ( .D(n2023), .C(inClock), .Q(\u_decoder/fir_filter/Q_data_add_4_buff [11]) );
  DF3 \u_decoder/fir_filter/Q_data_add_4_buff_reg[10]  ( .D(n2024), .C(inClock), .Q(\u_decoder/fir_filter/Q_data_add_4_buff [10]) );
  DF3 \u_decoder/fir_filter/Q_data_add_4_buff_reg[9]  ( .D(n2025), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_4_buff [9]) );
  DF3 \u_decoder/fir_filter/Q_data_add_4_buff_reg[8]  ( .D(n2026), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_4_buff [8]) );
  DF3 \u_decoder/fir_filter/Q_data_add_4_buff_reg[7]  ( .D(n2027), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_4_buff [7]) );
  DF3 \u_decoder/fir_filter/Q_data_add_4_buff_reg[6]  ( .D(n2028), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_4_buff [6]) );
  DF3 \u_decoder/fir_filter/Q_data_add_4_buff_reg[5]  ( .D(n2029), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_4_buff [5]) );
  DF3 \u_decoder/fir_filter/Q_data_add_4_buff_reg[4]  ( .D(n2030), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_4_buff [4]) );
  DF3 \u_decoder/fir_filter/Q_data_add_4_buff_reg[3]  ( .D(n2031), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_4_buff [3]) );
  DF3 \u_decoder/fir_filter/Q_data_add_4_buff_reg[2]  ( .D(n2032), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_4_buff [2]) );
  DF3 \u_decoder/fir_filter/Q_data_add_4_buff_reg[1]  ( .D(n2033), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_4_buff [1]) );
  DF3 \u_decoder/fir_filter/Q_data_add_4_buff_reg[0]  ( .D(n2034), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_4_buff [0]), .QN(n98) );
  DF3 \u_decoder/fir_filter/Q_data_add_5_buff_reg[14]  ( .D(n2035), .C(inClock), .Q(\u_decoder/fir_filter/Q_data_add_5_buff [14]) );
  DF3 \u_decoder/fir_filter/Q_data_add_5_buff_reg[13]  ( .D(n2036), .C(inClock), .Q(\u_decoder/fir_filter/Q_data_add_5_buff [13]) );
  DF3 \u_decoder/fir_filter/Q_data_add_5_buff_reg[12]  ( .D(n2037), .C(inClock), .Q(\u_decoder/fir_filter/Q_data_add_5_buff [12]) );
  DF3 \u_decoder/fir_filter/Q_data_add_5_buff_reg[11]  ( .D(n2038), .C(inClock), .Q(\u_decoder/fir_filter/Q_data_add_5_buff [11]) );
  DF3 \u_decoder/fir_filter/Q_data_add_5_buff_reg[10]  ( .D(n2039), .C(inClock), .Q(\u_decoder/fir_filter/Q_data_add_5_buff [10]) );
  DF3 \u_decoder/fir_filter/Q_data_add_5_buff_reg[9]  ( .D(n2040), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_5_buff [9]) );
  DF3 \u_decoder/fir_filter/Q_data_add_5_buff_reg[8]  ( .D(n2041), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_5_buff [8]) );
  DF3 \u_decoder/fir_filter/Q_data_add_5_buff_reg[7]  ( .D(n2042), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_5_buff [7]) );
  DF3 \u_decoder/fir_filter/Q_data_add_5_buff_reg[6]  ( .D(n2043), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_5_buff [6]) );
  DF3 \u_decoder/fir_filter/Q_data_add_5_buff_reg[5]  ( .D(n2044), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_5_buff [5]) );
  DF3 \u_decoder/fir_filter/Q_data_add_5_buff_reg[4]  ( .D(n2045), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_5_buff [4]) );
  DF3 \u_decoder/fir_filter/Q_data_add_5_buff_reg[3]  ( .D(n2046), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_5_buff [3]) );
  DF3 \u_decoder/fir_filter/Q_data_add_5_buff_reg[2]  ( .D(n2047), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_5_buff [2]) );
  DF3 \u_decoder/fir_filter/Q_data_add_5_buff_reg[1]  ( .D(n2048), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_5_buff [1]) );
  DF3 \u_decoder/fir_filter/Q_data_add_5_buff_reg[0]  ( .D(n2049), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_5_buff [0]), .QN(n97) );
  DF3 \u_decoder/fir_filter/Q_data_add_6_buff_reg[14]  ( .D(n2050), .C(inClock), .Q(\u_decoder/fir_filter/Q_data_add_6_buff [14]) );
  DF3 \u_decoder/fir_filter/Q_data_add_6_buff_reg[13]  ( .D(n2051), .C(inClock), .Q(\u_decoder/fir_filter/Q_data_add_6_buff [13]) );
  DF3 \u_decoder/fir_filter/Q_data_add_6_buff_reg[12]  ( .D(n2052), .C(inClock), .Q(\u_decoder/fir_filter/Q_data_add_6_buff [12]) );
  DF3 \u_decoder/fir_filter/Q_data_add_6_buff_reg[11]  ( .D(n2053), .C(inClock), .Q(\u_decoder/fir_filter/Q_data_add_6_buff [11]) );
  DF3 \u_decoder/fir_filter/Q_data_add_6_buff_reg[10]  ( .D(n2054), .C(inClock), .Q(\u_decoder/fir_filter/Q_data_add_6_buff [10]) );
  DF3 \u_decoder/fir_filter/Q_data_add_6_buff_reg[9]  ( .D(n2055), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_6_buff [9]) );
  DF3 \u_decoder/fir_filter/Q_data_add_6_buff_reg[8]  ( .D(n2056), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_6_buff [8]) );
  DF3 \u_decoder/fir_filter/Q_data_add_6_buff_reg[7]  ( .D(n2057), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_6_buff [7]) );
  DF3 \u_decoder/fir_filter/Q_data_add_6_buff_reg[6]  ( .D(n2058), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_6_buff [6]) );
  DF3 \u_decoder/fir_filter/Q_data_add_6_buff_reg[5]  ( .D(n2059), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_6_buff [5]) );
  DF3 \u_decoder/fir_filter/Q_data_add_6_buff_reg[4]  ( .D(n2060), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_6_buff [4]) );
  DF3 \u_decoder/fir_filter/Q_data_add_6_buff_reg[3]  ( .D(n2061), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_6_buff [3]) );
  DF3 \u_decoder/fir_filter/Q_data_add_6_buff_reg[2]  ( .D(n2062), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_6_buff [2]) );
  DF3 \u_decoder/fir_filter/Q_data_add_6_buff_reg[1]  ( .D(n2063), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_6_buff [1]) );
  DF3 \u_decoder/fir_filter/Q_data_add_6_buff_reg[0]  ( .D(n2064), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_6_buff [0]), .QN(n96) );
  DF3 \u_decoder/fir_filter/Q_data_add_7_buff_reg[14]  ( .D(n2065), .C(inClock), .Q(\u_decoder/fir_filter/Q_data_add_7_buff [14]) );
  DF3 \u_decoder/fir_filter/Q_data_add_7_buff_reg[13]  ( .D(n2066), .C(inClock), .Q(\u_decoder/fir_filter/Q_data_add_7_buff [13]) );
  DF3 \u_decoder/fir_filter/Q_data_add_7_buff_reg[12]  ( .D(n2067), .C(inClock), .Q(\u_decoder/fir_filter/Q_data_add_7_buff [12]) );
  DF3 \u_decoder/fir_filter/Q_data_add_7_buff_reg[11]  ( .D(n2068), .C(inClock), .Q(\u_decoder/fir_filter/Q_data_add_7_buff [11]) );
  DF3 \u_decoder/fir_filter/Q_data_add_7_buff_reg[10]  ( .D(n2069), .C(inClock), .Q(\u_decoder/fir_filter/Q_data_add_7_buff [10]) );
  DF3 \u_decoder/fir_filter/Q_data_add_7_buff_reg[9]  ( .D(n2070), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_7_buff [9]) );
  DF3 \u_decoder/fir_filter/Q_data_add_7_buff_reg[8]  ( .D(n2071), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_7_buff [8]) );
  DF3 \u_decoder/fir_filter/Q_data_add_7_buff_reg[7]  ( .D(n2072), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_7_buff [7]) );
  DF3 \u_decoder/fir_filter/Q_data_add_7_buff_reg[6]  ( .D(n2073), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_7_buff [6]) );
  DF3 \u_decoder/fir_filter/Q_data_add_7_buff_reg[5]  ( .D(n2074), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_7_buff [5]) );
  DF3 \u_decoder/fir_filter/Q_data_add_7_buff_reg[4]  ( .D(n2075), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_7_buff [4]) );
  DF3 \u_decoder/fir_filter/Q_data_add_7_buff_reg[3]  ( .D(n2076), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_7_buff [3]) );
  DF3 \u_decoder/fir_filter/Q_data_add_7_buff_reg[2]  ( .D(n2077), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_7_buff [2]) );
  DF3 \u_decoder/fir_filter/Q_data_add_7_buff_reg[1]  ( .D(n2078), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_7_buff [1]) );
  DF3 \u_decoder/fir_filter/Q_data_add_7_buff_reg[0]  ( .D(n2079), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_7_buff [0]), .QN(n95) );
  DF3 \u_decoder/fir_filter/Q_data_mult_8_buff_reg[0]  ( .D(
        \u_decoder/fir_filter/n1155 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_8_buff [0]), .QN(n88) );
  DF3 \u_decoder/fir_filter/Q_data_mult_8_buff_reg[1]  ( .D(
        \u_decoder/fir_filter/n1156 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_8_buff [1]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_8_buff_reg[2]  ( .D(
        \u_decoder/fir_filter/n1157 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_8_buff [2]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_8_buff_reg[3]  ( .D(
        \u_decoder/fir_filter/n1158 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_8_buff [3]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_8_buff_reg[4]  ( .D(
        \u_decoder/fir_filter/n1159 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_8_buff [4]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_8_buff_reg[5]  ( .D(
        \u_decoder/fir_filter/n1160 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_8_buff [5]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_8_buff_reg[6]  ( .D(
        \u_decoder/fir_filter/n1161 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_8_buff [6]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_8_buff_reg[7]  ( .D(
        \u_decoder/fir_filter/n1162 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_8_buff [7]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_8_buff_reg[8]  ( .D(
        \u_decoder/fir_filter/n1163 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_8_buff [8]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_8_buff_reg[9]  ( .D(
        \u_decoder/fir_filter/n1164 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_8_buff [9]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_8_buff_reg[10]  ( .D(
        \u_decoder/fir_filter/n1165 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_8_buff [10]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_8_buff_reg[11]  ( .D(
        \u_decoder/fir_filter/n1166 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_8_buff [11]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_8_buff_reg[12]  ( .D(
        \u_decoder/fir_filter/n1167 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_8_buff [12]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_8_buff_reg[13]  ( .D(
        \u_decoder/fir_filter/n1168 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_8_buff [13]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_8_buff_reg[14]  ( .D(
        \u_decoder/fir_filter/n1169 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_8_buff [14]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_8_delay_reg[0]  ( .D(
        \u_decoder/fir_filter/n1176 ), .C(inClock), .QN(
        \u_decoder/fir_filter/n442 ) );
  DF3 \u_decoder/fir_filter/Q_data_mult_8_delay_reg[1]  ( .D(
        \u_decoder/fir_filter/n1177 ), .C(inClock), .QN(
        \u_decoder/fir_filter/n441 ) );
  DF3 \u_decoder/fir_filter/Q_data_mult_8_delay_reg[2]  ( .D(
        \u_decoder/fir_filter/n1178 ), .C(inClock), .QN(
        \u_decoder/fir_filter/n440 ) );
  DF3 \u_decoder/fir_filter/Q_data_mult_8_delay_reg[3]  ( .D(
        \u_decoder/fir_filter/n1179 ), .C(inClock), .QN(
        \u_decoder/fir_filter/n439 ) );
  DF3 \u_decoder/fir_filter/Q_data_mult_8_delay_reg[4]  ( .D(
        \u_decoder/fir_filter/n1180 ), .C(inClock), .QN(
        \u_decoder/fir_filter/n438 ) );
  DF3 \u_decoder/fir_filter/Q_data_mult_8_delay_reg[5]  ( .D(
        \u_decoder/fir_filter/n1181 ), .C(inClock), .QN(
        \u_decoder/fir_filter/n437 ) );
  DF3 \u_decoder/fir_filter/Q_data_mult_8_delay_reg[6]  ( .D(
        \u_decoder/fir_filter/n1182 ), .C(inClock), .QN(
        \u_decoder/fir_filter/n436 ) );
  DF3 \u_decoder/fir_filter/Q_data_mult_8_delay_reg[7]  ( .D(
        \u_decoder/fir_filter/n1183 ), .C(inClock), .QN(
        \u_decoder/fir_filter/n435 ) );
  DF3 \u_decoder/fir_filter/Q_data_mult_8_delay_reg[8]  ( .D(
        \u_decoder/fir_filter/n1184 ), .C(inClock), .QN(
        \u_decoder/fir_filter/n434 ) );
  DF3 \u_decoder/fir_filter/Q_data_mult_8_delay_reg[9]  ( .D(
        \u_decoder/fir_filter/n1185 ), .C(inClock), .QN(
        \u_decoder/fir_filter/n433 ) );
  DF3 \u_decoder/fir_filter/Q_data_mult_8_delay_reg[10]  ( .D(
        \u_decoder/fir_filter/n1186 ), .C(inClock), .QN(
        \u_decoder/fir_filter/n432 ) );
  DF3 \u_decoder/fir_filter/Q_data_mult_8_delay_reg[11]  ( .D(
        \u_decoder/fir_filter/n1187 ), .C(inClock), .QN(
        \u_decoder/fir_filter/n431 ) );
  DF3 \u_decoder/fir_filter/Q_data_mult_8_delay_reg[12]  ( .D(
        \u_decoder/fir_filter/n1188 ), .C(inClock), .QN(
        \u_decoder/fir_filter/n430 ) );
  DF3 \u_decoder/fir_filter/Q_data_mult_8_delay_reg[13]  ( .D(
        \u_decoder/fir_filter/n1189 ), .C(inClock), .QN(
        \u_decoder/fir_filter/n429 ) );
  DF3 \u_decoder/fir_filter/Q_data_mult_8_delay_reg[14]  ( .D(
        \u_decoder/fir_filter/n1190 ), .C(inClock), .QN(
        \u_decoder/fir_filter/n428 ) );
  DF3 \u_decoder/fir_filter/Q_data_mult_7_buff_reg[0]  ( .D(
        \u_decoder/fir_filter/n1192 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_7_buff [0]), .QN(n10) );
  DF3 \u_decoder/fir_filter/Q_data_mult_7_buff_reg[1]  ( .D(
        \u_decoder/fir_filter/n1193 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_7_buff [1]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_7_buff_reg[2]  ( .D(
        \u_decoder/fir_filter/n1194 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_7_buff [2]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_7_buff_reg[3]  ( .D(
        \u_decoder/fir_filter/n1195 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_7_buff [3]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_7_buff_reg[4]  ( .D(
        \u_decoder/fir_filter/n1196 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_7_buff [4]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_7_buff_reg[5]  ( .D(
        \u_decoder/fir_filter/n1197 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_7_buff [5]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_7_buff_reg[6]  ( .D(
        \u_decoder/fir_filter/n1198 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_7_buff [6]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_7_buff_reg[7]  ( .D(
        \u_decoder/fir_filter/n1199 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_7_buff [7]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_7_buff_reg[8]  ( .D(
        \u_decoder/fir_filter/n1200 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_7_buff [8]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_7_buff_reg[9]  ( .D(
        \u_decoder/fir_filter/n1201 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_7_buff [9]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_7_buff_reg[10]  ( .D(
        \u_decoder/fir_filter/n1202 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_7_buff [10]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_7_buff_reg[11]  ( .D(
        \u_decoder/fir_filter/n1203 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_7_buff [11]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_7_buff_reg[12]  ( .D(
        \u_decoder/fir_filter/n1204 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_7_buff [12]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_7_buff_reg[13]  ( .D(
        \u_decoder/fir_filter/n1205 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_7_buff [13]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_7_buff_reg[14]  ( .D(
        \u_decoder/fir_filter/n1206 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_7_buff [14]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_6_buff_reg[0]  ( .D(n2080), .C(inClock), .Q(\u_decoder/fir_filter/Q_data_mult_6_buff [0]), .QN(n16) );
  DF3 \u_decoder/fir_filter/Q_data_mult_6_buff_reg[1]  ( .D(
        \u_decoder/fir_filter/n1209 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_6_buff [1]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_6_buff_reg[2]  ( .D(
        \u_decoder/fir_filter/n1210 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_6_buff [2]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_6_buff_reg[3]  ( .D(
        \u_decoder/fir_filter/n1211 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_6_buff [3]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_6_buff_reg[4]  ( .D(
        \u_decoder/fir_filter/n1212 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_6_buff [4]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_6_buff_reg[5]  ( .D(
        \u_decoder/fir_filter/n1213 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_6_buff [5]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_6_buff_reg[6]  ( .D(
        \u_decoder/fir_filter/n1214 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_6_buff [6]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_6_buff_reg[7]  ( .D(
        \u_decoder/fir_filter/n1215 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_6_buff [7]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_6_buff_reg[8]  ( .D(
        \u_decoder/fir_filter/n1216 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_6_buff [8]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_6_buff_reg[9]  ( .D(
        \u_decoder/fir_filter/n1217 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_6_buff [9]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_6_buff_reg[10]  ( .D(
        \u_decoder/fir_filter/n1218 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_6_buff [10]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_6_buff_reg[11]  ( .D(
        \u_decoder/fir_filter/n1219 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_6_buff [11]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_6_buff_reg[12]  ( .D(
        \u_decoder/fir_filter/n1220 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_6_buff [12]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_6_buff_reg[13]  ( .D(
        \u_decoder/fir_filter/n1221 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_6_buff [13]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_6_buff_reg[14]  ( .D(
        \u_decoder/fir_filter/n1222 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_6_buff [14]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_5_buff_reg[0]  ( .D(
        \u_decoder/fir_filter/n1224 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_5_buff [0]), .QN(n17) );
  DF3 \u_decoder/fir_filter/Q_data_mult_5_buff_reg[1]  ( .D(
        \u_decoder/fir_filter/n1225 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_5_buff [1]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_5_buff_reg[2]  ( .D(
        \u_decoder/fir_filter/n1226 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_5_buff [2]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_5_buff_reg[3]  ( .D(
        \u_decoder/fir_filter/n1227 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_5_buff [3]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_5_buff_reg[4]  ( .D(
        \u_decoder/fir_filter/n1228 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_5_buff [4]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_5_buff_reg[5]  ( .D(
        \u_decoder/fir_filter/n1229 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_5_buff [5]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_5_buff_reg[6]  ( .D(
        \u_decoder/fir_filter/n1230 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_5_buff [6]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_5_buff_reg[7]  ( .D(
        \u_decoder/fir_filter/n1231 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_5_buff [7]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_5_buff_reg[8]  ( .D(
        \u_decoder/fir_filter/n1232 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_5_buff [8]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_5_buff_reg[9]  ( .D(
        \u_decoder/fir_filter/n1233 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_5_buff [9]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_5_buff_reg[10]  ( .D(
        \u_decoder/fir_filter/n1234 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_5_buff [10]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_5_buff_reg[11]  ( .D(
        \u_decoder/fir_filter/n1235 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_5_buff [11]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_5_buff_reg[12]  ( .D(
        \u_decoder/fir_filter/n1236 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_5_buff [12]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_5_buff_reg[13]  ( .D(
        \u_decoder/fir_filter/n1237 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_5_buff [13]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_5_buff_reg[14]  ( .D(
        \u_decoder/fir_filter/n1238 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_5_buff [14]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_4_buff_reg[0]  ( .D(n1889), .C(inClock), .Q(\u_decoder/fir_filter/Q_data_mult_4_buff [0]), .QN(n22) );
  DF3 \u_decoder/fir_filter/Q_data_mult_4_buff_reg[1]  ( .D(n1932), .C(inClock), .Q(\u_decoder/fir_filter/Q_data_mult_4_buff [1]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_4_buff_reg[2]  ( .D(n1934), .C(inClock), .Q(\u_decoder/fir_filter/Q_data_mult_4_buff [2]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_4_buff_reg[3]  ( .D(n1907), .C(inClock), .Q(\u_decoder/fir_filter/Q_data_mult_4_buff [3]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_4_buff_reg[4]  ( .D(n1906), .C(inClock), .Q(\u_decoder/fir_filter/Q_data_mult_4_buff [4]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_4_buff_reg[5]  ( .D(n1905), .C(inClock), .Q(\u_decoder/fir_filter/Q_data_mult_4_buff [5]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_4_buff_reg[6]  ( .D(n1904), .C(inClock), .Q(\u_decoder/fir_filter/Q_data_mult_4_buff [6]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_4_buff_reg[7]  ( .D(n1903), .C(inClock), .Q(\u_decoder/fir_filter/Q_data_mult_4_buff [7]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_4_buff_reg[8]  ( .D(n1902), .C(inClock), .Q(\u_decoder/fir_filter/Q_data_mult_4_buff [8]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_4_buff_reg[9]  ( .D(n1901), .C(inClock), .Q(\u_decoder/fir_filter/Q_data_mult_4_buff [9]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_4_buff_reg[10]  ( .D(n1899), .C(
        inClock), .Q(\u_decoder/fir_filter/Q_data_mult_4_buff [10]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_4_buff_reg[11]  ( .D(n1895), .C(
        inClock), .Q(\u_decoder/fir_filter/Q_data_mult_4_buff [11]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_4_buff_reg[12]  ( .D(n1890), .C(
        inClock), .Q(\u_decoder/fir_filter/Q_data_mult_4_buff [12]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_4_buff_reg[13]  ( .D(n1892), .C(
        inClock), .Q(\u_decoder/fir_filter/Q_data_mult_4_buff [13]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_4_buff_reg[14]  ( .D(n1893), .C(
        inClock), .Q(\u_decoder/fir_filter/Q_data_mult_4_buff [14]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_3_buff_reg[0]  ( .D(
        \u_decoder/fir_filter/n1240 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_3_buff [0]), .QN(n18) );
  DF3 \u_decoder/fir_filter/Q_data_mult_3_buff_reg[1]  ( .D(
        \u_decoder/fir_filter/n1241 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_3_buff [1]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_3_buff_reg[2]  ( .D(
        \u_decoder/fir_filter/n1242 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_3_buff [2]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_3_buff_reg[3]  ( .D(
        \u_decoder/fir_filter/n1243 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_3_buff [3]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_3_buff_reg[4]  ( .D(
        \u_decoder/fir_filter/n1244 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_3_buff [4]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_3_buff_reg[5]  ( .D(
        \u_decoder/fir_filter/n1245 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_3_buff [5]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_3_buff_reg[6]  ( .D(
        \u_decoder/fir_filter/n1246 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_3_buff [6]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_3_buff_reg[7]  ( .D(
        \u_decoder/fir_filter/n1247 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_3_buff [7]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_3_buff_reg[8]  ( .D(
        \u_decoder/fir_filter/n1248 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_3_buff [8]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_3_buff_reg[9]  ( .D(
        \u_decoder/fir_filter/n1249 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_3_buff [9]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_3_buff_reg[10]  ( .D(
        \u_decoder/fir_filter/n1250 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_3_buff [10]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_3_buff_reg[11]  ( .D(
        \u_decoder/fir_filter/n1251 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_3_buff [11]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_3_buff_reg[12]  ( .D(
        \u_decoder/fir_filter/n1252 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_3_buff [12]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_3_buff_reg[13]  ( .D(
        \u_decoder/fir_filter/n1253 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_3_buff [13]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_3_buff_reg[14]  ( .D(
        \u_decoder/fir_filter/n1254 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_3_buff [14]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_2_buff_reg[0]  ( .D(n2081), .C(inClock), .Q(\u_decoder/fir_filter/Q_data_mult_2_buff [0]), .QN(n19) );
  DF3 \u_decoder/fir_filter/Q_data_mult_2_buff_reg[1]  ( .D(
        \u_decoder/fir_filter/n1257 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_2_buff [1]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_2_buff_reg[2]  ( .D(
        \u_decoder/fir_filter/n1258 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_2_buff [2]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_2_buff_reg[3]  ( .D(
        \u_decoder/fir_filter/n1259 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_2_buff [3]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_2_buff_reg[4]  ( .D(
        \u_decoder/fir_filter/n1260 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_2_buff [4]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_2_buff_reg[5]  ( .D(
        \u_decoder/fir_filter/n1261 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_2_buff [5]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_2_buff_reg[6]  ( .D(
        \u_decoder/fir_filter/n1262 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_2_buff [6]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_2_buff_reg[7]  ( .D(
        \u_decoder/fir_filter/n1263 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_2_buff [7]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_2_buff_reg[8]  ( .D(
        \u_decoder/fir_filter/n1264 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_2_buff [8]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_2_buff_reg[9]  ( .D(
        \u_decoder/fir_filter/n1265 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_2_buff [9]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_2_buff_reg[10]  ( .D(
        \u_decoder/fir_filter/n1266 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_2_buff [10]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_2_buff_reg[11]  ( .D(
        \u_decoder/fir_filter/n1267 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_2_buff [11]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_2_buff_reg[12]  ( .D(
        \u_decoder/fir_filter/n1268 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_2_buff [12]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_2_buff_reg[13]  ( .D(
        \u_decoder/fir_filter/n1269 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_2_buff [13]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_2_buff_reg[14]  ( .D(
        \u_decoder/fir_filter/n1270 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_2_buff [14]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_1_buff_reg[0]  ( .D(
        \u_decoder/fir_filter/n1272 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_1_buff [0]), .QN(n20) );
  DF3 \u_decoder/fir_filter/Q_data_mult_1_buff_reg[1]  ( .D(
        \u_decoder/fir_filter/n1273 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_1_buff [1]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_1_buff_reg[2]  ( .D(
        \u_decoder/fir_filter/n1274 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_1_buff [2]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_1_buff_reg[3]  ( .D(
        \u_decoder/fir_filter/n1275 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_1_buff [3]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_1_buff_reg[4]  ( .D(
        \u_decoder/fir_filter/n1276 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_1_buff [4]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_1_buff_reg[5]  ( .D(
        \u_decoder/fir_filter/n1277 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_1_buff [5]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_1_buff_reg[6]  ( .D(
        \u_decoder/fir_filter/n1278 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_1_buff [6]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_1_buff_reg[7]  ( .D(
        \u_decoder/fir_filter/n1279 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_1_buff [7]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_1_buff_reg[8]  ( .D(
        \u_decoder/fir_filter/n1280 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_1_buff [8]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_1_buff_reg[9]  ( .D(
        \u_decoder/fir_filter/n1281 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_1_buff [9]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_1_buff_reg[10]  ( .D(
        \u_decoder/fir_filter/n1282 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_1_buff [10]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_1_buff_reg[11]  ( .D(
        \u_decoder/fir_filter/n1283 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_1_buff [11]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_1_buff_reg[12]  ( .D(
        \u_decoder/fir_filter/n1284 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_1_buff [12]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_1_buff_reg[13]  ( .D(
        \u_decoder/fir_filter/n1285 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_1_buff [13]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_1_buff_reg[14]  ( .D(
        \u_decoder/fir_filter/n1286 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_1_buff [14]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_0_buff_reg[0]  ( .D(
        \u_decoder/fir_filter/n1288 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_0_buff [0]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_0_buff_reg[1]  ( .D(
        \u_decoder/fir_filter/n1289 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_0_buff [1]), .QN(n73) );
  DF3 \u_decoder/fir_filter/Q_data_mult_0_buff_reg[2]  ( .D(
        \u_decoder/fir_filter/n1290 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_0_buff [2]), .QN(n71) );
  DF3 \u_decoder/fir_filter/Q_data_mult_0_buff_reg[3]  ( .D(
        \u_decoder/fir_filter/n1291 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_0_buff [3]), .QN(n112) );
  DF3 \u_decoder/fir_filter/Q_data_mult_0_buff_reg[4]  ( .D(
        \u_decoder/fir_filter/n1292 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_0_buff [4]), .QN(n128) );
  DF3 \u_decoder/fir_filter/Q_data_mult_0_buff_reg[5]  ( .D(
        \u_decoder/fir_filter/n1293 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_0_buff [5]), .QN(n129) );
  DF3 \u_decoder/fir_filter/Q_data_mult_0_buff_reg[6]  ( .D(
        \u_decoder/fir_filter/n1294 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_0_buff [6]), .QN(n142) );
  DF3 \u_decoder/fir_filter/Q_data_mult_0_buff_reg[7]  ( .D(
        \u_decoder/fir_filter/n1295 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_0_buff [7]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_0_buff_reg[8]  ( .D(
        \u_decoder/fir_filter/n1296 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_0_buff [8]), .QN(n198) );
  DF3 \u_decoder/fir_filter/Q_data_mult_0_buff_reg[9]  ( .D(
        \u_decoder/fir_filter/n1297 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_0_buff [9]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_0_buff_reg[10]  ( .D(
        \u_decoder/fir_filter/n1298 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_0_buff [10]), .QN(n258) );
  DF3 \u_decoder/fir_filter/Q_data_mult_0_buff_reg[11]  ( .D(
        \u_decoder/fir_filter/n1299 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_0_buff [11]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_0_buff_reg[12]  ( .D(
        \u_decoder/fir_filter/n1300 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_0_buff [12]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_0_buff_reg[13]  ( .D(
        \u_decoder/fir_filter/n1301 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_0_buff [13]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_0_buff_reg[14]  ( .D(
        \u_decoder/fir_filter/n1302 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_0_buff [14]) );
  DF3 \u_decoder/fir_filter/o_I_postfilter_reg[3]  ( .D(n2082), .C(inClock), 
        .Q(sig_decod_outI[3]) );
  DF3 \u_decoder/fir_filter/o_I_postfilter_reg[2]  ( .D(n2083), .C(inClock), 
        .Q(sig_decod_outI[2]) );
  DF3 \u_decoder/fir_filter/o_I_postfilter_reg[1]  ( .D(n2084), .C(inClock), 
        .Q(sig_decod_outI[1]) );
  DF3 \u_decoder/fir_filter/o_I_postfilter_reg[0]  ( .D(n2085), .C(inClock), 
        .Q(sig_decod_outI[0]) );
  DF3 \u_decoder/fir_filter/I_data_add_1_buff_reg[14]  ( .D(n2086), .C(inClock), .Q(\u_decoder/fir_filter/I_data_add_1_buff [14]) );
  DF3 \u_decoder/fir_filter/I_data_add_1_buff_reg[13]  ( .D(n2087), .C(inClock), .Q(\u_decoder/fir_filter/I_data_add_1_buff [13]) );
  DF3 \u_decoder/fir_filter/I_data_add_1_buff_reg[12]  ( .D(n2088), .C(inClock), .Q(\u_decoder/fir_filter/I_data_add_1_buff [12]) );
  DF3 \u_decoder/fir_filter/I_data_add_1_buff_reg[11]  ( .D(n2089), .C(inClock), .Q(\u_decoder/fir_filter/I_data_add_1_buff [11]) );
  DF3 \u_decoder/fir_filter/I_data_add_1_buff_reg[10]  ( .D(n2090), .C(inClock), .Q(\u_decoder/fir_filter/I_data_add_1_buff [10]) );
  DF3 \u_decoder/fir_filter/I_data_add_1_buff_reg[9]  ( .D(n2093), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_1_buff [9]) );
  DF3 \u_decoder/fir_filter/I_data_add_1_buff_reg[8]  ( .D(n2094), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_1_buff [8]) );
  DF3 \u_decoder/fir_filter/I_data_add_1_buff_reg[7]  ( .D(n2097), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_1_buff [7]) );
  DF3 \u_decoder/fir_filter/I_data_add_1_buff_reg[6]  ( .D(n2098), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_1_buff [6]) );
  DF3 \u_decoder/fir_filter/I_data_add_1_buff_reg[5]  ( .D(n2100), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_1_buff [5]) );
  DF3 \u_decoder/fir_filter/I_data_add_1_buff_reg[4]  ( .D(n2102), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_1_buff [4]) );
  DF3 \u_decoder/fir_filter/I_data_add_1_buff_reg[3]  ( .D(n2104), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_1_buff [3]) );
  DF3 \u_decoder/fir_filter/I_data_add_1_buff_reg[2]  ( .D(n2106), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_1_buff [2]) );
  DF3 \u_decoder/fir_filter/I_data_add_1_buff_reg[1]  ( .D(n2108), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_1_buff [1]), .QN(n8) );
  DF3 \u_decoder/fir_filter/I_data_add_1_buff_reg[0]  ( .D(n2109), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_1_buff [0]) );
  DF3 \u_decoder/fir_filter/I_data_add_2_buff_reg[14]  ( .D(n2110), .C(inClock), .Q(\u_decoder/fir_filter/I_data_add_2_buff [14]) );
  DF3 \u_decoder/fir_filter/I_data_add_2_buff_reg[13]  ( .D(n2111), .C(inClock), .Q(\u_decoder/fir_filter/I_data_add_2_buff [13]) );
  DF3 \u_decoder/fir_filter/I_data_add_2_buff_reg[12]  ( .D(n2112), .C(inClock), .Q(\u_decoder/fir_filter/I_data_add_2_buff [12]) );
  DF3 \u_decoder/fir_filter/I_data_add_2_buff_reg[11]  ( .D(n2113), .C(inClock), .Q(\u_decoder/fir_filter/I_data_add_2_buff [11]) );
  DF3 \u_decoder/fir_filter/I_data_add_2_buff_reg[10]  ( .D(n2114), .C(inClock), .Q(\u_decoder/fir_filter/I_data_add_2_buff [10]) );
  DF3 \u_decoder/fir_filter/I_data_add_2_buff_reg[9]  ( .D(n2115), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_2_buff [9]) );
  DF3 \u_decoder/fir_filter/I_data_add_2_buff_reg[8]  ( .D(n2116), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_2_buff [8]) );
  DF3 \u_decoder/fir_filter/I_data_add_2_buff_reg[7]  ( .D(n2117), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_2_buff [7]) );
  DF3 \u_decoder/fir_filter/I_data_add_2_buff_reg[6]  ( .D(n2118), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_2_buff [6]) );
  DF3 \u_decoder/fir_filter/I_data_add_2_buff_reg[5]  ( .D(n2119), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_2_buff [5]) );
  DF3 \u_decoder/fir_filter/I_data_add_2_buff_reg[4]  ( .D(n2120), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_2_buff [4]) );
  DF3 \u_decoder/fir_filter/I_data_add_2_buff_reg[3]  ( .D(n2121), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_2_buff [3]) );
  DF3 \u_decoder/fir_filter/I_data_add_2_buff_reg[2]  ( .D(n2122), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_2_buff [2]) );
  DF3 \u_decoder/fir_filter/I_data_add_2_buff_reg[1]  ( .D(n2123), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_2_buff [1]) );
  DF3 \u_decoder/fir_filter/I_data_add_2_buff_reg[0]  ( .D(n2124), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_2_buff [0]), .QN(n94) );
  DF3 \u_decoder/fir_filter/I_data_add_3_buff_reg[14]  ( .D(n2125), .C(inClock), .Q(\u_decoder/fir_filter/I_data_add_3_buff [14]) );
  DF3 \u_decoder/fir_filter/I_data_add_3_buff_reg[13]  ( .D(n2126), .C(inClock), .Q(\u_decoder/fir_filter/I_data_add_3_buff [13]) );
  DF3 \u_decoder/fir_filter/I_data_add_3_buff_reg[12]  ( .D(n2127), .C(inClock), .Q(\u_decoder/fir_filter/I_data_add_3_buff [12]) );
  DF3 \u_decoder/fir_filter/I_data_add_3_buff_reg[11]  ( .D(n2128), .C(inClock), .Q(\u_decoder/fir_filter/I_data_add_3_buff [11]) );
  DF3 \u_decoder/fir_filter/I_data_add_3_buff_reg[10]  ( .D(n2129), .C(inClock), .Q(\u_decoder/fir_filter/I_data_add_3_buff [10]) );
  DF3 \u_decoder/fir_filter/I_data_add_3_buff_reg[9]  ( .D(n2130), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_3_buff [9]) );
  DF3 \u_decoder/fir_filter/I_data_add_3_buff_reg[8]  ( .D(n2131), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_3_buff [8]) );
  DF3 \u_decoder/fir_filter/I_data_add_3_buff_reg[7]  ( .D(n2132), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_3_buff [7]) );
  DF3 \u_decoder/fir_filter/I_data_add_3_buff_reg[6]  ( .D(n2133), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_3_buff [6]) );
  DF3 \u_decoder/fir_filter/I_data_add_3_buff_reg[5]  ( .D(n2134), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_3_buff [5]) );
  DF3 \u_decoder/fir_filter/I_data_add_3_buff_reg[4]  ( .D(n2135), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_3_buff [4]) );
  DF3 \u_decoder/fir_filter/I_data_add_3_buff_reg[3]  ( .D(n2136), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_3_buff [3]) );
  DF3 \u_decoder/fir_filter/I_data_add_3_buff_reg[2]  ( .D(n2137), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_3_buff [2]) );
  DF3 \u_decoder/fir_filter/I_data_add_3_buff_reg[1]  ( .D(n2138), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_3_buff [1]) );
  DF3 \u_decoder/fir_filter/I_data_add_3_buff_reg[0]  ( .D(n2139), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_3_buff [0]), .QN(n93) );
  DF3 \u_decoder/fir_filter/I_data_add_4_buff_reg[14]  ( .D(n2140), .C(inClock), .Q(\u_decoder/fir_filter/I_data_add_4_buff [14]) );
  DF3 \u_decoder/fir_filter/I_data_add_4_buff_reg[13]  ( .D(n2141), .C(inClock), .Q(\u_decoder/fir_filter/I_data_add_4_buff [13]) );
  DF3 \u_decoder/fir_filter/I_data_add_4_buff_reg[12]  ( .D(n2142), .C(inClock), .Q(\u_decoder/fir_filter/I_data_add_4_buff [12]) );
  DF3 \u_decoder/fir_filter/I_data_add_4_buff_reg[11]  ( .D(n2143), .C(inClock), .Q(\u_decoder/fir_filter/I_data_add_4_buff [11]) );
  DF3 \u_decoder/fir_filter/I_data_add_4_buff_reg[10]  ( .D(n2144), .C(inClock), .Q(\u_decoder/fir_filter/I_data_add_4_buff [10]) );
  DF3 \u_decoder/fir_filter/I_data_add_4_buff_reg[9]  ( .D(n2145), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_4_buff [9]) );
  DF3 \u_decoder/fir_filter/I_data_add_4_buff_reg[8]  ( .D(n2146), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_4_buff [8]) );
  DF3 \u_decoder/fir_filter/I_data_add_4_buff_reg[7]  ( .D(n2147), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_4_buff [7]) );
  DF3 \u_decoder/fir_filter/I_data_add_4_buff_reg[6]  ( .D(n2148), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_4_buff [6]) );
  DF3 \u_decoder/fir_filter/I_data_add_4_buff_reg[5]  ( .D(n2149), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_4_buff [5]) );
  DF3 \u_decoder/fir_filter/I_data_add_4_buff_reg[4]  ( .D(n2150), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_4_buff [4]) );
  DF3 \u_decoder/fir_filter/I_data_add_4_buff_reg[3]  ( .D(n2151), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_4_buff [3]) );
  DF3 \u_decoder/fir_filter/I_data_add_4_buff_reg[2]  ( .D(n2152), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_4_buff [2]) );
  DF3 \u_decoder/fir_filter/I_data_add_4_buff_reg[1]  ( .D(n2153), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_4_buff [1]) );
  DF3 \u_decoder/fir_filter/I_data_add_4_buff_reg[0]  ( .D(n2154), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_4_buff [0]), .QN(n92) );
  DF3 \u_decoder/fir_filter/I_data_add_5_buff_reg[14]  ( .D(n2155), .C(inClock), .Q(\u_decoder/fir_filter/I_data_add_5_buff [14]) );
  DF3 \u_decoder/fir_filter/I_data_add_5_buff_reg[13]  ( .D(n2156), .C(inClock), .Q(\u_decoder/fir_filter/I_data_add_5_buff [13]) );
  DF3 \u_decoder/fir_filter/I_data_add_5_buff_reg[12]  ( .D(n2157), .C(inClock), .Q(\u_decoder/fir_filter/I_data_add_5_buff [12]) );
  DF3 \u_decoder/fir_filter/I_data_add_5_buff_reg[11]  ( .D(n2158), .C(inClock), .Q(\u_decoder/fir_filter/I_data_add_5_buff [11]) );
  DF3 \u_decoder/fir_filter/I_data_add_5_buff_reg[10]  ( .D(n2159), .C(inClock), .Q(\u_decoder/fir_filter/I_data_add_5_buff [10]) );
  DF3 \u_decoder/fir_filter/I_data_add_5_buff_reg[9]  ( .D(n2160), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_5_buff [9]) );
  DF3 \u_decoder/fir_filter/I_data_add_5_buff_reg[8]  ( .D(n2161), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_5_buff [8]) );
  DF3 \u_decoder/fir_filter/I_data_add_5_buff_reg[7]  ( .D(n2162), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_5_buff [7]) );
  DF3 \u_decoder/fir_filter/I_data_add_5_buff_reg[6]  ( .D(n2163), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_5_buff [6]) );
  DF3 \u_decoder/fir_filter/I_data_add_5_buff_reg[5]  ( .D(n2164), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_5_buff [5]) );
  DF3 \u_decoder/fir_filter/I_data_add_5_buff_reg[4]  ( .D(n2165), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_5_buff [4]) );
  DF3 \u_decoder/fir_filter/I_data_add_5_buff_reg[3]  ( .D(n2166), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_5_buff [3]) );
  DF3 \u_decoder/fir_filter/I_data_add_5_buff_reg[2]  ( .D(n2167), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_5_buff [2]) );
  DF3 \u_decoder/fir_filter/I_data_add_5_buff_reg[1]  ( .D(n2168), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_5_buff [1]) );
  DF3 \u_decoder/fir_filter/I_data_add_5_buff_reg[0]  ( .D(n2169), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_5_buff [0]), .QN(n91) );
  DF3 \u_decoder/fir_filter/I_data_add_6_buff_reg[14]  ( .D(n2170), .C(inClock), .Q(\u_decoder/fir_filter/I_data_add_6_buff [14]) );
  DF3 \u_decoder/fir_filter/I_data_add_6_buff_reg[13]  ( .D(n2171), .C(inClock), .Q(\u_decoder/fir_filter/I_data_add_6_buff [13]) );
  DF3 \u_decoder/fir_filter/I_data_add_6_buff_reg[12]  ( .D(n2172), .C(inClock), .Q(\u_decoder/fir_filter/I_data_add_6_buff [12]) );
  DF3 \u_decoder/fir_filter/I_data_add_6_buff_reg[11]  ( .D(n2173), .C(inClock), .Q(\u_decoder/fir_filter/I_data_add_6_buff [11]) );
  DF3 \u_decoder/fir_filter/I_data_add_6_buff_reg[10]  ( .D(n2174), .C(inClock), .Q(\u_decoder/fir_filter/I_data_add_6_buff [10]) );
  DF3 \u_decoder/fir_filter/I_data_add_6_buff_reg[9]  ( .D(n2175), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_6_buff [9]) );
  DF3 \u_decoder/fir_filter/I_data_add_6_buff_reg[8]  ( .D(n2176), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_6_buff [8]) );
  DF3 \u_decoder/fir_filter/I_data_add_6_buff_reg[7]  ( .D(n2177), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_6_buff [7]) );
  DF3 \u_decoder/fir_filter/I_data_add_6_buff_reg[6]  ( .D(n2178), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_6_buff [6]) );
  DF3 \u_decoder/fir_filter/I_data_add_6_buff_reg[5]  ( .D(n2179), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_6_buff [5]) );
  DF3 \u_decoder/fir_filter/I_data_add_6_buff_reg[4]  ( .D(n2180), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_6_buff [4]) );
  DF3 \u_decoder/fir_filter/I_data_add_6_buff_reg[3]  ( .D(n2181), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_6_buff [3]) );
  DF3 \u_decoder/fir_filter/I_data_add_6_buff_reg[2]  ( .D(n2182), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_6_buff [2]) );
  DF3 \u_decoder/fir_filter/I_data_add_6_buff_reg[1]  ( .D(n2183), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_6_buff [1]) );
  DF3 \u_decoder/fir_filter/I_data_add_6_buff_reg[0]  ( .D(n2184), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_6_buff [0]), .QN(n90) );
  DF3 \u_decoder/fir_filter/I_data_add_7_buff_reg[14]  ( .D(n2185), .C(inClock), .Q(\u_decoder/fir_filter/I_data_add_7_buff [14]) );
  DF3 \u_decoder/fir_filter/I_data_add_7_buff_reg[13]  ( .D(n2186), .C(inClock), .Q(\u_decoder/fir_filter/I_data_add_7_buff [13]) );
  DF3 \u_decoder/fir_filter/I_data_add_7_buff_reg[12]  ( .D(n2187), .C(inClock), .Q(\u_decoder/fir_filter/I_data_add_7_buff [12]) );
  DF3 \u_decoder/fir_filter/I_data_add_7_buff_reg[11]  ( .D(n2188), .C(inClock), .Q(\u_decoder/fir_filter/I_data_add_7_buff [11]) );
  DF3 \u_decoder/fir_filter/I_data_add_7_buff_reg[10]  ( .D(n2189), .C(inClock), .Q(\u_decoder/fir_filter/I_data_add_7_buff [10]) );
  DF3 \u_decoder/fir_filter/I_data_add_7_buff_reg[9]  ( .D(n2190), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_7_buff [9]) );
  DF3 \u_decoder/fir_filter/I_data_add_7_buff_reg[8]  ( .D(n2191), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_7_buff [8]) );
  DF3 \u_decoder/fir_filter/I_data_add_7_buff_reg[7]  ( .D(n2192), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_7_buff [7]) );
  DF3 \u_decoder/fir_filter/I_data_add_7_buff_reg[6]  ( .D(n2193), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_7_buff [6]) );
  DF3 \u_decoder/fir_filter/I_data_add_7_buff_reg[5]  ( .D(n2194), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_7_buff [5]) );
  DF3 \u_decoder/fir_filter/I_data_add_7_buff_reg[4]  ( .D(n2195), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_7_buff [4]) );
  DF3 \u_decoder/fir_filter/I_data_add_7_buff_reg[3]  ( .D(n2196), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_7_buff [3]) );
  DF3 \u_decoder/fir_filter/I_data_add_7_buff_reg[2]  ( .D(n2197), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_7_buff [2]) );
  DF3 \u_decoder/fir_filter/I_data_add_7_buff_reg[1]  ( .D(n2198), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_7_buff [1]) );
  DF3 \u_decoder/fir_filter/I_data_add_7_buff_reg[0]  ( .D(n2199), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_7_buff [0]), .QN(n89) );
  DF3 \u_decoder/fir_filter/I_data_mult_8_buff_reg[0]  ( .D(
        \u_decoder/fir_filter/n1303 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_8_buff [0]), .QN(n87) );
  DF3 \u_decoder/fir_filter/I_data_mult_8_buff_reg[1]  ( .D(
        \u_decoder/fir_filter/n1304 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_8_buff [1]) );
  DF3 \u_decoder/fir_filter/I_data_mult_8_buff_reg[2]  ( .D(
        \u_decoder/fir_filter/n1305 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_8_buff [2]) );
  DF3 \u_decoder/fir_filter/I_data_mult_8_buff_reg[3]  ( .D(
        \u_decoder/fir_filter/n1306 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_8_buff [3]) );
  DF3 \u_decoder/fir_filter/I_data_mult_8_buff_reg[4]  ( .D(
        \u_decoder/fir_filter/n1307 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_8_buff [4]) );
  DF3 \u_decoder/fir_filter/I_data_mult_8_buff_reg[5]  ( .D(
        \u_decoder/fir_filter/n1308 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_8_buff [5]) );
  DF3 \u_decoder/fir_filter/I_data_mult_8_buff_reg[6]  ( .D(
        \u_decoder/fir_filter/n1309 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_8_buff [6]) );
  DF3 \u_decoder/fir_filter/I_data_mult_8_buff_reg[7]  ( .D(
        \u_decoder/fir_filter/n1310 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_8_buff [7]) );
  DF3 \u_decoder/fir_filter/I_data_mult_8_buff_reg[8]  ( .D(
        \u_decoder/fir_filter/n1311 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_8_buff [8]) );
  DF3 \u_decoder/fir_filter/I_data_mult_8_buff_reg[9]  ( .D(
        \u_decoder/fir_filter/n1312 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_8_buff [9]) );
  DF3 \u_decoder/fir_filter/I_data_mult_8_buff_reg[10]  ( .D(
        \u_decoder/fir_filter/n1313 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_8_buff [10]) );
  DF3 \u_decoder/fir_filter/I_data_mult_8_buff_reg[11]  ( .D(
        \u_decoder/fir_filter/n1314 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_8_buff [11]) );
  DF3 \u_decoder/fir_filter/I_data_mult_8_buff_reg[12]  ( .D(
        \u_decoder/fir_filter/n1315 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_8_buff [12]) );
  DF3 \u_decoder/fir_filter/I_data_mult_8_buff_reg[13]  ( .D(
        \u_decoder/fir_filter/n1316 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_8_buff [13]) );
  DF3 \u_decoder/fir_filter/I_data_mult_8_buff_reg[14]  ( .D(
        \u_decoder/fir_filter/n1317 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_8_buff [14]) );
  DF3 \u_decoder/fir_filter/I_data_mult_8_delay_reg[0]  ( .D(
        \u_decoder/fir_filter/n1324 ), .C(inClock), .QN(
        \u_decoder/fir_filter/n426 ) );
  DF3 \u_decoder/fir_filter/I_data_mult_8_delay_reg[1]  ( .D(
        \u_decoder/fir_filter/n1325 ), .C(inClock), .QN(
        \u_decoder/fir_filter/n425 ) );
  DF3 \u_decoder/fir_filter/I_data_mult_8_delay_reg[2]  ( .D(
        \u_decoder/fir_filter/n1326 ), .C(inClock), .QN(
        \u_decoder/fir_filter/n424 ) );
  DF3 \u_decoder/fir_filter/I_data_mult_8_delay_reg[3]  ( .D(
        \u_decoder/fir_filter/n1327 ), .C(inClock), .QN(
        \u_decoder/fir_filter/n423 ) );
  DF3 \u_decoder/fir_filter/I_data_mult_8_delay_reg[4]  ( .D(
        \u_decoder/fir_filter/n1328 ), .C(inClock), .QN(
        \u_decoder/fir_filter/n422 ) );
  DF3 \u_decoder/fir_filter/I_data_mult_8_delay_reg[5]  ( .D(
        \u_decoder/fir_filter/n1329 ), .C(inClock), .QN(
        \u_decoder/fir_filter/n421 ) );
  DF3 \u_decoder/fir_filter/I_data_mult_8_delay_reg[6]  ( .D(
        \u_decoder/fir_filter/n1330 ), .C(inClock), .QN(
        \u_decoder/fir_filter/n420 ) );
  DF3 \u_decoder/fir_filter/I_data_mult_8_delay_reg[7]  ( .D(
        \u_decoder/fir_filter/n1331 ), .C(inClock), .QN(
        \u_decoder/fir_filter/n419 ) );
  DF3 \u_decoder/fir_filter/I_data_mult_8_delay_reg[8]  ( .D(
        \u_decoder/fir_filter/n1332 ), .C(inClock), .QN(
        \u_decoder/fir_filter/n418 ) );
  DF3 \u_decoder/fir_filter/I_data_mult_8_delay_reg[9]  ( .D(
        \u_decoder/fir_filter/n1333 ), .C(inClock), .QN(
        \u_decoder/fir_filter/n417 ) );
  DF3 \u_decoder/fir_filter/I_data_mult_8_delay_reg[10]  ( .D(
        \u_decoder/fir_filter/n1334 ), .C(inClock), .QN(
        \u_decoder/fir_filter/n416 ) );
  DF3 \u_decoder/fir_filter/I_data_mult_8_delay_reg[11]  ( .D(
        \u_decoder/fir_filter/n1335 ), .C(inClock), .QN(
        \u_decoder/fir_filter/n415 ) );
  DF3 \u_decoder/fir_filter/I_data_mult_8_delay_reg[12]  ( .D(
        \u_decoder/fir_filter/n1336 ), .C(inClock), .QN(
        \u_decoder/fir_filter/n414 ) );
  DF3 \u_decoder/fir_filter/I_data_mult_8_delay_reg[13]  ( .D(
        \u_decoder/fir_filter/n1337 ), .C(inClock), .QN(
        \u_decoder/fir_filter/n413 ) );
  DF3 \u_decoder/fir_filter/I_data_mult_8_delay_reg[14]  ( .D(
        \u_decoder/fir_filter/n1338 ), .C(inClock), .QN(
        \u_decoder/fir_filter/n412 ) );
  DF3 \u_decoder/fir_filter/I_data_mult_7_buff_reg[0]  ( .D(
        \u_decoder/fir_filter/n1340 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_7_buff [0]), .QN(n9) );
  DF3 \u_decoder/fir_filter/I_data_mult_7_buff_reg[1]  ( .D(
        \u_decoder/fir_filter/n1341 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_7_buff [1]) );
  DF3 \u_decoder/fir_filter/I_data_mult_7_buff_reg[2]  ( .D(
        \u_decoder/fir_filter/n1342 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_7_buff [2]) );
  DF3 \u_decoder/fir_filter/I_data_mult_7_buff_reg[3]  ( .D(
        \u_decoder/fir_filter/n1343 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_7_buff [3]) );
  DF3 \u_decoder/fir_filter/I_data_mult_7_buff_reg[4]  ( .D(
        \u_decoder/fir_filter/n1344 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_7_buff [4]) );
  DF3 \u_decoder/fir_filter/I_data_mult_7_buff_reg[5]  ( .D(
        \u_decoder/fir_filter/n1345 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_7_buff [5]) );
  DF3 \u_decoder/fir_filter/I_data_mult_7_buff_reg[6]  ( .D(
        \u_decoder/fir_filter/n1346 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_7_buff [6]) );
  DF3 \u_decoder/fir_filter/I_data_mult_7_buff_reg[7]  ( .D(
        \u_decoder/fir_filter/n1347 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_7_buff [7]) );
  DF3 \u_decoder/fir_filter/I_data_mult_7_buff_reg[8]  ( .D(
        \u_decoder/fir_filter/n1348 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_7_buff [8]) );
  DF3 \u_decoder/fir_filter/I_data_mult_7_buff_reg[9]  ( .D(
        \u_decoder/fir_filter/n1349 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_7_buff [9]) );
  DF3 \u_decoder/fir_filter/I_data_mult_7_buff_reg[10]  ( .D(
        \u_decoder/fir_filter/n1350 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_7_buff [10]) );
  DF3 \u_decoder/fir_filter/I_data_mult_7_buff_reg[11]  ( .D(
        \u_decoder/fir_filter/n1351 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_7_buff [11]) );
  DF3 \u_decoder/fir_filter/I_data_mult_7_buff_reg[12]  ( .D(
        \u_decoder/fir_filter/n1352 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_7_buff [12]) );
  DF3 \u_decoder/fir_filter/I_data_mult_7_buff_reg[13]  ( .D(
        \u_decoder/fir_filter/n1353 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_7_buff [13]) );
  DF3 \u_decoder/fir_filter/I_data_mult_7_buff_reg[14]  ( .D(
        \u_decoder/fir_filter/n1354 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_7_buff [14]) );
  DF3 \u_decoder/fir_filter/I_data_mult_6_buff_reg[0]  ( .D(n2200), .C(inClock), .Q(\u_decoder/fir_filter/I_data_mult_6_buff [0]), .QN(n11) );
  DF3 \u_decoder/fir_filter/I_data_mult_6_buff_reg[1]  ( .D(
        \u_decoder/fir_filter/n1357 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_6_buff [1]) );
  DF3 \u_decoder/fir_filter/I_data_mult_6_buff_reg[2]  ( .D(
        \u_decoder/fir_filter/n1358 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_6_buff [2]) );
  DF3 \u_decoder/fir_filter/I_data_mult_6_buff_reg[3]  ( .D(
        \u_decoder/fir_filter/n1359 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_6_buff [3]) );
  DF3 \u_decoder/fir_filter/I_data_mult_6_buff_reg[4]  ( .D(
        \u_decoder/fir_filter/n1360 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_6_buff [4]) );
  DF3 \u_decoder/fir_filter/I_data_mult_6_buff_reg[5]  ( .D(
        \u_decoder/fir_filter/n1361 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_6_buff [5]) );
  DF3 \u_decoder/fir_filter/I_data_mult_6_buff_reg[6]  ( .D(
        \u_decoder/fir_filter/n1362 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_6_buff [6]) );
  DF3 \u_decoder/fir_filter/I_data_mult_6_buff_reg[7]  ( .D(
        \u_decoder/fir_filter/n1363 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_6_buff [7]) );
  DF3 \u_decoder/fir_filter/I_data_mult_6_buff_reg[8]  ( .D(
        \u_decoder/fir_filter/n1364 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_6_buff [8]) );
  DF3 \u_decoder/fir_filter/I_data_mult_6_buff_reg[9]  ( .D(
        \u_decoder/fir_filter/n1365 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_6_buff [9]) );
  DF3 \u_decoder/fir_filter/I_data_mult_6_buff_reg[10]  ( .D(
        \u_decoder/fir_filter/n1366 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_6_buff [10]) );
  DF3 \u_decoder/fir_filter/I_data_mult_6_buff_reg[11]  ( .D(
        \u_decoder/fir_filter/n1367 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_6_buff [11]) );
  DF3 \u_decoder/fir_filter/I_data_mult_6_buff_reg[12]  ( .D(
        \u_decoder/fir_filter/n1368 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_6_buff [12]) );
  DF3 \u_decoder/fir_filter/I_data_mult_6_buff_reg[13]  ( .D(
        \u_decoder/fir_filter/n1369 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_6_buff [13]) );
  DF3 \u_decoder/fir_filter/I_data_mult_6_buff_reg[14]  ( .D(
        \u_decoder/fir_filter/n1370 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_6_buff [14]) );
  DF3 \u_decoder/fir_filter/I_data_mult_5_buff_reg[0]  ( .D(
        \u_decoder/fir_filter/n1372 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_5_buff [0]), .QN(n12) );
  DF3 \u_decoder/fir_filter/I_data_mult_5_buff_reg[1]  ( .D(
        \u_decoder/fir_filter/n1373 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_5_buff [1]) );
  DF3 \u_decoder/fir_filter/I_data_mult_5_buff_reg[2]  ( .D(
        \u_decoder/fir_filter/n1374 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_5_buff [2]) );
  DF3 \u_decoder/fir_filter/I_data_mult_5_buff_reg[3]  ( .D(
        \u_decoder/fir_filter/n1375 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_5_buff [3]) );
  DF3 \u_decoder/fir_filter/I_data_mult_5_buff_reg[4]  ( .D(
        \u_decoder/fir_filter/n1376 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_5_buff [4]) );
  DF3 \u_decoder/fir_filter/I_data_mult_5_buff_reg[5]  ( .D(
        \u_decoder/fir_filter/n1377 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_5_buff [5]) );
  DF3 \u_decoder/fir_filter/I_data_mult_5_buff_reg[6]  ( .D(
        \u_decoder/fir_filter/n1378 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_5_buff [6]) );
  DF3 \u_decoder/fir_filter/I_data_mult_5_buff_reg[7]  ( .D(
        \u_decoder/fir_filter/n1379 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_5_buff [7]) );
  DF3 \u_decoder/fir_filter/I_data_mult_5_buff_reg[8]  ( .D(
        \u_decoder/fir_filter/n1380 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_5_buff [8]) );
  DF3 \u_decoder/fir_filter/I_data_mult_5_buff_reg[9]  ( .D(
        \u_decoder/fir_filter/n1381 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_5_buff [9]) );
  DF3 \u_decoder/fir_filter/I_data_mult_5_buff_reg[10]  ( .D(
        \u_decoder/fir_filter/n1382 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_5_buff [10]) );
  DF3 \u_decoder/fir_filter/I_data_mult_5_buff_reg[11]  ( .D(
        \u_decoder/fir_filter/n1383 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_5_buff [11]) );
  DF3 \u_decoder/fir_filter/I_data_mult_5_buff_reg[12]  ( .D(
        \u_decoder/fir_filter/n1384 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_5_buff [12]) );
  DF3 \u_decoder/fir_filter/I_data_mult_5_buff_reg[13]  ( .D(
        \u_decoder/fir_filter/n1385 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_5_buff [13]) );
  DF3 \u_decoder/fir_filter/I_data_mult_5_buff_reg[14]  ( .D(
        \u_decoder/fir_filter/n1386 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_5_buff [14]) );
  DF3 \u_decoder/fir_filter/I_data_mult_4_buff_reg[0]  ( .D(n1818), .C(inClock), .Q(\u_decoder/fir_filter/I_data_mult_4_buff [0]), .QN(n21) );
  DF3 \u_decoder/fir_filter/I_data_mult_4_buff_reg[1]  ( .D(n1861), .C(inClock), .Q(\u_decoder/fir_filter/I_data_mult_4_buff [1]) );
  DF3 \u_decoder/fir_filter/I_data_mult_4_buff_reg[2]  ( .D(n1863), .C(inClock), .Q(\u_decoder/fir_filter/I_data_mult_4_buff [2]) );
  DF3 \u_decoder/fir_filter/I_data_mult_4_buff_reg[3]  ( .D(n1836), .C(inClock), .Q(\u_decoder/fir_filter/I_data_mult_4_buff [3]) );
  DF3 \u_decoder/fir_filter/I_data_mult_4_buff_reg[4]  ( .D(n1835), .C(inClock), .Q(\u_decoder/fir_filter/I_data_mult_4_buff [4]) );
  DF3 \u_decoder/fir_filter/I_data_mult_4_buff_reg[5]  ( .D(n1834), .C(inClock), .Q(\u_decoder/fir_filter/I_data_mult_4_buff [5]) );
  DF3 \u_decoder/fir_filter/I_data_mult_4_buff_reg[6]  ( .D(n1833), .C(inClock), .Q(\u_decoder/fir_filter/I_data_mult_4_buff [6]) );
  DF3 \u_decoder/fir_filter/I_data_mult_4_buff_reg[7]  ( .D(n1832), .C(inClock), .Q(\u_decoder/fir_filter/I_data_mult_4_buff [7]) );
  DF3 \u_decoder/fir_filter/I_data_mult_4_buff_reg[8]  ( .D(n1831), .C(inClock), .Q(\u_decoder/fir_filter/I_data_mult_4_buff [8]) );
  DF3 \u_decoder/fir_filter/I_data_mult_4_buff_reg[9]  ( .D(n1830), .C(inClock), .Q(\u_decoder/fir_filter/I_data_mult_4_buff [9]) );
  DF3 \u_decoder/fir_filter/I_data_mult_4_buff_reg[10]  ( .D(n1828), .C(
        inClock), .Q(\u_decoder/fir_filter/I_data_mult_4_buff [10]) );
  DF3 \u_decoder/fir_filter/I_data_mult_4_buff_reg[11]  ( .D(n1824), .C(
        inClock), .Q(\u_decoder/fir_filter/I_data_mult_4_buff [11]) );
  DF3 \u_decoder/fir_filter/I_data_mult_4_buff_reg[12]  ( .D(n1819), .C(
        inClock), .Q(\u_decoder/fir_filter/I_data_mult_4_buff [12]) );
  DF3 \u_decoder/fir_filter/I_data_mult_4_buff_reg[13]  ( .D(n1821), .C(
        inClock), .Q(\u_decoder/fir_filter/I_data_mult_4_buff [13]) );
  DF3 \u_decoder/fir_filter/I_data_mult_4_buff_reg[14]  ( .D(n1822), .C(
        inClock), .Q(\u_decoder/fir_filter/I_data_mult_4_buff [14]) );
  DF3 \u_decoder/fir_filter/I_data_mult_3_buff_reg[0]  ( .D(
        \u_decoder/fir_filter/n1388 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_3_buff [0]), .QN(n13) );
  DF3 \u_decoder/fir_filter/I_data_mult_3_buff_reg[1]  ( .D(
        \u_decoder/fir_filter/n1389 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_3_buff [1]) );
  DF3 \u_decoder/fir_filter/I_data_mult_3_buff_reg[2]  ( .D(
        \u_decoder/fir_filter/n1390 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_3_buff [2]) );
  DF3 \u_decoder/fir_filter/I_data_mult_3_buff_reg[3]  ( .D(
        \u_decoder/fir_filter/n1391 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_3_buff [3]) );
  DF3 \u_decoder/fir_filter/I_data_mult_3_buff_reg[4]  ( .D(
        \u_decoder/fir_filter/n1392 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_3_buff [4]) );
  DF3 \u_decoder/fir_filter/I_data_mult_3_buff_reg[5]  ( .D(
        \u_decoder/fir_filter/n1393 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_3_buff [5]) );
  DF3 \u_decoder/fir_filter/I_data_mult_3_buff_reg[6]  ( .D(
        \u_decoder/fir_filter/n1394 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_3_buff [6]) );
  DF3 \u_decoder/fir_filter/I_data_mult_3_buff_reg[7]  ( .D(
        \u_decoder/fir_filter/n1395 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_3_buff [7]) );
  DF3 \u_decoder/fir_filter/I_data_mult_3_buff_reg[8]  ( .D(
        \u_decoder/fir_filter/n1396 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_3_buff [8]) );
  DF3 \u_decoder/fir_filter/I_data_mult_3_buff_reg[9]  ( .D(
        \u_decoder/fir_filter/n1397 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_3_buff [9]) );
  DF3 \u_decoder/fir_filter/I_data_mult_3_buff_reg[10]  ( .D(
        \u_decoder/fir_filter/n1398 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_3_buff [10]) );
  DF3 \u_decoder/fir_filter/I_data_mult_3_buff_reg[11]  ( .D(
        \u_decoder/fir_filter/n1399 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_3_buff [11]) );
  DF3 \u_decoder/fir_filter/I_data_mult_3_buff_reg[12]  ( .D(
        \u_decoder/fir_filter/n1400 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_3_buff [12]) );
  DF3 \u_decoder/fir_filter/I_data_mult_3_buff_reg[13]  ( .D(
        \u_decoder/fir_filter/n1401 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_3_buff [13]) );
  DF3 \u_decoder/fir_filter/I_data_mult_3_buff_reg[14]  ( .D(
        \u_decoder/fir_filter/n1402 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_3_buff [14]) );
  DF3 \u_decoder/fir_filter/I_data_mult_2_buff_reg[0]  ( .D(n2201), .C(inClock), .Q(\u_decoder/fir_filter/I_data_mult_2_buff [0]), .QN(n14) );
  DF3 \u_decoder/fir_filter/I_data_mult_2_buff_reg[1]  ( .D(
        \u_decoder/fir_filter/n1405 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_2_buff [1]) );
  DF3 \u_decoder/fir_filter/I_data_mult_2_buff_reg[2]  ( .D(
        \u_decoder/fir_filter/n1406 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_2_buff [2]) );
  DF3 \u_decoder/fir_filter/I_data_mult_2_buff_reg[3]  ( .D(
        \u_decoder/fir_filter/n1407 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_2_buff [3]) );
  DF3 \u_decoder/fir_filter/I_data_mult_2_buff_reg[4]  ( .D(
        \u_decoder/fir_filter/n1408 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_2_buff [4]) );
  DF3 \u_decoder/fir_filter/I_data_mult_2_buff_reg[5]  ( .D(
        \u_decoder/fir_filter/n1409 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_2_buff [5]) );
  DF3 \u_decoder/fir_filter/I_data_mult_2_buff_reg[6]  ( .D(
        \u_decoder/fir_filter/n1410 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_2_buff [6]) );
  DF3 \u_decoder/fir_filter/I_data_mult_2_buff_reg[7]  ( .D(
        \u_decoder/fir_filter/n1411 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_2_buff [7]) );
  DF3 \u_decoder/fir_filter/I_data_mult_2_buff_reg[8]  ( .D(
        \u_decoder/fir_filter/n1412 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_2_buff [8]) );
  DF3 \u_decoder/fir_filter/I_data_mult_2_buff_reg[9]  ( .D(
        \u_decoder/fir_filter/n1413 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_2_buff [9]) );
  DF3 \u_decoder/fir_filter/I_data_mult_2_buff_reg[10]  ( .D(
        \u_decoder/fir_filter/n1414 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_2_buff [10]) );
  DF3 \u_decoder/fir_filter/I_data_mult_2_buff_reg[11]  ( .D(
        \u_decoder/fir_filter/n1415 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_2_buff [11]) );
  DF3 \u_decoder/fir_filter/I_data_mult_2_buff_reg[12]  ( .D(
        \u_decoder/fir_filter/n1416 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_2_buff [12]) );
  DF3 \u_decoder/fir_filter/I_data_mult_2_buff_reg[13]  ( .D(
        \u_decoder/fir_filter/n1417 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_2_buff [13]) );
  DF3 \u_decoder/fir_filter/I_data_mult_2_buff_reg[14]  ( .D(
        \u_decoder/fir_filter/n1418 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_2_buff [14]) );
  DF3 \u_decoder/fir_filter/I_data_mult_1_buff_reg[0]  ( .D(
        \u_decoder/fir_filter/n1420 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_1_buff [0]), .QN(n15) );
  DF3 \u_decoder/fir_filter/I_data_mult_1_buff_reg[1]  ( .D(
        \u_decoder/fir_filter/n1421 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_1_buff [1]) );
  DF3 \u_decoder/fir_filter/I_data_mult_1_buff_reg[2]  ( .D(
        \u_decoder/fir_filter/n1422 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_1_buff [2]) );
  DF3 \u_decoder/fir_filter/I_data_mult_1_buff_reg[3]  ( .D(
        \u_decoder/fir_filter/n1423 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_1_buff [3]) );
  DF3 \u_decoder/fir_filter/I_data_mult_1_buff_reg[4]  ( .D(
        \u_decoder/fir_filter/n1424 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_1_buff [4]) );
  DF3 \u_decoder/fir_filter/I_data_mult_1_buff_reg[5]  ( .D(
        \u_decoder/fir_filter/n1425 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_1_buff [5]) );
  DF3 \u_decoder/fir_filter/I_data_mult_1_buff_reg[6]  ( .D(
        \u_decoder/fir_filter/n1426 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_1_buff [6]) );
  DF3 \u_decoder/fir_filter/I_data_mult_1_buff_reg[7]  ( .D(
        \u_decoder/fir_filter/n1427 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_1_buff [7]) );
  DF3 \u_decoder/fir_filter/I_data_mult_1_buff_reg[8]  ( .D(
        \u_decoder/fir_filter/n1428 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_1_buff [8]) );
  DF3 \u_decoder/fir_filter/I_data_mult_1_buff_reg[9]  ( .D(
        \u_decoder/fir_filter/n1429 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_1_buff [9]) );
  DF3 \u_decoder/fir_filter/I_data_mult_1_buff_reg[10]  ( .D(
        \u_decoder/fir_filter/n1430 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_1_buff [10]) );
  DF3 \u_decoder/fir_filter/I_data_mult_1_buff_reg[11]  ( .D(
        \u_decoder/fir_filter/n1431 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_1_buff [11]) );
  DF3 \u_decoder/fir_filter/I_data_mult_1_buff_reg[12]  ( .D(
        \u_decoder/fir_filter/n1432 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_1_buff [12]) );
  DF3 \u_decoder/fir_filter/I_data_mult_1_buff_reg[13]  ( .D(
        \u_decoder/fir_filter/n1433 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_1_buff [13]) );
  DF3 \u_decoder/fir_filter/I_data_mult_1_buff_reg[14]  ( .D(
        \u_decoder/fir_filter/n1434 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_1_buff [14]) );
  DF3 \u_decoder/fir_filter/I_data_mult_0_buff_reg[0]  ( .D(
        \u_decoder/fir_filter/n1436 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_0_buff [0]) );
  DF3 \u_decoder/fir_filter/I_data_mult_0_buff_reg[1]  ( .D(
        \u_decoder/fir_filter/n1437 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_0_buff [1]), .QN(n74) );
  DF3 \u_decoder/fir_filter/I_data_mult_0_buff_reg[2]  ( .D(
        \u_decoder/fir_filter/n1438 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_0_buff [2]), .QN(n72) );
  DF3 \u_decoder/fir_filter/I_data_mult_0_buff_reg[3]  ( .D(
        \u_decoder/fir_filter/n1439 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_0_buff [3]), .QN(n113) );
  DF3 \u_decoder/fir_filter/I_data_mult_0_buff_reg[4]  ( .D(
        \u_decoder/fir_filter/n1440 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_0_buff [4]), .QN(n130) );
  DF3 \u_decoder/fir_filter/I_data_mult_0_buff_reg[5]  ( .D(
        \u_decoder/fir_filter/n1441 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_0_buff [5]), .QN(n131) );
  DF3 \u_decoder/fir_filter/I_data_mult_0_buff_reg[6]  ( .D(
        \u_decoder/fir_filter/n1442 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_0_buff [6]), .QN(n143) );
  DF3 \u_decoder/fir_filter/I_data_mult_0_buff_reg[7]  ( .D(
        \u_decoder/fir_filter/n1443 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_0_buff [7]) );
  DF3 \u_decoder/fir_filter/I_data_mult_0_buff_reg[8]  ( .D(
        \u_decoder/fir_filter/n1444 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_0_buff [8]), .QN(n199) );
  DF3 \u_decoder/fir_filter/I_data_mult_0_buff_reg[9]  ( .D(
        \u_decoder/fir_filter/n1445 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_0_buff [9]) );
  DF3 \u_decoder/fir_filter/I_data_mult_0_buff_reg[10]  ( .D(
        \u_decoder/fir_filter/n1446 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_0_buff [10]), .QN(n259) );
  DF3 \u_decoder/fir_filter/I_data_mult_0_buff_reg[11]  ( .D(
        \u_decoder/fir_filter/n1447 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_0_buff [11]) );
  DF3 \u_decoder/fir_filter/I_data_mult_0_buff_reg[12]  ( .D(
        \u_decoder/fir_filter/n1448 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_0_buff [12]) );
  DF3 \u_decoder/fir_filter/I_data_mult_0_buff_reg[13]  ( .D(
        \u_decoder/fir_filter/n1449 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_0_buff [13]) );
  DF3 \u_decoder/fir_filter/I_data_mult_0_buff_reg[14]  ( .D(
        \u_decoder/fir_filter/n1450 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_0_buff [14]) );
  DF3 \u_decoder/fir_filter/o_postfilter_ready_reg  ( .D(
        \u_decoder/fir_filter/n1451 ), .C(inClock), .Q(\sig_MUX_inMUX8[0] ) );
  DF3 \u_decoder/fir_filter/state_reg[0]  ( .D(\u_decoder/fir_filter/N11 ), 
        .C(inClock), .Q(\u_decoder/fir_filter/state [0]), .QN(
        \u_decoder/fir_filter/n410 ) );
  DF3 \u_decoder/fir_filter/state_reg[1]  ( .D(\u_decoder/fir_filter/N12 ), 
        .C(inClock), .Q(\u_decoder/fir_filter/state [1]) );
  DF3 \u_cordic/mycordic/o_angle_reg[15]  ( .D(n1542), .C(inClock), .Q(
        \u_cordic/cordic_to_rotation [15]) );
  DF3 \u_cordic/mycordic/o_angle_reg[14]  ( .D(n1543), .C(inClock), .Q(
        \u_cordic/cordic_to_rotation [14]) );
  DF3 \u_cordic/mycordic/o_angle_reg[13]  ( .D(n1544), .C(inClock), .Q(
        \u_cordic/cordic_to_rotation [13]) );
  DF3 \u_cordic/mycordic/o_angle_reg[12]  ( .D(n1545), .C(inClock), .Q(
        \u_cordic/cordic_to_rotation [12]) );
  DF3 \u_cordic/mycordic/o_angle_reg[11]  ( .D(n1546), .C(inClock), .Q(
        \u_cordic/cordic_to_rotation [11]) );
  DF3 \u_cordic/mycordic/o_angle_reg[10]  ( .D(n1547), .C(inClock), .Q(
        \u_cordic/cordic_to_rotation [10]) );
  DF3 \u_cordic/mycordic/o_angle_reg[9]  ( .D(n1548), .C(inClock), .Q(
        \u_cordic/cordic_to_rotation [9]) );
  DF3 \u_cordic/mycordic/o_angle_reg[8]  ( .D(n1549), .C(inClock), .Q(
        \u_cordic/cordic_to_rotation [8]) );
  DF3 \u_cordic/mycordic/o_angle_reg[7]  ( .D(n1550), .C(inClock), .Q(
        \u_cordic/cordic_to_rotation [7]) );
  DF3 \u_cordic/mycordic/o_angle_reg[6]  ( .D(n1551), .C(inClock), .Q(
        \u_cordic/cordic_to_rotation [6]) );
  DF3 \u_cordic/mycordic/o_angle_reg[5]  ( .D(n1552), .C(inClock), .Q(
        \u_cordic/cordic_to_rotation [5]) );
  DF3 \u_cordic/mycordic/o_angle_reg[4]  ( .D(n1553), .C(inClock), .Q(
        \u_cordic/cordic_to_rotation [4]) );
  DF3 \u_cordic/mycordic/o_angle_reg[3]  ( .D(n1554), .C(inClock), .Q(
        \u_cordic/cordic_to_rotation [3]) );
  DF3 \u_cordic/mycordic/o_angle_reg[2]  ( .D(n1556), .C(inClock), .Q(
        \u_cordic/cordic_to_rotation [2]) );
  DF3 \u_cordic/mycordic/o_angle_reg[1]  ( .D(n1567), .C(inClock), .Q(
        \u_cordic/cordic_to_rotation [1]) );
  DF3 \u_cordic/mycordic/o_angle_reg[0]  ( .D(n1576), .C(inClock), .Q(
        \u_cordic/cordic_to_rotation [0]) );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[6][15]  ( .D(n1194), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[6][15] ) );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[6][14]  ( .D(n1193), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[6][14] ), .QN(n279) );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[6][13]  ( .D(n1192), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[6][13] ), .QN(n260) );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[6][12]  ( .D(n1191), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[6][12] ), .QN(n235) );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[6][11]  ( .D(n1190), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[6][11] ), .QN(n234) );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[6][10]  ( .D(n1189), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[6][10] ), .QN(n200) );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[6][9]  ( .D(n1188), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[6][9] ), .QN(n169)
         );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[6][8]  ( .D(n1187), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[6][8] ), .QN(n144)
         );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[6][7]  ( .D(n1186), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[6][7] ), .QN(n377)
         );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[6][6]  ( .D(n1185), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[6][6] ), .QN(n132)
         );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[6][5]  ( .D(n1184), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[6][5] ), .QN(n382)
         );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[6][4]  ( .D(n1183), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[6][4] ), .QN(n385)
         );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[6][3]  ( .D(n1182), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[6][3] ), .QN(n303)
         );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[6][2]  ( .D(n1181), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[6][2] ), .QN(n75)
         );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[6][1]  ( .D(n1180), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[6][1] ), .QN(n311)
         );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[6][0]  ( .D(n1179), .C(
        inClock), .Q(\u_cordic/mycordic/N615 ), .QN(n310) );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[5][15]  ( .D(n1254), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[5][15] ) );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[5][14]  ( .D(n1253), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[5][14] ), .QN(n307) );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[5][13]  ( .D(n1252), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[5][13] ), .QN(n288) );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[5][12]  ( .D(n1251), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[5][12] ), .QN(n265) );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[5][11]  ( .D(n1250), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[5][11] ), .QN(n240) );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[5][10]  ( .D(n1249), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[5][10] ), .QN(n207) );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[5][9]  ( .D(n1248), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[5][9] ), .QN(n208)
         );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[5][8]  ( .D(n1247), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[5][8] ), .QN(n177)
         );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[5][7]  ( .D(n1246), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[5][7] ), .QN(n149)
         );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[5][6]  ( .D(n1245), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[5][6] ), .QN(n138)
         );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[5][5]  ( .D(n1244), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[5][5] ), .QN(n122)
         );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[5][4]  ( .D(n1243), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[5][4] ), .QN(n121)
         );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[5][3]  ( .D(n1242), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[5][3] ), .QN(n86)
         );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[5][2]  ( .D(n1241), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[5][2] ), .QN(n62)
         );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[5][1]  ( .D(n1240), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[5][1] ), .QN(n301)
         );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[5][0]  ( .D(n1239), .C(
        inClock), .Q(\u_cordic/mycordic/N550 ) );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[4][15]  ( .D(n1278), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[4][15] ) );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[4][14]  ( .D(n1277), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[4][14] ), .QN(n306) );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[4][13]  ( .D(n1276), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[4][13] ), .QN(n284) );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[4][12]  ( .D(n1275), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[4][12] ), .QN(n264) );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[4][11]  ( .D(n1274), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[4][11] ), .QN(n239) );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[4][10]  ( .D(n1273), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[4][10] ), .QN(n206) );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[4][9]  ( .D(n1272), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[4][9] ), .QN(n205)
         );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[4][8]  ( .D(n1271), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[4][8] ), .QN(n176)
         );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[4][7]  ( .D(n1270), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[4][7] ), .QN(n148)
         );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[4][6]  ( .D(n1269), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[4][6] ), .QN(n137)
         );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[4][5]  ( .D(n1268), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[4][5] ), .QN(n120)
         );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[4][4]  ( .D(n1267), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[4][4] ), .QN(n119)
         );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[4][3]  ( .D(n1266), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[4][3] ), .QN(n85)
         );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[4][2]  ( .D(n1265), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[4][2] ), .QN(n63)
         );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[4][1]  ( .D(n1264), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[4][1] ), .QN(n78)
         );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[4][0]  ( .D(n1263), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[4][0] ), .QN(n300)
         );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[3][15]  ( .D(n1303), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[3][15] ) );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[3][14]  ( .D(n1302), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[3][14] ), .QN(n287) );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[3][13]  ( .D(n1301), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[3][13] ), .QN(n283) );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[3][12]  ( .D(n1300), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[3][12] ), .QN(n263) );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[3][11]  ( .D(n1299), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[3][11] ), .QN(n238) );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[3][10]  ( .D(n1298), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[3][10] ), .QN(n204) );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[3][9]  ( .D(n1297), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[3][9] ), .QN(n175)
         );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[3][8]  ( .D(n1296), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[3][8] ), .QN(n174)
         );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[3][7]  ( .D(n1295), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[3][7] ), .QN(n147)
         );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[3][6]  ( .D(n1294), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[3][6] ), .QN(n136)
         );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[3][5]  ( .D(n1293), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[3][5] ), .QN(n118)
         );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[3][4]  ( .D(n1292), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[3][4] ), .QN(n84)
         );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[3][3]  ( .D(n1291), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[3][3] ), .QN(n83)
         );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[3][2]  ( .D(n1290), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[3][2] ), .QN(n79)
         );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[3][1]  ( .D(n1289), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[3][1] ), .QN(n81)
         );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[3][0]  ( .D(n1288), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[3][0] ), .QN(n299)
         );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[2][15]  ( .D(n1210), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[2][15] ) );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[2][14]  ( .D(n1209), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[2][14] ), .QN(n286) );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[2][13]  ( .D(n1208), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[2][13] ), .QN(n282) );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[2][12]  ( .D(n1207), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[2][12] ), .QN(n262) );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[2][11]  ( .D(n1206), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[2][11] ), .QN(n237) );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[2][10]  ( .D(n1205), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[2][10] ), .QN(n203) );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[2][9]  ( .D(n1204), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[2][9] ), .QN(n173)
         );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[2][8]  ( .D(n1203), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[2][8] ), .QN(n172)
         );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[2][7]  ( .D(n1202), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[2][7] ), .QN(n146)
         );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[2][6]  ( .D(n1201), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[2][6] ), .QN(n135)
         );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[2][5]  ( .D(n1200), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[2][5] ), .QN(n117)
         );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[2][4]  ( .D(n1199), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[2][4] ), .QN(n82)
         );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[2][3]  ( .D(n1198), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[2][3] ), .QN(n114)
         );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[2][2]  ( .D(n1197), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[2][2] ), .QN(n80)
         );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[2][1]  ( .D(n1196), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[2][1] ), .QN(n297)
         );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[2][0]  ( .D(n1195), .C(
        inClock), .Q(\u_cordic/mycordic/N428 ) );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[1][15]  ( .D(n1579), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[1][15] ) );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[1][14]  ( .D(n1579), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[1][14] ), .QN(n285) );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[1][13]  ( .D(n1579), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[1][13] ), .QN(n281) );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[1][12]  ( .D(n1579), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[1][12] ), .QN(n261) );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[1][11]  ( .D(n1579), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[1][11] ), .QN(n236) );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[1][10]  ( .D(n1579), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[1][10] ), .QN(n202) );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[1][9]  ( .D(n1579), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[1][9] ), .QN(n171)
         );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[1][8]  ( .D(n1579), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[1][8] ), .QN(n170)
         );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[1][7]  ( .D(n1579), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[1][7] ), .QN(n145)
         );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[1][6]  ( .D(n1579), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[1][6] ), .QN(n134)
         );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[1][5]  ( .D(n787), .C(inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[1][5] ), .QN(n116) );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[1][4]  ( .D(n1579), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[1][4] ), .QN(n133)
         );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[1][3]  ( .D(n787), .C(inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[1][3] ), .QN(n115) );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[1][2]  ( .D(n787), .C(inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[1][2] ), .QN(n4) );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[1][1]  ( .D(n1579), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[1][1] ), .QN(n77)
         );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[1][0]  ( .D(n1227), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[1][0] ), .QN(n298)
         );
  DF3 \u_cordic/mycordic/present_C_table_reg[7][0]  ( .D(n1558), .C(inClock), 
        .Q(\u_cordic/mycordic/present_C_table[7][0] ) );
  DF3 \u_cordic/mycordic/present_C_table_reg[6][0]  ( .D(n1561), .C(inClock), 
        .Q(\u_cordic/mycordic/present_C_table[6][0] ) );
  DF3 \u_cordic/mycordic/present_C_table_reg[5][0]  ( .D(n1564), .C(inClock), 
        .Q(\u_cordic/mycordic/present_C_table[5][0] ) );
  DF3 \u_cordic/mycordic/present_C_table_reg[4][0]  ( .D(n1568), .C(inClock), 
        .Q(\u_cordic/mycordic/present_C_table[4][0] ) );
  DF3 \u_cordic/mycordic/present_C_table_reg[3][0]  ( .D(n1571), .C(inClock), 
        .Q(\u_cordic/mycordic/present_C_table[3][0] ) );
  DF3 \u_cordic/mycordic/present_C_table_reg[2][0]  ( .D(n1574), .C(inClock), 
        .Q(\u_cordic/mycordic/present_C_table[2][0] ) );
  DF3 \u_cordic/mycordic/present_C_table_reg[1][0]  ( .D(n1168), .C(inClock), 
        .Q(\u_cordic/mycordic/present_C_table[1][0] ) );
  DF3 \u_cordic/mycordic/present_C_table_reg[7][1]  ( .D(n1557), .C(inClock), 
        .Q(\u_cordic/mycordic/present_C_table[7][1] ), .QN(
        \u_cordic/mycordic/n110 ) );
  DF3 \u_cordic/mycordic/present_C_table_reg[6][1]  ( .D(n1560), .C(inClock), 
        .Q(\u_cordic/mycordic/present_C_table[6][1] ) );
  DF3 \u_cordic/mycordic/present_C_table_reg[5][1]  ( .D(n1563), .C(inClock), 
        .Q(\u_cordic/mycordic/present_C_table[5][1] ) );
  DF3 \u_cordic/mycordic/present_C_table_reg[4][1]  ( .D(n1566), .C(inClock), 
        .Q(\u_cordic/mycordic/present_C_table[4][1] ) );
  DF3 \u_cordic/mycordic/present_C_table_reg[3][1]  ( .D(n1570), .C(inClock), 
        .Q(\u_cordic/mycordic/present_C_table[3][1] ) );
  DF3 \u_cordic/mycordic/present_C_table_reg[2][1]  ( .D(n1573), .C(inClock), 
        .Q(\u_cordic/mycordic/present_C_table[2][1] ) );
  DF3 \u_cordic/mycordic/present_C_table_reg[1][1]  ( .D(
        \u_cordic/mycordic/N211 ), .C(inClock), .Q(
        \u_cordic/mycordic/present_C_table[1][1] ) );
  DF3 \u_cordic/mycordic/present_C_table_reg[7][2]  ( .D(n1555), .C(inClock), 
        .QN(\u_cordic/mycordic/n108 ) );
  DF3 \u_cordic/mycordic/present_C_table_reg[6][2]  ( .D(n1559), .C(inClock), 
        .Q(\u_cordic/mycordic/present_C_table[6][2] ) );
  DF3 \u_cordic/mycordic/present_C_table_reg[5][2]  ( .D(n1562), .C(inClock), 
        .Q(\u_cordic/mycordic/present_C_table[5][2] ) );
  DF3 \u_cordic/mycordic/present_C_table_reg[4][2]  ( .D(n1565), .C(inClock), 
        .Q(\u_cordic/mycordic/present_C_table[4][2] ) );
  DF3 \u_cordic/mycordic/present_C_table_reg[3][2]  ( .D(n1569), .C(inClock), 
        .Q(\u_cordic/mycordic/present_C_table[3][2] ) );
  DF3 \u_cordic/mycordic/present_C_table_reg[2][2]  ( .D(n1572), .C(inClock), 
        .Q(\u_cordic/mycordic/present_C_table[2][2] ) );
  DF3 \u_cordic/mycordic/present_C_table_reg[1][2]  ( .D(
        \u_cordic/mycordic/N212 ), .C(inClock), .Q(
        \u_cordic/mycordic/present_C_table[1][2] ) );
  DF3 \u_cordic/mycordic/present_Q_table_reg[6][7]  ( .D(n1238), .C(inClock), 
        .Q(\u_cordic/mycordic/present_Q_table[6][7] ) );
  DF3 \u_cordic/mycordic/present_Q_table_reg[5][7]  ( .D(n1262), .C(inClock), 
        .Q(\u_cordic/mycordic/present_Q_table[5][7] ) );
  DF3 \u_cordic/mycordic/present_Q_table_reg[5][6]  ( .D(n1261), .C(inClock), 
        .Q(\u_cordic/mycordic/present_Q_table[5][6] ), .QN(n269) );
  DF3 \u_cordic/mycordic/present_Q_table_reg[5][5]  ( .D(n1260), .C(inClock), 
        .Q(\u_cordic/mycordic/present_Q_table[5][5] ) );
  DF3 \u_cordic/mycordic/present_Q_table_reg[5][4]  ( .D(n1259), .C(inClock), 
        .Q(\u_cordic/mycordic/present_Q_table[5][4] ), .QN(n217) );
  DF3 \u_cordic/mycordic/present_Q_table_reg[5][3]  ( .D(n1258), .C(inClock), 
        .Q(\u_cordic/mycordic/present_Q_table[5][3] ) );
  DF3 \u_cordic/mycordic/present_Q_table_reg[5][2]  ( .D(n1257), .C(inClock), 
        .Q(\u_cordic/mycordic/present_Q_table[5][2] ), .QN(n156) );
  DF3 \u_cordic/mycordic/present_Q_table_reg[5][1]  ( .D(n1256), .C(inClock), 
        .Q(\u_cordic/mycordic/present_Q_table[5][1] ), .QN(n168) );
  DF3 \u_cordic/mycordic/present_Q_table_reg[5][0]  ( .D(n1255), .C(inClock), 
        .Q(\u_cordic/mycordic/present_Q_table[5][0] ), .QN(n150) );
  DF3 \u_cordic/mycordic/present_I_table_reg[5][7]  ( .D(n1282), .C(inClock), 
        .Q(\u_cordic/mycordic/present_I_table[5][7] ), .QN(n182) );
  DF3 \u_cordic/mycordic/present_I_table_reg[5][6]  ( .D(n1281), .C(inClock), 
        .Q(\u_cordic/mycordic/present_I_table[5][6] ) );
  DF3 \u_cordic/mycordic/present_I_table_reg[5][5]  ( .D(n1280), .C(inClock), 
        .Q(\u_cordic/mycordic/present_I_table[5][5] ), .QN(n32) );
  DF3 \u_cordic/mycordic/present_I_table_reg[5][4]  ( .D(n1279), .C(inClock), 
        .Q(\u_cordic/mycordic/present_I_table[5][4] ) );
  DF3 \u_cordic/mycordic/present_Q_table_reg[4][3]  ( .D(n1283), .C(inClock), 
        .Q(\u_cordic/mycordic/present_Q_table[4][3] ), .QN(n167) );
  DF3 \u_cordic/mycordic/present_Q_table_reg[4][4]  ( .D(n1284), .C(inClock), 
        .Q(\u_cordic/mycordic/present_Q_table[4][4] ) );
  DF3 \u_cordic/mycordic/present_Q_table_reg[4][5]  ( .D(n1285), .C(inClock), 
        .Q(\u_cordic/mycordic/present_Q_table[4][5] ), .QN(n231) );
  DF3 \u_cordic/mycordic/present_Q_table_reg[4][6]  ( .D(n1286), .C(inClock), 
        .Q(\u_cordic/mycordic/present_Q_table[4][6] ) );
  DF3 \u_cordic/mycordic/present_Q_table_reg[4][7]  ( .D(n1287), .C(inClock), 
        .Q(\u_cordic/mycordic/present_Q_table[4][7] ), .QN(n180) );
  DF3 \u_cordic/mycordic/present_I_table_reg[4][0]  ( .D(n1304), .C(inClock), 
        .Q(\u_cordic/mycordic/present_I_table[4][0] ) );
  DF3 \u_cordic/mycordic/present_I_table_reg[4][1]  ( .D(n1305), .C(inClock), 
        .Q(\u_cordic/mycordic/present_I_table[4][1] ), .QN(n201) );
  DF3 \u_cordic/mycordic/present_I_table_reg[4][2]  ( .D(n1306), .C(inClock), 
        .Q(\u_cordic/mycordic/present_I_table[4][2] ), .QN(n232) );
  DF3 \u_cordic/mycordic/present_I_table_reg[4][3]  ( .D(n1307), .C(inClock), 
        .Q(\u_cordic/mycordic/present_I_table[4][3] ), .QN(n155) );
  DF3 \u_cordic/mycordic/present_I_table_reg[4][4]  ( .D(n1308), .C(inClock), 
        .Q(\u_cordic/mycordic/present_I_table[4][4] ), .QN(n184) );
  DF3 \u_cordic/mycordic/present_I_table_reg[4][5]  ( .D(n1309), .C(inClock), 
        .Q(\u_cordic/mycordic/present_I_table[4][5] ), .QN(n183) );
  DF3 \u_cordic/mycordic/present_I_table_reg[4][6]  ( .D(n1310), .C(inClock), 
        .Q(\u_cordic/mycordic/present_I_table[4][6] ), .QN(n218) );
  DF3 \u_cordic/mycordic/present_I_table_reg[4][7]  ( .D(n1311), .C(inClock), 
        .Q(\u_cordic/mycordic/present_I_table[4][7] ), .QN(n214) );
  DF3 \u_cordic/mycordic/present_Q_table_reg[4][0]  ( .D(n1312), .C(inClock), 
        .Q(\u_cordic/mycordic/present_Q_table[4][0] ), .QN(n212) );
  DF3 \u_cordic/mycordic/present_Q_table_reg[4][1]  ( .D(n1313), .C(inClock), 
        .Q(\u_cordic/mycordic/present_Q_table[4][1] ) );
  DF3 \u_cordic/mycordic/present_Q_table_reg[4][2]  ( .D(n1314), .C(inClock), 
        .Q(\u_cordic/mycordic/present_Q_table[4][2] ) );
  DF3 \u_cordic/mycordic/present_Q_table_reg[3][7]  ( .D(n1226), .C(inClock), 
        .Q(\u_cordic/mycordic/present_Q_table[3][7] ), .QN(n242) );
  DF3 \u_cordic/mycordic/present_Q_table_reg[3][6]  ( .D(n1225), .C(inClock), 
        .Q(\u_cordic/mycordic/present_Q_table[3][6] ), .QN(n244) );
  DF3 \u_cordic/mycordic/present_Q_table_reg[3][5]  ( .D(n1224), .C(inClock), 
        .Q(\u_cordic/mycordic/present_Q_table[3][5] ), .QN(n219) );
  DF3 \u_cordic/mycordic/present_Q_table_reg[3][4]  ( .D(n1223), .C(inClock), 
        .Q(\u_cordic/mycordic/present_Q_table[3][4] ), .QN(n185) );
  DF3 \u_cordic/mycordic/present_Q_table_reg[3][3]  ( .D(n1222), .C(inClock), 
        .Q(\u_cordic/mycordic/present_Q_table[3][3] ), .QN(n186) );
  DF3 \u_cordic/mycordic/present_Q_table_reg[3][2]  ( .D(n1221), .C(inClock), 
        .Q(\u_cordic/mycordic/present_Q_table[3][2] ), .QN(n158) );
  DF3 \u_cordic/mycordic/present_Q_table_reg[3][1]  ( .D(n1220), .C(inClock), 
        .Q(\u_cordic/mycordic/present_Q_table[3][1] ) );
  DF3 \u_cordic/mycordic/present_Q_table_reg[3][0]  ( .D(n1219), .C(inClock), 
        .Q(\u_cordic/mycordic/present_Q_table[3][0] ), .QN(n210) );
  DF3 \u_cordic/mycordic/present_I_table_reg[3][7]  ( .D(n1218), .C(inClock), 
        .Q(\u_cordic/mycordic/present_I_table[3][7] ), .QN(n243) );
  DF3 \u_cordic/mycordic/present_I_table_reg[3][6]  ( .D(n1217), .C(inClock), 
        .Q(\u_cordic/mycordic/present_I_table[3][6] ), .QN(n245) );
  DF3 \u_cordic/mycordic/present_I_table_reg[3][5]  ( .D(n1216), .C(inClock), 
        .Q(\u_cordic/mycordic/present_I_table[3][5] ), .QN(n220) );
  DF3 \u_cordic/mycordic/present_I_table_reg[3][4]  ( .D(n1215), .C(inClock), 
        .Q(\u_cordic/mycordic/present_I_table[3][4] ), .QN(n187) );
  DF3 \u_cordic/mycordic/present_I_table_reg[3][3]  ( .D(n1214), .C(inClock), 
        .Q(\u_cordic/mycordic/present_I_table[3][3] ), .QN(n188) );
  DF3 \u_cordic/mycordic/present_I_table_reg[3][2]  ( .D(n1213), .C(inClock), 
        .Q(\u_cordic/mycordic/present_I_table[3][2] ), .QN(n157) );
  DF3 \u_cordic/mycordic/present_I_table_reg[3][1]  ( .D(n1212), .C(inClock), 
        .Q(\u_cordic/mycordic/present_I_table[3][1] ) );
  DF3 \u_cordic/mycordic/present_I_table_reg[3][0]  ( .D(n1211), .C(inClock), 
        .Q(\u_cordic/mycordic/present_I_table[3][0] ), .QN(n209) );
  DF3 \u_cordic/mycordic/present_I_table_reg[2][7]  ( .D(n1232), .C(inClock), 
        .Q(\u_cordic/mycordic/present_I_table[2][7] ), .QN(n270) );
  DF3 \u_cordic/mycordic/present_I_table_reg[2][6]  ( .D(n1231), .C(inClock), 
        .Q(\u_cordic/mycordic/present_I_table[2][6] ), .QN(n248) );
  DF3 \u_cordic/mycordic/present_I_table_reg[2][5]  ( .D(n1230), .C(inClock), 
        .Q(\u_cordic/mycordic/present_I_table[2][5] ), .QN(n249) );
  DF3 \u_cordic/mycordic/present_I_table_reg[2][4]  ( .D(n1229), .C(inClock), 
        .Q(\u_cordic/mycordic/present_I_table[2][4] ), .QN(n222) );
  DF3 \u_cordic/mycordic/present_I_table_reg[2][3]  ( .D(n1228), .C(inClock), 
        .Q(\u_cordic/mycordic/present_I_table[2][3] ), .QN(n191) );
  DF3 \u_cordic/mycordic/present_I_table_reg[2][2]  ( .D(n2), .C(inClock), .Q(
        \u_cordic/mycordic/present_I_table[2][2] ), .QN(n192) );
  DF3 \u_cordic/mycordic/present_I_table_reg[2][1]  ( .D(n2), .C(inClock), .Q(
        \u_cordic/mycordic/present_I_table[2][1] ), .QN(n160) );
  DF3 \u_cordic/mycordic/present_I_table_reg[2][0]  ( .D(n2), .C(inClock), .Q(
        \u_cordic/mycordic/present_I_table[2][0] ), .QN(n178) );
  DF3 \u_cordic/mycordic/present_Q_table_reg[2][7]  ( .D(n1237), .C(inClock), 
        .Q(\u_cordic/mycordic/present_Q_table[2][7] ), .QN(n268) );
  DF3 \u_cordic/mycordic/present_Q_table_reg[2][6]  ( .D(n1236), .C(inClock), 
        .Q(\u_cordic/mycordic/present_Q_table[2][6] ), .QN(n246) );
  DF3 \u_cordic/mycordic/present_Q_table_reg[2][5]  ( .D(n1235), .C(inClock), 
        .Q(\u_cordic/mycordic/present_Q_table[2][5] ), .QN(n247) );
  DF3 \u_cordic/mycordic/present_Q_table_reg[2][4]  ( .D(n1234), .C(inClock), 
        .Q(\u_cordic/mycordic/present_Q_table[2][4] ), .QN(n221) );
  DF3 \u_cordic/mycordic/present_Q_table_reg[2][3]  ( .D(n1233), .C(inClock), 
        .Q(\u_cordic/mycordic/present_Q_table[2][3] ), .QN(n189) );
  DF3 \u_cordic/mycordic/present_Q_table_reg[2][2]  ( .D(n2), .C(inClock), .Q(
        \u_cordic/mycordic/present_Q_table[2][2] ), .QN(n190) );
  DF3 \u_cordic/mycordic/present_Q_table_reg[2][1]  ( .D(n2), .C(inClock), .Q(
        \u_cordic/mycordic/present_Q_table[2][1] ), .QN(n159) );
  DF3 \u_cordic/mycordic/present_Q_table_reg[2][0]  ( .D(n2), .C(inClock), .Q(
        \u_cordic/mycordic/present_Q_table[2][0] ), .QN(n211) );
  DF3 \u_cordic/mycordic/present_Q_table_reg[1][7]  ( .D(n1178), .C(inClock), 
        .Q(\u_cordic/mycordic/present_Q_table[1][7] ), .QN(n277) );
  DF3 \u_cordic/mycordic/present_Q_table_reg[1][6]  ( .D(n1177), .C(inClock), 
        .Q(\u_cordic/mycordic/present_Q_table[1][6] ), .QN(n274) );
  DF3 \u_cordic/mycordic/present_Q_table_reg[1][5]  ( .D(n1176), .C(inClock), 
        .Q(\u_cordic/mycordic/present_Q_table[1][5] ), .QN(n252) );
  DF3 \u_cordic/mycordic/present_Q_table_reg[1][4]  ( .D(n1175), .C(inClock), 
        .Q(\u_cordic/mycordic/present_Q_table[1][4] ), .QN(n253) );
  DF3 \u_cordic/mycordic/present_Q_table_reg[1][3]  ( .D(n1174), .C(inClock), 
        .Q(\u_cordic/mycordic/present_Q_table[1][3] ), .QN(n224) );
  DF3 \u_cordic/mycordic/present_Q_table_reg[0][3]  ( .D(\u_cordic/Q [0]), .C(
        inClock), .Q(\u_cordic/mycordic/present_Q_table[0][3] ), .QN(n254) );
  DF3 \u_cordic/mycordic/present_Q_table_reg[0][4]  ( .D(\u_cordic/Q [1]), .C(
        inClock), .Q(\u_cordic/mycordic/present_Q_table[0][4] ), .QN(n43) );
  DF3 \u_cordic/mycordic/present_Q_table_reg[0][5]  ( .D(\u_cordic/Q [2]), .C(
        inClock), .Q(\u_cordic/mycordic/present_Q_table[0][5] ), .QN(n42) );
  DF3 \u_cordic/mycordic/present_Q_table_reg[0][6]  ( .D(\u_cordic/Q [3]), .C(
        inClock), .Q(\u_cordic/mycordic/present_Q_table[0][6] ), .QN(n41) );
  DF3 \u_cordic/mycordic/present_Q_table_reg[0][7]  ( .D(\u_cordic/Q [3]), .C(
        inClock), .Q(\u_cordic/mycordic/present_Q_table[0][7] ) );
  DF3 \u_cordic/mycordic/present_I_table_reg[1][7]  ( .D(
        \u_cordic/mycordic/N44 ), .C(inClock), .Q(
        \u_cordic/mycordic/present_I_table[1][7] ), .QN(n280) );
  DF3 \u_cordic/mycordic/present_I_table_reg[1][6]  ( .D(n1173), .C(inClock), 
        .Q(\u_cordic/mycordic/present_I_table[1][6] ), .QN(n272) );
  DF3 \u_cordic/mycordic/present_I_table_reg[1][5]  ( .D(n1172), .C(inClock), 
        .Q(\u_cordic/mycordic/present_I_table[1][5] ), .QN(n273) );
  DF3 \u_cordic/mycordic/present_I_table_reg[1][4]  ( .D(n1171), .C(inClock), 
        .Q(\u_cordic/mycordic/present_I_table[1][4] ), .QN(n251) );
  DF3 \u_cordic/mycordic/present_I_table_reg[1][3]  ( .D(n1170), .C(inClock), 
        .Q(\u_cordic/mycordic/present_I_table[1][3] ), .QN(n223) );
  DF3 \u_cordic/mycordic/present_I_table_reg[0][3]  ( .D(\u_cordic/I [0]), .C(
        inClock), .Q(\u_cordic/mycordic/present_I_table[0][3] ), .QN(n257) );
  DF3 \u_cordic/mycordic/present_I_table_reg[0][4]  ( .D(\u_cordic/I [1]), .C(
        inClock), .Q(\u_cordic/mycordic/present_I_table[0][4] ), .QN(n46) );
  DF3 \u_cordic/mycordic/present_I_table_reg[0][5]  ( .D(\u_cordic/I [2]), .C(
        inClock), .Q(\u_cordic/mycordic/present_I_table[0][5] ), .QN(n45) );
  DF3 \u_cordic/mycordic/present_I_table_reg[0][6]  ( .D(\u_cordic/I [3]), .C(
        inClock), .Q(\u_cordic/mycordic/present_I_table[0][6] ), .QN(n44) );
  DF3 \u_cordic/mycordic/present_I_table_reg[0][7]  ( .D(\u_cordic/I [3]), .C(
        inClock), .Q(\u_cordic/mycordic/present_I_table[0][7] ), .QN(n305) );
  DF3 \u_cordic/my_rotation/present_direction_reg  ( .D(n1529), .C(inClock), 
        .Q(\u_cordic/dir ) );
  DF3 \u_cordic/my_rotation/present_delta_reg[15]  ( .D(n1513), .C(inClock), 
        .Q(\u_cordic/my_rotation/N39 ), .QN(n33) );
  DF3 \u_cordic/my_rotation/present_delta_reg[14]  ( .D(n1514), .C(inClock), 
        .Q(\u_cordic/my_rotation/present_delta [14]), .QN(n267) );
  DF3 \u_cordic/my_rotation/present_delta_reg[13]  ( .D(n1515), .C(inClock), 
        .Q(\u_cordic/my_rotation/present_delta [13]), .QN(n241) );
  DF3 \u_cordic/my_rotation/present_delta_reg[12]  ( .D(n1516), .C(inClock), 
        .Q(\u_cordic/my_rotation/present_delta [12]), .QN(n213) );
  DF3 \u_cordic/my_rotation/present_delta_reg[11]  ( .D(n1517), .C(inClock), 
        .Q(\u_cordic/my_rotation/present_delta [11]), .QN(n179) );
  DF3 \u_cordic/my_rotation/present_delta_reg[10]  ( .D(n1518), .C(inClock), 
        .Q(\u_cordic/my_rotation/present_delta [10]), .QN(n152) );
  DF3 \u_cordic/my_rotation/present_delta_reg[9]  ( .D(n1519), .C(inClock), 
        .Q(\u_cordic/my_rotation/present_delta [9]), .QN(n151) );
  DF3 \u_cordic/my_rotation/present_delta_reg[8]  ( .D(n1520), .C(inClock), 
        .Q(\u_cordic/my_rotation/present_delta [8]) );
  DF3 \u_cordic/my_rotation/present_delta_reg[7]  ( .D(n1521), .C(inClock), 
        .Q(\u_cordic/my_rotation/present_delta [7]), .QN(n123) );
  DF3 \u_cordic/my_rotation/present_delta_reg[6]  ( .D(n1522), .C(inClock), 
        .Q(\u_cordic/my_rotation/present_delta [6]) );
  DF3 \u_cordic/my_rotation/present_delta_reg[5]  ( .D(n1523), .C(inClock), 
        .Q(\u_cordic/my_rotation/present_delta [5]) );
  DF3 \u_cordic/my_rotation/present_delta_reg[4]  ( .D(n1524), .C(inClock), 
        .Q(\u_cordic/my_rotation/present_delta [4]), .QN(n64) );
  DF3 \u_cordic/my_rotation/present_delta_reg[3]  ( .D(n1525), .C(inClock), 
        .Q(\u_cordic/my_rotation/present_delta [3]), .QN(n266) );
  DF3 \u_cordic/my_rotation/present_delta_reg[2]  ( .D(n1526), .C(inClock), 
        .Q(\u_cordic/my_rotation/present_delta [2]) );
  DF3 \u_cordic/my_rotation/present_delta_reg[1]  ( .D(n1527), .C(inClock), 
        .Q(\u_cordic/my_rotation/present_delta [1]) );
  DF3 \u_cordic/my_rotation/present_delta_reg[0]  ( .D(n1528), .C(inClock), 
        .Q(\u_cordic/my_rotation/N41 ) );
  DF3 \u_cordic/my_rotation/present_angle_reg[0][0]  ( .D(n1512), .C(inClock), 
        .Q(\u_cordic/my_rotation/present_angle[0][0] ) );
  DF3 \u_cordic/my_rotation/present_angle_reg[0][1]  ( .D(n1511), .C(inClock), 
        .Q(\u_cordic/my_rotation/present_angle[0][1] ) );
  DF3 \u_cordic/my_rotation/present_angle_reg[0][2]  ( .D(n1510), .C(inClock), 
        .Q(\u_cordic/my_rotation/present_angle[0][2] ) );
  DF3 \u_cordic/my_rotation/present_angle_reg[0][3]  ( .D(n1509), .C(inClock), 
        .Q(\u_cordic/my_rotation/present_angle[0][3] ) );
  DF3 \u_cordic/my_rotation/present_angle_reg[0][4]  ( .D(n1541), .C(inClock), 
        .Q(\u_cordic/my_rotation/present_angle[0][4] ) );
  DF3 \u_cordic/my_rotation/present_angle_reg[0][5]  ( .D(n1540), .C(inClock), 
        .Q(\u_cordic/my_rotation/present_angle[0][5] ) );
  DF3 \u_cordic/my_rotation/present_angle_reg[0][6]  ( .D(n1539), .C(inClock), 
        .Q(\u_cordic/my_rotation/present_angle[0][6] ) );
  DF3 \u_cordic/my_rotation/present_angle_reg[0][7]  ( .D(n1538), .C(inClock), 
        .Q(\u_cordic/my_rotation/present_angle[0][7] ) );
  DF3 \u_cordic/my_rotation/present_angle_reg[0][8]  ( .D(n1537), .C(inClock), 
        .Q(\u_cordic/my_rotation/present_angle[0][8] ) );
  DF3 \u_cordic/my_rotation/present_angle_reg[0][9]  ( .D(n1536), .C(inClock), 
        .Q(\u_cordic/my_rotation/present_angle[0][9] ) );
  DF3 \u_cordic/my_rotation/present_angle_reg[0][10]  ( .D(n1535), .C(inClock), 
        .Q(\u_cordic/my_rotation/present_angle[0][10] ) );
  DF3 \u_cordic/my_rotation/present_angle_reg[0][11]  ( .D(n1534), .C(inClock), 
        .Q(\u_cordic/my_rotation/present_angle[0][11] ) );
  DF3 \u_cordic/my_rotation/present_angle_reg[0][12]  ( .D(n1533), .C(inClock), 
        .Q(\u_cordic/my_rotation/present_angle[0][12] ) );
  DF3 \u_cordic/my_rotation/present_angle_reg[0][13]  ( .D(n1532), .C(inClock), 
        .Q(\u_cordic/my_rotation/present_angle[0][13] ) );
  DF3 \u_cordic/my_rotation/present_angle_reg[0][14]  ( .D(n1531), .C(inClock), 
        .Q(\u_cordic/my_rotation/present_angle[0][14] ) );
  DF3 \u_cordic/my_rotation/present_angle_reg[0][15]  ( .D(n1530), .C(inClock), 
        .Q(\u_cordic/my_rotation/present_angle[0][15] ) );
  DF3 \u_cdr/div1/o_nb_P_reg[2]  ( .D(\u_cdr/div1/n36 ), .C(inClock), .Q(
        \u_cdr/w_nb_P [2]), .QN(\u_cdr/div1/n9 ) );
  DF3 \u_cdr/div1/o_nb_P_reg[1]  ( .D(\u_cdr/div1/n37 ), .C(inClock), .Q(
        \u_cdr/w_nb_P [1]), .QN(\u_cdr/div1/n10 ) );
  DF3 \u_cdr/div1/o_nb_P_reg[3]  ( .D(\u_cdr/div1/n35 ), .C(inClock), .Q(
        \u_cdr/w_nb_P [3]), .QN(\u_cdr/div1/n8 ) );
  DF3 \u_cdr/div1/o_nb_P_reg[4]  ( .D(\u_cdr/div1/n34 ), .C(inClock), .Q(
        \u_cdr/w_nb_P [4]), .QN(n124) );
  DF3 \u_cdr/div1/o_nb_P_reg[5]  ( .D(\u_cdr/div1/n38 ), .C(inClock), .Q(
        \u_cdr/w_nb_P [5]), .QN(\u_cdr/div1/n7 ) );
  DF3 \u_cdr/div1/o_nb_P_reg[0]  ( .D(\u_cdr/div1/n39 ), .C(inClock), .Q(
        \u_cdr/div1/N34 ), .QN(n29) );
  DF3 \u_cdr/phd1/o_T_reg  ( .D(\u_cdr/phd1/n20 ), .C(inClock), .Q(
        \u_cdr/w_sT ), .QN(\u_cdr/phd1/n10 ) );
  DF3 \u_cdr/phd1/o_E_reg  ( .D(\u_cdr/phd1/n21 ), .C(inClock), .Q(
        \u_cdr/w_sE ), .QN(\u_cdr/phd1/n9 ) );
  DF3 \u_cdr/dec1/o_data_reg  ( .D(n1508), .C(inClock), .Q(
        \sig_MUX_inMUX13[0] ), .QN(\u_cdr/dec1/n20 ) );
  DF3 \u_cdr/dec1/o_flag_reg  ( .D(\u_cdr/dec1/N73 ), .C(inClock), .Q(
        \sig_MUX_inMUX12[0] ), .QN(n40) );
  DF3 \u_cdr/dec1/cnt_r_reg[1]  ( .D(n1163), .C(inClock), .Q(
        \u_cdr/dec1/cnt_r [1]) );
  DF3 \u_cdr/dec1/cnt_r_reg[2]  ( .D(n1164), .C(inClock), .Q(
        \u_cdr/dec1/cnt_r [2]) );
  DF3 \u_cdr/dec1/cnt_r_reg[3]  ( .D(n1165), .C(inClock), .Q(
        \u_cdr/dec1/cnt_r [3]) );
  DF3 \u_cdr/dec1/cnt_r_reg[4]  ( .D(n1166), .C(inClock), .Q(
        \u_cdr/dec1/cnt_r [4]) );
  DF3 \u_cdr/dec1/cnt_r_reg[5]  ( .D(n1162), .C(inClock), .Q(
        \u_cdr/dec1/cnt_r [5]), .QN(n304) );
  DF3 \u_cdr/dec1/cnt_r_reg[0]  ( .D(n1161), .C(inClock), .Q(
        \u_cdr/dec1/cnt_r [0]), .QN(n250) );
  DF3 \u_inFIFO/os1/dff1/s_qout_reg  ( .D(n1507), .C(inClock), .Q(
        \u_inFIFO/os1/sigQout1 ), .QN(n293) );
  DF3 \u_decoder/iq_demod/cossin_dig/o_cos_reg[0]  ( .D(n2243), .C(inClock), 
        .Q(\u_decoder/iq_demod/cos_out [0]), .QN(n27) );
  DF3 \u_decoder/iq_demod/cossin_dig/o_cos_reg[1]  ( .D(
        \u_decoder/iq_demod/cossin_dig/n49 ), .C(inClock), .Q(
        \u_decoder/iq_demod/cos_out [1]), .QN(n23) );
  DF3 \u_decoder/iq_demod/cossin_dig/o_cos_reg[2]  ( .D(
        \u_decoder/iq_demod/cossin_dig/n50 ), .C(inClock), .Q(
        \u_decoder/iq_demod/cos_out [2]), .QN(n25) );
  DF3 \u_decoder/iq_demod/cossin_dig/o_cos_reg[3]  ( .D(n2244), .C(inClock), 
        .Q(\u_decoder/iq_demod/cos_out [3]), .QN(n5) );
  DF3 \u_decoder/iq_demod/cossin_dig/o_sin_reg[0]  ( .D(
        \u_decoder/iq_demod/cossin_dig/n51 ), .C(inClock), .Q(
        \u_decoder/iq_demod/sin_out [0]), .QN(n24) );
  DF3 \u_decoder/iq_demod/cossin_dig/o_sin_reg[1]  ( .D(n2245), .C(inClock), 
        .Q(\u_decoder/iq_demod/sin_out [1]), .QN(n26) );
  DF3 \u_decoder/iq_demod/cossin_dig/o_sin_reg[2]  ( .D(n2246), .C(inClock), 
        .Q(\u_decoder/iq_demod/sin_out [2]), .QN(n28) );
  DF3 \u_decoder/iq_demod/cossin_dig/o_sin_reg[3]  ( .D(n2247), .C(inClock), 
        .Q(\u_decoder/iq_demod/sin_out [3]), .QN(n6) );
  DF3 \u_decoder/iq_demod/cossin_dig/val_counter_reg[2]  ( .D(n1505), .C(
        inClock), .Q(\u_decoder/iq_demod/cossin_dig/val_counter [2]) );
  DF3 \u_decoder/iq_demod/cossin_dig/val_counter_reg[1]  ( .D(
        \u_decoder/iq_demod/cossin_dig/n52 ), .C(inClock), .Q(
        \u_decoder/iq_demod/cossin_dig/val_counter [1]), .QN(
        \u_decoder/iq_demod/cossin_dig/n19 ) );
  DF3 \u_decoder/iq_demod/cossin_dig/val_counter_reg[0]  ( .D(
        \u_decoder/iq_demod/cossin_dig/n53 ), .C(inClock), .Q(
        \u_decoder/iq_demod/cossin_dig/N55 ), .QN(
        \u_decoder/iq_demod/cossin_dig/n21 ) );
  DF3 \u_decoder/iq_demod/cossin_dig/state_reg[1]  ( .D(
        \u_decoder/iq_demod/cossin_dig/N42 ), .C(inClock), .QN(
        \u_decoder/iq_demod/cossin_dig/n23 ) );
  DF3 \u_decoder/iq_demod/cossin_dig/counter_reg[2]  ( .D(
        \u_decoder/iq_demod/cossin_dig/N22 ), .C(inClock), .Q(
        \u_decoder/iq_demod/cossin_dig/counter [2]), .QN(
        \u_decoder/iq_demod/cossin_dig/n10 ) );
  DF3 \u_decoder/iq_demod/cossin_dig/counter_reg[1]  ( .D(
        \u_decoder/iq_demod/cossin_dig/N21 ), .C(inClock), .Q(
        \u_decoder/iq_demod/cossin_dig/counter [1]) );
  DF3 \u_decoder/iq_demod/cossin_dig/counter_reg[0]  ( .D(
        \u_decoder/iq_demod/cossin_dig/N20 ), .C(inClock), .Q(
        \u_decoder/iq_demod/cossin_dig/counter [0]) );
  DF3 \u_decoder/iq_demod/cossin_dig/state_reg[0]  ( .D(
        \u_decoder/iq_demod/cossin_dig/N41 ), .C(inClock), .Q(
        \u_decoder/iq_demod/cossin_dig/state[0] ) );
  DF3 \u_cdr/div1/cnt_div/o_en_freq_synch_reg  ( .D(n1503), .C(inClock), .Q(
        \u_cdr/div1/w_en_freq_synch ) );
  DF3 \u_cdr/div1/cnt_div/cnt_reg[1]  ( .D(n1157), .C(inClock), .Q(
        \u_cdr/div1/cnt_div/cnt [1]) );
  DF3 \u_cdr/div1/cnt_div/cnt_reg[2]  ( .D(n1158), .C(inClock), .Q(
        \u_cdr/div1/cnt_div/cnt [2]) );
  DF3 \u_cdr/div1/cnt_div/cnt_reg[3]  ( .D(n1159), .C(inClock), .Q(
        \u_cdr/div1/cnt_div/cnt [3]) );
  DF3 \u_cdr/div1/cnt_div/cnt_reg[4]  ( .D(n1160), .C(inClock), .Q(
        \u_cdr/div1/cnt_div/cnt [4]) );
  DF3 \u_cdr/div1/cnt_div/cnt_reg[5]  ( .D(n1156), .C(inClock), .Q(
        \u_cdr/div1/cnt_div/cnt [5]) );
  DF3 \u_cdr/div1/cnt_div/cnt_reg[0]  ( .D(n1155), .C(inClock), .Q(
        \u_cdr/div1/cnt_div/cnt [0]), .QN(n197) );
  DF3 \u_cdr/phd1/f1/o_Q_reg  ( .D(n1502), .C(inClock), .Q(\u_cdr/phd1/w_s1 )
         );
  DF3 \u_outFIFO/os2/dff2/s_qout_reg  ( .D(n1501), .C(inClock), .Q(
        \u_outFIFO/os2/sigQout2 ) );
  DF3 \u_outFIFO/os2/dff1/s_qout_reg  ( .D(n1500), .C(inClock), .Q(
        \u_outFIFO/os2/sigQout1 ), .QN(n291) );
  DF3 \u_outFIFO/os1/dff2/s_qout_reg  ( .D(n1499), .C(inClock), .Q(
        \u_outFIFO/os1/sigQout2 ) );
  DF3 \u_outFIFO/os1/dff1/s_qout_reg  ( .D(n1498), .C(inClock), .Q(
        \u_outFIFO/os1/sigQout1 ), .QN(n292) );
  DF3 \u_inFIFO/os2/dff2/s_qout_reg  ( .D(n1497), .C(inClock), .Q(
        \u_inFIFO/os2/sigQout2 ) );
  DF3 \u_inFIFO/os2/dff1/s_qout_reg  ( .D(n1496), .C(inClock), .Q(
        \u_inFIFO/os2/sigQout1 ), .QN(n290) );
  DF3 \u_inFIFO/os1/dff2/s_qout_reg  ( .D(n1495), .C(inClock), .Q(
        \u_inFIFO/os1/sigQout2 ) );
  DF3 \u_cdr/dec1/cnt_dec/o_en_dec_reg  ( .D(n1494), .C(inClock), .Q(
        \u_cdr/dec1/w_en_dec ), .QN(n308) );
  DF3 \u_cdr/dec1/cnt_dec/cnt_reg[1]  ( .D(n1151), .C(inClock), .Q(
        \u_cdr/dec1/cnt_dec/cnt [1]), .QN(n278) );
  DF3 \u_cdr/dec1/cnt_dec/cnt_reg[2]  ( .D(n1152), .C(inClock), .Q(
        \u_cdr/dec1/cnt_dec/cnt [2]) );
  DF3 \u_cdr/dec1/cnt_dec/cnt_reg[3]  ( .D(n1153), .C(inClock), .Q(
        \u_cdr/dec1/cnt_dec/cnt [3]) );
  DF3 \u_cdr/dec1/cnt_dec/cnt_reg[4]  ( .D(n1154), .C(inClock), .Q(
        \u_cdr/dec1/cnt_dec/cnt [4]) );
  DF3 \u_cdr/dec1/cnt_dec/cnt_reg[5]  ( .D(n1150), .C(inClock), .Q(
        \u_cdr/dec1/cnt_dec/cnt [5]) );
  DF3 \u_cdr/dec1/cnt_dec/cnt_reg[0]  ( .D(n1149), .C(inClock), .Q(
        \u_cdr/dec1/cnt_dec/cnt [0]), .QN(n196) );
  DF3 \u_cdr/phd1/cnt_phd/o_en_reg  ( .D(n1491), .C(inClock), .QN(n312) );
  DF3 \u_cdr/phd1/cnt_phd/o_en_f_reg  ( .D(n1492), .C(inClock), .Q(
        \u_cdr/phd1/w_en_f ), .QN(n302) );
  DF3 \u_cdr/phd1/cnt_phd/o_en_m_reg  ( .D(n1493), .C(inClock), .Q(
        \u_cdr/phd1/w_en_m ), .QN(n313) );
  DF3 \u_cdr/phd1/cnt_phd/o_en_d_reg  ( .D(\u_cdr/phd1/cnt_phd/N92 ), .C(
        inClock), .Q(\u_cdr/phd1/w_en_d ) );
  DF3 \u_cdr/phd1/cnt_phd/cnt_reg[1]  ( .D(n1145), .C(inClock), .Q(
        \u_cdr/phd1/cnt_phd/cnt [1]), .QN(n276) );
  DF3 \u_cdr/phd1/cnt_phd/cnt_reg[2]  ( .D(n1146), .C(inClock), .Q(
        \u_cdr/phd1/cnt_phd/cnt [2]) );
  DF3 \u_cdr/phd1/cnt_phd/cnt_reg[3]  ( .D(n1147), .C(inClock), .Q(
        \u_cdr/phd1/cnt_phd/cnt [3]) );
  DF3 \u_cdr/phd1/cnt_phd/cnt_reg[4]  ( .D(n1148), .C(inClock), .Q(
        \u_cdr/phd1/cnt_phd/cnt [4]) );
  DF3 \u_cdr/phd1/cnt_phd/cnt_reg[5]  ( .D(n1144), .C(inClock), .Q(
        \u_cdr/phd1/cnt_phd/cnt [5]), .QN(n271) );
  DF3 \u_cdr/phd1/cnt_phd/cnt_reg[0]  ( .D(n1143), .C(inClock), .Q(
        \u_cdr/phd1/cnt_phd/cnt [0]), .QN(n2620) );
  DF3 \u_cdr/dec1/ffd_retard/o_Q_reg  ( .D(n1490), .C(inClock), .Q(
        \u_cdr/dec1/w_s_r ), .QN(n289) );
  DF3 \u_cdr/phd1/f4/o_Q_reg  ( .D(n1489), .C(inClock), .Q(\u_cdr/phd1/w_s4 )
         );
  DF3 \u_cdr/phd1/f3/o_Q_reg  ( .D(n1488), .C(inClock), .Q(\u_cdr/phd1/w_s3 )
         );
  DF3 \u_cdr/phd1/f2/o_Q_reg  ( .D(n1487), .C(inClock), .Q(\u_cdr/phd1/w_s2 )
         );
  DFE1 \u_cdr/dir_f_reg  ( .D(n1586), .E(\u_cdr/n44 ), .C(inClock), .QN(
        \u_cdr/n3 ) );
  DFE1 \u_cdr/dir_d_reg  ( .D(n1586), .E(\u_cdr/n30 ), .C(inClock), .QN(
        \u_cdr/n18 ) );
  DFE1 \u_cdr/dir_m_reg  ( .D(n1586), .E(\u_cdr/n27 ), .C(inClock), .QN(
        \u_cdr/n19 ) );
  DFE1 \u_cordic/my_rotation/present_angle_reg[1][14]  ( .D(
        \u_cordic/my_rotation/present_angle[0][14] ), .E(n979), .C(inClock), 
        .QN(n296) );
  DFE1 \u_cordic/my_rotation/present_angle_reg[1][15]  ( .D(
        \u_cordic/my_rotation/present_angle[0][15] ), .E(n978), .C(inClock), 
        .QN(n309) );
  DFE1 \u_inFIFO/FIFO_reg[2][0]  ( .D(n1611), .E(n1649), .C(inClock), .Q(
        \u_inFIFO/FIFO[2][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[2][1]  ( .D(n1612), .E(n1649), .C(inClock), .Q(
        \u_inFIFO/FIFO[2][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[2][2]  ( .D(n1613), .E(n1649), .C(inClock), .Q(
        \u_inFIFO/FIFO[2][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[2][3]  ( .D(n1614), .E(n1649), .C(inClock), .Q(
        \u_inFIFO/FIFO[2][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[6][0]  ( .D(n1611), .E(n1645), .C(inClock), .Q(
        \u_inFIFO/FIFO[6][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[6][1]  ( .D(n1612), .E(n1645), .C(inClock), .Q(
        \u_inFIFO/FIFO[6][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[6][2]  ( .D(n1613), .E(n1645), .C(inClock), .Q(
        \u_inFIFO/FIFO[6][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[6][3]  ( .D(n1614), .E(n1645), .C(inClock), .Q(
        \u_inFIFO/FIFO[6][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[10][0]  ( .D(n1611), .E(n1641), .C(inClock), .Q(
        \u_inFIFO/FIFO[10][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[10][1]  ( .D(n1612), .E(n1641), .C(inClock), .Q(
        \u_inFIFO/FIFO[10][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[10][2]  ( .D(n1613), .E(n1641), .C(inClock), .Q(
        \u_inFIFO/FIFO[10][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[10][3]  ( .D(n1614), .E(n1641), .C(inClock), .Q(
        \u_inFIFO/FIFO[10][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[14][0]  ( .D(n1611), .E(n1637), .C(inClock), .Q(
        \u_inFIFO/FIFO[14][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[14][1]  ( .D(n1612), .E(n1637), .C(inClock), .Q(
        \u_inFIFO/FIFO[14][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[14][2]  ( .D(n1613), .E(n1637), .C(inClock), .Q(
        \u_inFIFO/FIFO[14][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[14][3]  ( .D(n1614), .E(n1637), .C(inClock), .Q(
        \u_inFIFO/FIFO[14][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[18][0]  ( .D(n1611), .E(n1633), .C(inClock), .Q(
        \u_inFIFO/FIFO[18][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[18][1]  ( .D(n1612), .E(n1633), .C(inClock), .Q(
        \u_inFIFO/FIFO[18][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[18][2]  ( .D(n1613), .E(n1633), .C(inClock), .Q(
        \u_inFIFO/FIFO[18][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[18][3]  ( .D(n1614), .E(n1633), .C(inClock), .Q(
        \u_inFIFO/FIFO[18][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[22][0]  ( .D(n1611), .E(n1629), .C(inClock), .Q(
        \u_inFIFO/FIFO[22][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[22][1]  ( .D(n1612), .E(n1629), .C(inClock), .Q(
        \u_inFIFO/FIFO[22][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[22][2]  ( .D(n1613), .E(n1629), .C(inClock), .Q(
        \u_inFIFO/FIFO[22][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[22][3]  ( .D(n1614), .E(n1629), .C(inClock), .Q(
        \u_inFIFO/FIFO[22][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[26][0]  ( .D(n1611), .E(n1625), .C(inClock), .Q(
        \u_inFIFO/FIFO[26][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[26][1]  ( .D(n1612), .E(n1625), .C(inClock), .Q(
        \u_inFIFO/FIFO[26][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[26][2]  ( .D(n1613), .E(n1625), .C(inClock), .Q(
        \u_inFIFO/FIFO[26][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[26][3]  ( .D(n1614), .E(n1625), .C(inClock), .Q(
        \u_inFIFO/FIFO[26][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[30][0]  ( .D(n1611), .E(n1621), .C(inClock), .Q(
        \u_inFIFO/FIFO[30][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[30][1]  ( .D(n1612), .E(n1621), .C(inClock), .Q(
        \u_inFIFO/FIFO[30][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[30][2]  ( .D(n1613), .E(n1621), .C(inClock), .Q(
        \u_inFIFO/FIFO[30][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[30][3]  ( .D(n1614), .E(n1621), .C(inClock), .Q(
        \u_inFIFO/FIFO[30][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[0][0]  ( .D(n1611), .E(n1651), .C(inClock), .Q(
        \u_inFIFO/FIFO[0][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[0][1]  ( .D(n1612), .E(n1651), .C(inClock), .Q(
        \u_inFIFO/FIFO[0][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[0][2]  ( .D(n1613), .E(n1651), .C(inClock), .Q(
        \u_inFIFO/FIFO[0][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[0][3]  ( .D(n1614), .E(n1651), .C(inClock), .Q(
        \u_inFIFO/FIFO[0][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[1][0]  ( .D(n1611), .E(n1650), .C(inClock), .Q(
        \u_inFIFO/FIFO[1][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[1][1]  ( .D(n1612), .E(n1650), .C(inClock), .Q(
        \u_inFIFO/FIFO[1][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[1][2]  ( .D(n1613), .E(n1650), .C(inClock), .Q(
        \u_inFIFO/FIFO[1][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[1][3]  ( .D(n1614), .E(n1650), .C(inClock), .Q(
        \u_inFIFO/FIFO[1][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[3][0]  ( .D(n1611), .E(n1648), .C(inClock), .Q(
        \u_inFIFO/FIFO[3][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[3][1]  ( .D(n1612), .E(n1648), .C(inClock), .Q(
        \u_inFIFO/FIFO[3][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[3][2]  ( .D(n1613), .E(n1648), .C(inClock), .Q(
        \u_inFIFO/FIFO[3][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[3][3]  ( .D(n1614), .E(n1648), .C(inClock), .Q(
        \u_inFIFO/FIFO[3][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[4][0]  ( .D(n1611), .E(n1647), .C(inClock), .Q(
        \u_inFIFO/FIFO[4][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[4][1]  ( .D(n1612), .E(n1647), .C(inClock), .Q(
        \u_inFIFO/FIFO[4][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[4][2]  ( .D(n1613), .E(n1647), .C(inClock), .Q(
        \u_inFIFO/FIFO[4][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[4][3]  ( .D(n1614), .E(n1647), .C(inClock), .Q(
        \u_inFIFO/FIFO[4][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[5][0]  ( .D(n1611), .E(n1646), .C(inClock), .Q(
        \u_inFIFO/FIFO[5][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[5][1]  ( .D(n1612), .E(n1646), .C(inClock), .Q(
        \u_inFIFO/FIFO[5][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[5][2]  ( .D(n1613), .E(n1646), .C(inClock), .Q(
        \u_inFIFO/FIFO[5][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[5][3]  ( .D(n1614), .E(n1646), .C(inClock), .Q(
        \u_inFIFO/FIFO[5][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[7][0]  ( .D(n1611), .E(n1644), .C(inClock), .Q(
        \u_inFIFO/FIFO[7][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[7][1]  ( .D(n1612), .E(n1644), .C(inClock), .Q(
        \u_inFIFO/FIFO[7][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[7][2]  ( .D(n1613), .E(n1644), .C(inClock), .Q(
        \u_inFIFO/FIFO[7][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[7][3]  ( .D(n1614), .E(n1644), .C(inClock), .Q(
        \u_inFIFO/FIFO[7][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[8][0]  ( .D(n1611), .E(n1643), .C(inClock), .Q(
        \u_inFIFO/FIFO[8][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[8][1]  ( .D(n1612), .E(n1643), .C(inClock), .Q(
        \u_inFIFO/FIFO[8][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[8][2]  ( .D(n1613), .E(n1643), .C(inClock), .Q(
        \u_inFIFO/FIFO[8][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[8][3]  ( .D(n1614), .E(n1643), .C(inClock), .Q(
        \u_inFIFO/FIFO[8][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[9][0]  ( .D(n1611), .E(n1642), .C(inClock), .Q(
        \u_inFIFO/FIFO[9][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[9][1]  ( .D(n1612), .E(n1642), .C(inClock), .Q(
        \u_inFIFO/FIFO[9][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[9][2]  ( .D(n1613), .E(n1642), .C(inClock), .Q(
        \u_inFIFO/FIFO[9][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[9][3]  ( .D(n1614), .E(n1642), .C(inClock), .Q(
        \u_inFIFO/FIFO[9][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[11][0]  ( .D(n1611), .E(n1640), .C(inClock), .Q(
        \u_inFIFO/FIFO[11][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[11][1]  ( .D(n1612), .E(n1640), .C(inClock), .Q(
        \u_inFIFO/FIFO[11][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[11][2]  ( .D(n1613), .E(n1640), .C(inClock), .Q(
        \u_inFIFO/FIFO[11][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[11][3]  ( .D(n1614), .E(n1640), .C(inClock), .Q(
        \u_inFIFO/FIFO[11][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[12][0]  ( .D(n1611), .E(n1639), .C(inClock), .Q(
        \u_inFIFO/FIFO[12][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[12][1]  ( .D(n1612), .E(n1639), .C(inClock), .Q(
        \u_inFIFO/FIFO[12][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[12][2]  ( .D(n1613), .E(n1639), .C(inClock), .Q(
        \u_inFIFO/FIFO[12][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[12][3]  ( .D(n1614), .E(n1639), .C(inClock), .Q(
        \u_inFIFO/FIFO[12][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[13][0]  ( .D(n1611), .E(n1638), .C(inClock), .Q(
        \u_inFIFO/FIFO[13][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[13][1]  ( .D(n1612), .E(n1638), .C(inClock), .Q(
        \u_inFIFO/FIFO[13][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[13][2]  ( .D(n1613), .E(n1638), .C(inClock), .Q(
        \u_inFIFO/FIFO[13][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[13][3]  ( .D(n1614), .E(n1638), .C(inClock), .Q(
        \u_inFIFO/FIFO[13][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[15][0]  ( .D(n1611), .E(n1636), .C(inClock), .Q(
        \u_inFIFO/FIFO[15][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[15][1]  ( .D(n1612), .E(n1636), .C(inClock), .Q(
        \u_inFIFO/FIFO[15][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[15][2]  ( .D(n1613), .E(n1636), .C(inClock), .Q(
        \u_inFIFO/FIFO[15][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[15][3]  ( .D(n1614), .E(n1636), .C(inClock), .Q(
        \u_inFIFO/FIFO[15][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[16][0]  ( .D(n1611), .E(n1635), .C(inClock), .Q(
        \u_inFIFO/FIFO[16][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[16][1]  ( .D(n1612), .E(n1635), .C(inClock), .Q(
        \u_inFIFO/FIFO[16][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[16][2]  ( .D(n1613), .E(n1635), .C(inClock), .Q(
        \u_inFIFO/FIFO[16][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[16][3]  ( .D(n1614), .E(n1635), .C(inClock), .Q(
        \u_inFIFO/FIFO[16][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[17][0]  ( .D(n1611), .E(n1634), .C(inClock), .Q(
        \u_inFIFO/FIFO[17][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[17][1]  ( .D(n1612), .E(n1634), .C(inClock), .Q(
        \u_inFIFO/FIFO[17][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[17][2]  ( .D(n1613), .E(n1634), .C(inClock), .Q(
        \u_inFIFO/FIFO[17][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[17][3]  ( .D(n1614), .E(n1634), .C(inClock), .Q(
        \u_inFIFO/FIFO[17][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[19][0]  ( .D(n1611), .E(n1632), .C(inClock), .Q(
        \u_inFIFO/FIFO[19][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[19][1]  ( .D(n1612), .E(n1632), .C(inClock), .Q(
        \u_inFIFO/FIFO[19][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[19][2]  ( .D(n1613), .E(n1632), .C(inClock), .Q(
        \u_inFIFO/FIFO[19][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[19][3]  ( .D(n1614), .E(n1632), .C(inClock), .Q(
        \u_inFIFO/FIFO[19][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[20][0]  ( .D(n1611), .E(n1631), .C(inClock), .Q(
        \u_inFIFO/FIFO[20][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[20][1]  ( .D(n1612), .E(n1631), .C(inClock), .Q(
        \u_inFIFO/FIFO[20][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[20][2]  ( .D(n1613), .E(n1631), .C(inClock), .Q(
        \u_inFIFO/FIFO[20][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[20][3]  ( .D(n1614), .E(n1631), .C(inClock), .Q(
        \u_inFIFO/FIFO[20][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[21][0]  ( .D(n1611), .E(n1630), .C(inClock), .Q(
        \u_inFIFO/FIFO[21][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[21][1]  ( .D(n1612), .E(n1630), .C(inClock), .Q(
        \u_inFIFO/FIFO[21][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[21][2]  ( .D(n1613), .E(n1630), .C(inClock), .Q(
        \u_inFIFO/FIFO[21][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[21][3]  ( .D(n1614), .E(n1630), .C(inClock), .Q(
        \u_inFIFO/FIFO[21][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[23][0]  ( .D(n1611), .E(n1628), .C(inClock), .Q(
        \u_inFIFO/FIFO[23][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[23][1]  ( .D(n1612), .E(n1628), .C(inClock), .Q(
        \u_inFIFO/FIFO[23][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[23][2]  ( .D(n1613), .E(n1628), .C(inClock), .Q(
        \u_inFIFO/FIFO[23][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[23][3]  ( .D(n1614), .E(n1628), .C(inClock), .Q(
        \u_inFIFO/FIFO[23][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[24][0]  ( .D(n1611), .E(n1627), .C(inClock), .Q(
        \u_inFIFO/FIFO[24][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[24][1]  ( .D(n1612), .E(n1627), .C(inClock), .Q(
        \u_inFIFO/FIFO[24][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[24][2]  ( .D(n1613), .E(n1627), .C(inClock), .Q(
        \u_inFIFO/FIFO[24][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[24][3]  ( .D(n1614), .E(n1627), .C(inClock), .Q(
        \u_inFIFO/FIFO[24][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[25][0]  ( .D(n1611), .E(n1626), .C(inClock), .Q(
        \u_inFIFO/FIFO[25][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[25][1]  ( .D(n1612), .E(n1626), .C(inClock), .Q(
        \u_inFIFO/FIFO[25][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[25][2]  ( .D(n1613), .E(n1626), .C(inClock), .Q(
        \u_inFIFO/FIFO[25][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[25][3]  ( .D(n1614), .E(n1626), .C(inClock), .Q(
        \u_inFIFO/FIFO[25][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[27][0]  ( .D(n1611), .E(n1624), .C(inClock), .Q(
        \u_inFIFO/FIFO[27][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[27][1]  ( .D(n1612), .E(n1624), .C(inClock), .Q(
        \u_inFIFO/FIFO[27][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[27][2]  ( .D(n1613), .E(n1624), .C(inClock), .Q(
        \u_inFIFO/FIFO[27][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[27][3]  ( .D(n1614), .E(n1624), .C(inClock), .Q(
        \u_inFIFO/FIFO[27][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[28][0]  ( .D(n1611), .E(n1623), .C(inClock), .Q(
        \u_inFIFO/FIFO[28][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[28][1]  ( .D(n1612), .E(n1623), .C(inClock), .Q(
        \u_inFIFO/FIFO[28][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[28][2]  ( .D(n1613), .E(n1623), .C(inClock), .Q(
        \u_inFIFO/FIFO[28][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[28][3]  ( .D(n1614), .E(n1623), .C(inClock), .Q(
        \u_inFIFO/FIFO[28][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[29][0]  ( .D(n1611), .E(n1622), .C(inClock), .Q(
        \u_inFIFO/FIFO[29][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[29][1]  ( .D(n1612), .E(n1622), .C(inClock), .Q(
        \u_inFIFO/FIFO[29][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[29][2]  ( .D(n1613), .E(n1622), .C(inClock), .Q(
        \u_inFIFO/FIFO[29][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[29][3]  ( .D(n1614), .E(n1622), .C(inClock), .Q(
        \u_inFIFO/FIFO[29][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[31][0]  ( .D(n1611), .E(n1620), .C(inClock), .Q(
        \u_inFIFO/FIFO[31][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[31][1]  ( .D(n1612), .E(n1620), .C(inClock), .Q(
        \u_inFIFO/FIFO[31][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[31][2]  ( .D(n1613), .E(n1620), .C(inClock), .Q(
        \u_inFIFO/FIFO[31][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[31][3]  ( .D(n1614), .E(n1620), .C(inClock), .Q(
        \u_inFIFO/FIFO[31][3] ) );
  DFE1 \u_cordic/my_rotation/present_angle_reg[1][13]  ( .D(
        \u_cordic/my_rotation/present_angle[0][13] ), .E(n978), .C(inClock), 
        .QN(n275) );
  DFE1 \u_cordic/my_rotation/present_angle_reg[1][11]  ( .D(
        \u_cordic/my_rotation/present_angle[0][11] ), .E(n979), .C(inClock), 
        .QN(n256) );
  DFE1 \u_cordic/my_rotation/present_angle_reg[1][12]  ( .D(
        \u_cordic/my_rotation/present_angle[0][12] ), .E(n978), .C(inClock), 
        .QN(n255) );
  DFE1 \u_coder/my_clk_10M_reg  ( .D(\u_coder/clk_10M ), .E(n979), .C(inClock), 
        .Q(\u_coder/my_clk_10M ), .QN(\u_coder/n69 ) );
  DFE1 \u_cordic/my_rotation/present_angle_reg[1][10]  ( .D(
        \u_cordic/my_rotation/present_angle[0][10] ), .E(n979), .C(inClock), 
        .QN(n228) );
  DFE1 \u_cordic/my_rotation/present_angle_reg[1][8]  ( .D(
        \u_cordic/my_rotation/present_angle[0][8] ), .E(n979), .C(inClock), 
        .QN(n195) );
  DFE1 \u_cordic/my_rotation/present_angle_reg[1][9]  ( .D(
        \u_cordic/my_rotation/present_angle[0][9] ), .E(n979), .C(inClock), 
        .QN(n194) );
  DFE1 \u_cordic/my_rotation/present_angle_reg[1][7]  ( .D(
        \u_cordic/my_rotation/present_angle[0][7] ), .E(n979), .C(inClock), 
        .QN(n163) );
  DFE1 \u_cordic/my_rotation/present_angle_reg[1][5]  ( .D(
        \u_cordic/my_rotation/present_angle[0][5] ), .E(n979), .C(inClock), 
        .QN(n141) );
  DFE1 \u_cordic/my_rotation/present_angle_reg[1][6]  ( .D(
        \u_cordic/my_rotation/present_angle[0][6] ), .E(n979), .C(inClock), 
        .QN(n140) );
  DFE1 \u_cordic/my_rotation/present_angle_reg[1][4]  ( .D(
        \u_cordic/my_rotation/present_angle[0][4] ), .E(n979), .C(inClock), 
        .QN(n127) );
  DFE1 \u_cordic/my_rotation/present_angle_reg[1][2]  ( .D(
        \u_cordic/my_rotation/present_angle[0][2] ), .E(n979), .C(inClock), 
        .QN(n111) );
  DFE1 \u_cordic/my_rotation/present_angle_reg[1][3]  ( .D(
        \u_cordic/my_rotation/present_angle[0][3] ), .E(n979), .C(inClock), 
        .QN(n110) );
  DFE1 \u_cordic/my_rotation/present_angle_reg[1][0]  ( .D(
        \u_cordic/my_rotation/present_angle[0][0] ), .E(n979), .C(inClock), 
        .QN(n61) );
  DFE1 \u_cordic/my_rotation/present_angle_reg[1][1]  ( .D(
        \u_cordic/my_rotation/present_angle[0][1] ), .E(n979), .C(inClock), 
        .QN(n68) );
  NOR21 \u_decoder/iq_demod/cossin_dig/U49  ( .A(
        \u_decoder/iq_demod/cossin_dig/n21 ), .B(
        \u_decoder/iq_demod/cossin_dig/n19 ), .Q(
        \u_decoder/iq_demod/cossin_dig/N52 ) );
  NAND22 \u_cordic/mycordic/U560  ( .A(n303), .B(n751), .Q(
        \u_cordic/mycordic/n562 ) );
  NAND22 \u_cordic/mycordic/U558  ( .A(
        \u_cordic/mycordic/present_ANGLE_table[6][1] ), .B(n751), .Q(
        \u_cordic/mycordic/n558 ) );
  NAND22 \u_cordic/mycordic/U557  ( .A(\u_cordic/mycordic/N615 ), .B(n751), 
        .Q(\u_cordic/mycordic/n556 ) );
  NAND22 \u_cordic/mycordic/U559  ( .A(
        \u_cordic/mycordic/present_ANGLE_table[6][2] ), .B(n751), .Q(
        \u_cordic/mycordic/n560 ) );
  NAND22 \u_decoder/iq_demod/cossin_dig/U50  ( .A(
        \u_decoder/iq_demod/cossin_dig/N55 ), .B(
        \u_decoder/iq_demod/cossin_dig/n19 ), .Q(
        \u_decoder/iq_demod/cossin_dig/n55 ) );
  NOR21 \u_decoder/iq_demod/cossin_dig/U51  ( .A(
        \u_decoder/iq_demod/cossin_dig/N55 ), .B(
        \u_decoder/iq_demod/cossin_dig/n54 ), .Q(
        \u_decoder/iq_demod/cossin_dig/N60 ) );
  NAND22 \u_cordic/mycordic/U562  ( .A(\u_cordic/mycordic/N620 ), .B(n751), 
        .Q(\u_cordic/mycordic/n566 ) );
  NAND22 \u_cordic/mycordic/U561  ( .A(\u_cordic/mycordic/N619 ), .B(n751), 
        .Q(\u_cordic/mycordic/n564 ) );
  NAND22 \u_decoder/iq_demod/cossin_dig/U52  ( .A(
        \u_decoder/iq_demod/cossin_dig/n21 ), .B(
        \u_decoder/iq_demod/cossin_dig/n54 ), .Q(
        \u_decoder/iq_demod/cossin_dig/n56 ) );
  IMUX40 \u_outFIFO/U685  ( .A(\u_outFIFO/FIFO[4][0] ), .B(
        \u_outFIFO/FIFO[5][0] ), .C(\u_outFIFO/FIFO[6][0] ), .D(
        \u_outFIFO/FIFO[7][0] ), .S0(n35), .S1(\u_outFIFO/N36 ), .Q(
        \u_outFIFO/n700 ) );
  IMUX40 \u_outFIFO/U693  ( .A(\u_outFIFO/FIFO[4][1] ), .B(
        \u_outFIFO/FIFO[5][1] ), .C(\u_outFIFO/FIFO[6][1] ), .D(
        \u_outFIFO/FIFO[7][1] ), .S0(n35), .S1(\u_outFIFO/N36 ), .Q(
        \u_outFIFO/n710 ) );
  IMUX40 \u_outFIFO/U701  ( .A(\u_outFIFO/FIFO[4][2] ), .B(
        \u_outFIFO/FIFO[5][2] ), .C(\u_outFIFO/FIFO[6][2] ), .D(
        \u_outFIFO/FIFO[7][2] ), .S0(n942), .S1(\u_outFIFO/N36 ), .Q(
        \u_outFIFO/n720 ) );
  IMUX40 \u_outFIFO/U709  ( .A(\u_outFIFO/FIFO[4][3] ), .B(
        \u_outFIFO/FIFO[5][3] ), .C(\u_outFIFO/FIFO[6][3] ), .D(
        \u_outFIFO/FIFO[7][3] ), .S0(n942), .S1(\u_outFIFO/N36 ), .Q(
        \u_outFIFO/n730 ) );
  IMUX40 \u_outFIFO/U684  ( .A(\u_outFIFO/FIFO[8][0] ), .B(
        \u_outFIFO/FIFO[9][0] ), .C(\u_outFIFO/FIFO[10][0] ), .D(
        \u_outFIFO/FIFO[11][0] ), .S0(n35), .S1(\u_outFIFO/N36 ), .Q(
        \u_outFIFO/n699 ) );
  IMUX40 \u_outFIFO/U686  ( .A(\u_outFIFO/FIFO[0][0] ), .B(
        \u_outFIFO/FIFO[1][0] ), .C(\u_outFIFO/FIFO[2][0] ), .D(
        \u_outFIFO/FIFO[3][0] ), .S0(n35), .S1(\u_outFIFO/N36 ), .Q(
        \u_outFIFO/n698 ) );
  IMUX40 \u_outFIFO/U683  ( .A(\u_outFIFO/FIFO[12][0] ), .B(
        \u_outFIFO/FIFO[13][0] ), .C(\u_outFIFO/FIFO[14][0] ), .D(
        \u_outFIFO/FIFO[15][0] ), .S0(n35), .S1(\u_outFIFO/N36 ), .Q(
        \u_outFIFO/n701 ) );
  IMUX40 \u_outFIFO/U679  ( .A(\u_outFIFO/FIFO[28][0] ), .B(
        \u_outFIFO/FIFO[29][0] ), .C(\u_outFIFO/FIFO[30][0] ), .D(
        \u_outFIFO/FIFO[31][0] ), .S0(n35), .S1(n943), .Q(\u_outFIFO/n696 ) );
  IMUX40 \u_outFIFO/U692  ( .A(\u_outFIFO/FIFO[8][1] ), .B(
        \u_outFIFO/FIFO[9][1] ), .C(\u_outFIFO/FIFO[10][1] ), .D(
        \u_outFIFO/FIFO[11][1] ), .S0(n35), .S1(\u_outFIFO/N36 ), .Q(
        \u_outFIFO/n709 ) );
  IMUX40 \u_outFIFO/U694  ( .A(\u_outFIFO/FIFO[0][1] ), .B(
        \u_outFIFO/FIFO[1][1] ), .C(\u_outFIFO/FIFO[2][1] ), .D(
        \u_outFIFO/FIFO[3][1] ), .S0(n942), .S1(\u_outFIFO/N36 ), .Q(
        \u_outFIFO/n708 ) );
  IMUX40 \u_outFIFO/U691  ( .A(\u_outFIFO/FIFO[12][1] ), .B(
        \u_outFIFO/FIFO[13][1] ), .C(\u_outFIFO/FIFO[14][1] ), .D(
        \u_outFIFO/FIFO[15][1] ), .S0(n35), .S1(\u_outFIFO/N36 ), .Q(
        \u_outFIFO/n711 ) );
  IMUX40 \u_outFIFO/U700  ( .A(\u_outFIFO/FIFO[8][2] ), .B(
        \u_outFIFO/FIFO[9][2] ), .C(\u_outFIFO/FIFO[10][2] ), .D(
        \u_outFIFO/FIFO[11][2] ), .S0(n942), .S1(\u_outFIFO/N36 ), .Q(
        \u_outFIFO/n719 ) );
  IMUX40 \u_outFIFO/U702  ( .A(\u_outFIFO/FIFO[0][2] ), .B(
        \u_outFIFO/FIFO[1][2] ), .C(\u_outFIFO/FIFO[2][2] ), .D(
        \u_outFIFO/FIFO[3][2] ), .S0(n942), .S1(\u_outFIFO/N36 ), .Q(
        \u_outFIFO/n718 ) );
  IMUX40 \u_outFIFO/U699  ( .A(\u_outFIFO/FIFO[12][2] ), .B(
        \u_outFIFO/FIFO[13][2] ), .C(\u_outFIFO/FIFO[14][2] ), .D(
        \u_outFIFO/FIFO[15][2] ), .S0(n942), .S1(n943), .Q(\u_outFIFO/n721 )
         );
  IMUX40 \u_outFIFO/U708  ( .A(\u_outFIFO/FIFO[8][3] ), .B(
        \u_outFIFO/FIFO[9][3] ), .C(\u_outFIFO/FIFO[10][3] ), .D(
        \u_outFIFO/FIFO[11][3] ), .S0(n942), .S1(n943), .Q(\u_outFIFO/n729 )
         );
  IMUX40 \u_outFIFO/U710  ( .A(\u_outFIFO/FIFO[0][3] ), .B(
        \u_outFIFO/FIFO[1][3] ), .C(\u_outFIFO/FIFO[2][3] ), .D(
        \u_outFIFO/FIFO[3][3] ), .S0(n942), .S1(\u_outFIFO/N36 ), .Q(
        \u_outFIFO/n728 ) );
  IMUX40 \u_outFIFO/U707  ( .A(\u_outFIFO/FIFO[12][3] ), .B(
        \u_outFIFO/FIFO[13][3] ), .C(\u_outFIFO/FIFO[14][3] ), .D(
        \u_outFIFO/FIFO[15][3] ), .S0(n942), .S1(n943), .Q(\u_outFIFO/n731 )
         );
  IMUX40 \u_outFIFO/U682  ( .A(\u_outFIFO/FIFO[16][0] ), .B(
        \u_outFIFO/FIFO[17][0] ), .C(\u_outFIFO/FIFO[18][0] ), .D(
        \u_outFIFO/FIFO[19][0] ), .S0(n35), .S1(n943), .Q(\u_outFIFO/n693 ) );
  IMUX40 \u_outFIFO/U680  ( .A(\u_outFIFO/FIFO[24][0] ), .B(
        \u_outFIFO/FIFO[25][0] ), .C(\u_outFIFO/FIFO[26][0] ), .D(
        \u_outFIFO/FIFO[27][0] ), .S0(n35), .S1(n943), .Q(\u_outFIFO/n694 ) );
  IMUX40 \u_outFIFO/U681  ( .A(\u_outFIFO/FIFO[20][0] ), .B(
        \u_outFIFO/FIFO[21][0] ), .C(\u_outFIFO/FIFO[22][0] ), .D(
        \u_outFIFO/FIFO[23][0] ), .S0(n35), .S1(n943), .Q(\u_outFIFO/n695 ) );
  IMUX40 \u_outFIFO/U667  ( .A(\u_outFIFO/n693 ), .B(\u_outFIFO/n694 ), .C(
        \u_outFIFO/n695 ), .D(\u_outFIFO/n696 ), .S0(n775), .S1(n774), .Q(
        \u_outFIFO/n692 ) );
  IMUX21 \u_cordic/mycordic/U535  ( .A(\u_cordic/mycordic/n568 ), .B(n383), 
        .S(n782), .Q(\u_cordic/mycordic/n567 ) );
  MUX22 \u_cordic/mycordic/U536  ( .A(
        \u_cordic/mycordic/present_ANGLE_table[6][6] ), .B(
        \u_cordic/mycordic/n567 ), .S(n153), .Q(
        \u_cordic/mycordic/next_ANGLE_table[6][6] ) );
  IMUX21 \u_cordic/mycordic/U533  ( .A(\u_cordic/mycordic/n566 ), .B(n381), 
        .S(n783), .Q(\u_cordic/mycordic/n565 ) );
  MUX22 \u_cordic/mycordic/U534  ( .A(
        \u_cordic/mycordic/present_ANGLE_table[6][5] ), .B(
        \u_cordic/mycordic/n565 ), .S(n153), .Q(
        \u_cordic/mycordic/next_ANGLE_table[6][5] ) );
  IMUX21 \u_cordic/mycordic/U531  ( .A(\u_cordic/mycordic/n564 ), .B(n384), 
        .S(n781), .Q(\u_cordic/mycordic/n563 ) );
  MUX22 \u_cordic/mycordic/U532  ( .A(
        \u_cordic/mycordic/present_ANGLE_table[6][4] ), .B(
        \u_cordic/mycordic/n563 ), .S(n153), .Q(
        \u_cordic/mycordic/next_ANGLE_table[6][4] ) );
  IMUX21 \u_cordic/mycordic/U529  ( .A(\u_cordic/mycordic/n562 ), .B(n386), 
        .S(n782), .Q(\u_cordic/mycordic/n561 ) );
  MUX22 \u_cordic/mycordic/U530  ( .A(
        \u_cordic/mycordic/present_ANGLE_table[6][3] ), .B(
        \u_cordic/mycordic/n561 ), .S(n153), .Q(
        \u_cordic/mycordic/next_ANGLE_table[6][3] ) );
  IMUX21 \u_cordic/mycordic/U527  ( .A(\u_cordic/mycordic/n560 ), .B(
        \u_cordic/mycordic/present_ANGLE_table[6][2] ), .S(n783), .Q(
        \u_cordic/mycordic/n559 ) );
  MUX22 \u_cordic/mycordic/U528  ( .A(
        \u_cordic/mycordic/present_ANGLE_table[6][2] ), .B(
        \u_cordic/mycordic/n559 ), .S(n153), .Q(
        \u_cordic/mycordic/next_ANGLE_table[6][2] ) );
  IMUX21 \u_cordic/mycordic/U525  ( .A(\u_cordic/mycordic/n558 ), .B(n311), 
        .S(n781), .Q(\u_cordic/mycordic/n557 ) );
  MUX22 \u_cordic/mycordic/U526  ( .A(
        \u_cordic/mycordic/present_ANGLE_table[6][1] ), .B(
        \u_cordic/mycordic/n557 ), .S(n153), .Q(
        \u_cordic/mycordic/next_ANGLE_table[6][1] ) );
  IMUX21 \u_cordic/mycordic/U523  ( .A(\u_cordic/mycordic/n556 ), .B(n310), 
        .S(n782), .Q(\u_cordic/mycordic/n555 ) );
  MUX22 \u_cordic/mycordic/U524  ( .A(\u_cordic/mycordic/N615 ), .B(
        \u_cordic/mycordic/n555 ), .S(n153), .Q(
        \u_cordic/mycordic/next_ANGLE_table[6][0] ) );
  IMUX40 \u_inFIFO/U258  ( .A(\u_inFIFO/FIFO[4][1] ), .B(\u_inFIFO/FIFO[5][1] ), .C(\u_inFIFO/FIFO[6][1] ), .D(\u_inFIFO/FIFO[7][1] ), .S0(n34), .S1(
        \u_inFIFO/N34 ), .Q(\u_inFIFO/n273 ) );
  IMUX40 \u_inFIFO/U235  ( .A(\u_inFIFO/n266 ), .B(\u_inFIFO/n267 ), .C(
        \u_inFIFO/n268 ), .D(\u_inFIFO/n269 ), .S0(n780), .S1(n779), .Q(
        \u_inFIFO/n265 ) );
  IMUX40 \u_inFIFO/U236  ( .A(\u_inFIFO/n271 ), .B(\u_inFIFO/n272 ), .C(
        \u_inFIFO/n273 ), .D(\u_inFIFO/n274 ), .S0(n780), .S1(n779), .Q(
        \u_inFIFO/n270 ) );
  MUX22 \u_inFIFO/U237  ( .A(\u_inFIFO/n270 ), .B(\u_inFIFO/n265 ), .S(
        \u_inFIFO/N37 ), .Q(\u_inFIFO/N182 ) );
  IMUX40 \u_inFIFO/U274  ( .A(\u_inFIFO/FIFO[4][3] ), .B(\u_inFIFO/FIFO[5][3] ), .C(\u_inFIFO/FIFO[6][3] ), .D(\u_inFIFO/FIFO[7][3] ), .S0(n964), .S1(n965), 
        .Q(\u_inFIFO/n293 ) );
  IMUX40 \u_inFIFO/U241  ( .A(\u_inFIFO/n286 ), .B(\u_inFIFO/n287 ), .C(
        \u_inFIFO/n288 ), .D(\u_inFIFO/n289 ), .S0(n780), .S1(n779), .Q(
        \u_inFIFO/n285 ) );
  IMUX40 \u_inFIFO/U242  ( .A(\u_inFIFO/n291 ), .B(\u_inFIFO/n292 ), .C(
        \u_inFIFO/n293 ), .D(\u_inFIFO/n294 ), .S0(n780), .S1(n779), .Q(
        \u_inFIFO/n290 ) );
  MUX22 \u_inFIFO/U243  ( .A(\u_inFIFO/n290 ), .B(\u_inFIFO/n285 ), .S(
        \u_inFIFO/N37 ), .Q(\u_inFIFO/N180 ) );
  IMUX40 \u_inFIFO/U266  ( .A(\u_inFIFO/FIFO[4][2] ), .B(\u_inFIFO/FIFO[5][2] ), .C(\u_inFIFO/FIFO[6][2] ), .D(\u_inFIFO/FIFO[7][2] ), .S0(n964), .S1(n965), 
        .Q(\u_inFIFO/n283 ) );
  IMUX40 \u_inFIFO/U238  ( .A(\u_inFIFO/n276 ), .B(\u_inFIFO/n277 ), .C(
        \u_inFIFO/n278 ), .D(\u_inFIFO/n279 ), .S0(n780), .S1(n779), .Q(
        \u_inFIFO/n275 ) );
  IMUX40 \u_inFIFO/U239  ( .A(\u_inFIFO/n281 ), .B(\u_inFIFO/n282 ), .C(
        \u_inFIFO/n283 ), .D(\u_inFIFO/n284 ), .S0(n780), .S1(n779), .Q(
        \u_inFIFO/n280 ) );
  MUX22 \u_inFIFO/U240  ( .A(\u_inFIFO/n280 ), .B(\u_inFIFO/n275 ), .S(
        \u_inFIFO/N37 ), .Q(\u_inFIFO/N181 ) );
  MUX22 \u_inFIFO/U234  ( .A(\u_inFIFO/n260 ), .B(\u_inFIFO/n255 ), .S(
        \u_inFIFO/N37 ), .Q(\u_inFIFO/N183 ) );
  IMUX40 \u_outFIFO/U668  ( .A(\u_outFIFO/n698 ), .B(\u_outFIFO/n699 ), .C(
        \u_outFIFO/n700 ), .D(\u_outFIFO/n701 ), .S0(n775), .S1(n774), .Q(
        \u_outFIFO/n697 ) );
  MUX22 \u_outFIFO/U669  ( .A(\u_outFIFO/n697 ), .B(\u_outFIFO/n692 ), .S(
        \u_outFIFO/N39 ), .Q(\u_outFIFO/N185 ) );
  IMUX40 \u_outFIFO/U671  ( .A(\u_outFIFO/n708 ), .B(\u_outFIFO/n709 ), .C(
        \u_outFIFO/n710 ), .D(\u_outFIFO/n711 ), .S0(n775), .S1(n774), .Q(
        \u_outFIFO/n707 ) );
  MUX22 \u_outFIFO/U672  ( .A(\u_outFIFO/n707 ), .B(\u_outFIFO/n702 ), .S(
        \u_outFIFO/N39 ), .Q(\u_outFIFO/N184 ) );
  IMUX40 \u_outFIFO/U674  ( .A(\u_outFIFO/n718 ), .B(\u_outFIFO/n719 ), .C(
        \u_outFIFO/n720 ), .D(\u_outFIFO/n721 ), .S0(n775), .S1(n774), .Q(
        \u_outFIFO/n717 ) );
  MUX22 \u_outFIFO/U675  ( .A(\u_outFIFO/n717 ), .B(\u_outFIFO/n712 ), .S(
        \u_outFIFO/N39 ), .Q(\u_outFIFO/N183 ) );
  IMUX40 \u_outFIFO/U677  ( .A(\u_outFIFO/n728 ), .B(\u_outFIFO/n729 ), .C(
        \u_outFIFO/n730 ), .D(\u_outFIFO/n731 ), .S0(n775), .S1(n774), .Q(
        \u_outFIFO/n727 ) );
  MUX22 \u_outFIFO/U678  ( .A(\u_outFIFO/n727 ), .B(\u_outFIFO/n722 ), .S(
        \u_outFIFO/N39 ), .Q(\u_outFIFO/N182 ) );
  NAND22 \u_cordic/mycordic/U564  ( .A(\u_cordic/mycordic/N622 ), .B(n751), 
        .Q(\u_cordic/mycordic/n570 ) );
  NAND22 \u_cordic/mycordic/U563  ( .A(\u_cordic/mycordic/N621 ), .B(n751), 
        .Q(\u_cordic/mycordic/n568 ) );
  IMUX40 \u_inFIFO/U270  ( .A(\u_inFIFO/FIFO[20][3] ), .B(
        \u_inFIFO/FIFO[21][3] ), .C(\u_inFIFO/FIFO[22][3] ), .D(
        \u_inFIFO/FIFO[23][3] ), .S0(n964), .S1(n965), .Q(\u_inFIFO/n288 ) );
  IMUX40 \u_inFIFO/U262  ( .A(\u_inFIFO/FIFO[20][2] ), .B(
        \u_inFIFO/FIFO[21][2] ), .C(\u_inFIFO/FIFO[22][2] ), .D(
        \u_inFIFO/FIFO[23][2] ), .S0(n34), .S1(\u_inFIFO/N34 ), .Q(
        \u_inFIFO/n278 ) );
  IMUX40 \u_inFIFO/U254  ( .A(\u_inFIFO/FIFO[20][1] ), .B(
        \u_inFIFO/FIFO[21][1] ), .C(\u_inFIFO/FIFO[22][1] ), .D(
        \u_inFIFO/FIFO[23][1] ), .S0(n964), .S1(\u_inFIFO/N34 ), .Q(
        \u_inFIFO/n268 ) );
  IMUX40 \u_inFIFO/U248  ( .A(\u_inFIFO/FIFO[12][0] ), .B(
        \u_inFIFO/FIFO[13][0] ), .C(\u_inFIFO/FIFO[14][0] ), .D(
        \u_inFIFO/FIFO[15][0] ), .S0(n34), .S1(\u_inFIFO/N34 ), .Q(
        \u_inFIFO/n264 ) );
  IMUX40 \u_inFIFO/U244  ( .A(\u_inFIFO/FIFO[28][0] ), .B(
        \u_inFIFO/FIFO[29][0] ), .C(\u_inFIFO/FIFO[30][0] ), .D(
        \u_inFIFO/FIFO[31][0] ), .S0(n34), .S1(n965), .Q(\u_inFIFO/n259 ) );
  IMUX40 \u_inFIFO/U273  ( .A(\u_inFIFO/FIFO[8][3] ), .B(\u_inFIFO/FIFO[9][3] ), .C(\u_inFIFO/FIFO[10][3] ), .D(\u_inFIFO/FIFO[11][3] ), .S0(n964), .S1(n965), 
        .Q(\u_inFIFO/n292 ) );
  IMUX40 \u_inFIFO/U275  ( .A(\u_inFIFO/FIFO[0][3] ), .B(\u_inFIFO/FIFO[1][3] ), .C(\u_inFIFO/FIFO[2][3] ), .D(\u_inFIFO/FIFO[3][3] ), .S0(n964), .S1(
        \u_inFIFO/N34 ), .Q(\u_inFIFO/n291 ) );
  IMUX40 \u_inFIFO/U272  ( .A(\u_inFIFO/FIFO[12][3] ), .B(
        \u_inFIFO/FIFO[13][3] ), .C(\u_inFIFO/FIFO[14][3] ), .D(
        \u_inFIFO/FIFO[15][3] ), .S0(n964), .S1(n965), .Q(\u_inFIFO/n294 ) );
  IMUX40 \u_inFIFO/U269  ( .A(\u_inFIFO/FIFO[24][3] ), .B(
        \u_inFIFO/FIFO[25][3] ), .C(\u_inFIFO/FIFO[26][3] ), .D(
        \u_inFIFO/FIFO[27][3] ), .S0(n964), .S1(n965), .Q(\u_inFIFO/n287 ) );
  IMUX40 \u_inFIFO/U271  ( .A(\u_inFIFO/FIFO[16][3] ), .B(
        \u_inFIFO/FIFO[17][3] ), .C(\u_inFIFO/FIFO[18][3] ), .D(
        \u_inFIFO/FIFO[19][3] ), .S0(n964), .S1(n965), .Q(\u_inFIFO/n286 ) );
  IMUX40 \u_inFIFO/U268  ( .A(\u_inFIFO/FIFO[28][3] ), .B(
        \u_inFIFO/FIFO[29][3] ), .C(\u_inFIFO/FIFO[30][3] ), .D(
        \u_inFIFO/FIFO[31][3] ), .S0(n964), .S1(n965), .Q(\u_inFIFO/n289 ) );
  IMUX40 \u_inFIFO/U265  ( .A(\u_inFIFO/FIFO[8][2] ), .B(\u_inFIFO/FIFO[9][2] ), .C(\u_inFIFO/FIFO[10][2] ), .D(\u_inFIFO/FIFO[11][2] ), .S0(n964), .S1(n965), 
        .Q(\u_inFIFO/n282 ) );
  IMUX40 \u_inFIFO/U267  ( .A(\u_inFIFO/FIFO[0][2] ), .B(\u_inFIFO/FIFO[1][2] ), .C(\u_inFIFO/FIFO[2][2] ), .D(\u_inFIFO/FIFO[3][2] ), .S0(n964), .S1(n965), 
        .Q(\u_inFIFO/n281 ) );
  IMUX40 \u_inFIFO/U264  ( .A(\u_inFIFO/FIFO[12][2] ), .B(
        \u_inFIFO/FIFO[13][2] ), .C(\u_inFIFO/FIFO[14][2] ), .D(
        \u_inFIFO/FIFO[15][2] ), .S0(n964), .S1(n965), .Q(\u_inFIFO/n284 ) );
  IMUX40 \u_inFIFO/U261  ( .A(\u_inFIFO/FIFO[24][2] ), .B(
        \u_inFIFO/FIFO[25][2] ), .C(\u_inFIFO/FIFO[26][2] ), .D(
        \u_inFIFO/FIFO[27][2] ), .S0(n34), .S1(\u_inFIFO/N34 ), .Q(
        \u_inFIFO/n277 ) );
  IMUX40 \u_inFIFO/U263  ( .A(\u_inFIFO/FIFO[16][2] ), .B(
        \u_inFIFO/FIFO[17][2] ), .C(\u_inFIFO/FIFO[18][2] ), .D(
        \u_inFIFO/FIFO[19][2] ), .S0(n964), .S1(\u_inFIFO/N34 ), .Q(
        \u_inFIFO/n276 ) );
  IMUX40 \u_inFIFO/U260  ( .A(\u_inFIFO/FIFO[28][2] ), .B(
        \u_inFIFO/FIFO[29][2] ), .C(\u_inFIFO/FIFO[30][2] ), .D(
        \u_inFIFO/FIFO[31][2] ), .S0(n34), .S1(\u_inFIFO/N34 ), .Q(
        \u_inFIFO/n279 ) );
  IMUX40 \u_inFIFO/U257  ( .A(\u_inFIFO/FIFO[8][1] ), .B(\u_inFIFO/FIFO[9][1] ), .C(\u_inFIFO/FIFO[10][1] ), .D(\u_inFIFO/FIFO[11][1] ), .S0(n34), .S1(
        \u_inFIFO/N34 ), .Q(\u_inFIFO/n272 ) );
  IMUX40 \u_inFIFO/U259  ( .A(\u_inFIFO/FIFO[0][1] ), .B(\u_inFIFO/FIFO[1][1] ), .C(\u_inFIFO/FIFO[2][1] ), .D(\u_inFIFO/FIFO[3][1] ), .S0(n964), .S1(
        \u_inFIFO/N34 ), .Q(\u_inFIFO/n271 ) );
  IMUX40 \u_inFIFO/U256  ( .A(\u_inFIFO/FIFO[12][1] ), .B(
        \u_inFIFO/FIFO[13][1] ), .C(\u_inFIFO/FIFO[14][1] ), .D(
        \u_inFIFO/FIFO[15][1] ), .S0(n34), .S1(\u_inFIFO/N34 ), .Q(
        \u_inFIFO/n274 ) );
  IMUX40 \u_inFIFO/U253  ( .A(\u_inFIFO/FIFO[24][1] ), .B(
        \u_inFIFO/FIFO[25][1] ), .C(\u_inFIFO/FIFO[26][1] ), .D(
        \u_inFIFO/FIFO[27][1] ), .S0(n34), .S1(\u_inFIFO/N34 ), .Q(
        \u_inFIFO/n267 ) );
  IMUX40 \u_inFIFO/U255  ( .A(\u_inFIFO/FIFO[16][1] ), .B(
        \u_inFIFO/FIFO[17][1] ), .C(\u_inFIFO/FIFO[18][1] ), .D(
        \u_inFIFO/FIFO[19][1] ), .S0(n964), .S1(\u_inFIFO/N34 ), .Q(
        \u_inFIFO/n266 ) );
  IMUX40 \u_inFIFO/U252  ( .A(\u_inFIFO/FIFO[28][1] ), .B(
        \u_inFIFO/FIFO[29][1] ), .C(\u_inFIFO/FIFO[30][1] ), .D(
        \u_inFIFO/FIFO[31][1] ), .S0(n34), .S1(\u_inFIFO/N34 ), .Q(
        \u_inFIFO/n269 ) );
  IMUX40 \u_outFIFO/U687  ( .A(\u_outFIFO/FIFO[28][1] ), .B(
        \u_outFIFO/FIFO[29][1] ), .C(\u_outFIFO/FIFO[30][1] ), .D(
        \u_outFIFO/FIFO[31][1] ), .S0(n35), .S1(\u_outFIFO/N36 ), .Q(
        \u_outFIFO/n706 ) );
  IMUX40 \u_outFIFO/U695  ( .A(\u_outFIFO/FIFO[28][2] ), .B(
        \u_outFIFO/FIFO[29][2] ), .C(\u_outFIFO/FIFO[30][2] ), .D(
        \u_outFIFO/FIFO[31][2] ), .S0(n35), .S1(\u_outFIFO/N36 ), .Q(
        \u_outFIFO/n716 ) );
  IMUX40 \u_outFIFO/U703  ( .A(\u_outFIFO/FIFO[28][3] ), .B(
        \u_outFIFO/FIFO[29][3] ), .C(\u_outFIFO/FIFO[30][3] ), .D(
        \u_outFIFO/FIFO[31][3] ), .S0(n942), .S1(n943), .Q(\u_outFIFO/n726 )
         );
  IMUX40 \u_outFIFO/U690  ( .A(\u_outFIFO/FIFO[16][1] ), .B(
        \u_outFIFO/FIFO[17][1] ), .C(\u_outFIFO/FIFO[18][1] ), .D(
        \u_outFIFO/FIFO[19][1] ), .S0(n942), .S1(\u_outFIFO/N36 ), .Q(
        \u_outFIFO/n703 ) );
  IMUX40 \u_outFIFO/U688  ( .A(\u_outFIFO/FIFO[24][1] ), .B(
        \u_outFIFO/FIFO[25][1] ), .C(\u_outFIFO/FIFO[26][1] ), .D(
        \u_outFIFO/FIFO[27][1] ), .S0(n35), .S1(\u_outFIFO/N36 ), .Q(
        \u_outFIFO/n704 ) );
  IMUX40 \u_outFIFO/U689  ( .A(\u_outFIFO/FIFO[20][1] ), .B(
        \u_outFIFO/FIFO[21][1] ), .C(\u_outFIFO/FIFO[22][1] ), .D(
        \u_outFIFO/FIFO[23][1] ), .S0(n942), .S1(\u_outFIFO/N36 ), .Q(
        \u_outFIFO/n705 ) );
  IMUX40 \u_outFIFO/U670  ( .A(\u_outFIFO/n703 ), .B(\u_outFIFO/n704 ), .C(
        \u_outFIFO/n705 ), .D(\u_outFIFO/n706 ), .S0(n775), .S1(n774), .Q(
        \u_outFIFO/n702 ) );
  IMUX40 \u_outFIFO/U698  ( .A(\u_outFIFO/FIFO[16][2] ), .B(
        \u_outFIFO/FIFO[17][2] ), .C(\u_outFIFO/FIFO[18][2] ), .D(
        \u_outFIFO/FIFO[19][2] ), .S0(n942), .S1(\u_outFIFO/N36 ), .Q(
        \u_outFIFO/n713 ) );
  IMUX40 \u_outFIFO/U696  ( .A(\u_outFIFO/FIFO[24][2] ), .B(
        \u_outFIFO/FIFO[25][2] ), .C(\u_outFIFO/FIFO[26][2] ), .D(
        \u_outFIFO/FIFO[27][2] ), .S0(n35), .S1(\u_outFIFO/N36 ), .Q(
        \u_outFIFO/n714 ) );
  IMUX40 \u_outFIFO/U697  ( .A(\u_outFIFO/FIFO[20][2] ), .B(
        \u_outFIFO/FIFO[21][2] ), .C(\u_outFIFO/FIFO[22][2] ), .D(
        \u_outFIFO/FIFO[23][2] ), .S0(n35), .S1(\u_outFIFO/N36 ), .Q(
        \u_outFIFO/n715 ) );
  IMUX40 \u_outFIFO/U673  ( .A(\u_outFIFO/n713 ), .B(\u_outFIFO/n714 ), .C(
        \u_outFIFO/n715 ), .D(\u_outFIFO/n716 ), .S0(n775), .S1(n774), .Q(
        \u_outFIFO/n712 ) );
  IMUX40 \u_outFIFO/U706  ( .A(\u_outFIFO/FIFO[16][3] ), .B(
        \u_outFIFO/FIFO[17][3] ), .C(\u_outFIFO/FIFO[18][3] ), .D(
        \u_outFIFO/FIFO[19][3] ), .S0(n942), .S1(\u_outFIFO/N36 ), .Q(
        \u_outFIFO/n723 ) );
  IMUX40 \u_outFIFO/U704  ( .A(\u_outFIFO/FIFO[24][3] ), .B(
        \u_outFIFO/FIFO[25][3] ), .C(\u_outFIFO/FIFO[26][3] ), .D(
        \u_outFIFO/FIFO[27][3] ), .S0(n942), .S1(\u_outFIFO/N36 ), .Q(
        \u_outFIFO/n724 ) );
  IMUX40 \u_outFIFO/U705  ( .A(\u_outFIFO/FIFO[20][3] ), .B(
        \u_outFIFO/FIFO[21][3] ), .C(\u_outFIFO/FIFO[22][3] ), .D(
        \u_outFIFO/FIFO[23][3] ), .S0(n942), .S1(\u_outFIFO/N36 ), .Q(
        \u_outFIFO/n725 ) );
  IMUX40 \u_outFIFO/U676  ( .A(\u_outFIFO/n723 ), .B(\u_outFIFO/n724 ), .C(
        \u_outFIFO/n725 ), .D(\u_outFIFO/n726 ), .S0(n775), .S1(n774), .Q(
        \u_outFIFO/n722 ) );
  IMUX40 \u_inFIFO/U247  ( .A(\u_inFIFO/FIFO[16][0] ), .B(
        \u_inFIFO/FIFO[17][0] ), .C(\u_inFIFO/FIFO[18][0] ), .D(
        \u_inFIFO/FIFO[19][0] ), .S0(n34), .S1(n965), .Q(\u_inFIFO/n256 ) );
  IMUX40 \u_inFIFO/U245  ( .A(\u_inFIFO/FIFO[24][0] ), .B(
        \u_inFIFO/FIFO[25][0] ), .C(\u_inFIFO/FIFO[26][0] ), .D(
        \u_inFIFO/FIFO[27][0] ), .S0(n34), .S1(n965), .Q(\u_inFIFO/n257 ) );
  IMUX40 \u_inFIFO/U246  ( .A(\u_inFIFO/FIFO[20][0] ), .B(
        \u_inFIFO/FIFO[21][0] ), .C(\u_inFIFO/FIFO[22][0] ), .D(
        \u_inFIFO/FIFO[23][0] ), .S0(n34), .S1(n965), .Q(\u_inFIFO/n258 ) );
  IMUX40 \u_inFIFO/U232  ( .A(\u_inFIFO/n256 ), .B(\u_inFIFO/n257 ), .C(
        \u_inFIFO/n258 ), .D(\u_inFIFO/n259 ), .S0(n780), .S1(n779), .Q(
        \u_inFIFO/n255 ) );
  IMUX40 \u_inFIFO/U251  ( .A(\u_inFIFO/FIFO[0][0] ), .B(\u_inFIFO/FIFO[1][0] ), .C(\u_inFIFO/FIFO[2][0] ), .D(\u_inFIFO/FIFO[3][0] ), .S0(n34), .S1(
        \u_inFIFO/N34 ), .Q(\u_inFIFO/n261 ) );
  IMUX40 \u_inFIFO/U249  ( .A(\u_inFIFO/FIFO[8][0] ), .B(\u_inFIFO/FIFO[9][0] ), .C(\u_inFIFO/FIFO[10][0] ), .D(\u_inFIFO/FIFO[11][0] ), .S0(n34), .S1(
        \u_inFIFO/N34 ), .Q(\u_inFIFO/n262 ) );
  IMUX40 \u_inFIFO/U250  ( .A(\u_inFIFO/FIFO[4][0] ), .B(\u_inFIFO/FIFO[5][0] ), .C(\u_inFIFO/FIFO[6][0] ), .D(\u_inFIFO/FIFO[7][0] ), .S0(n34), .S1(
        \u_inFIFO/N34 ), .Q(\u_inFIFO/n263 ) );
  IMUX40 \u_inFIFO/U233  ( .A(\u_inFIFO/n261 ), .B(\u_inFIFO/n262 ), .C(
        \u_inFIFO/n263 ), .D(\u_inFIFO/n264 ), .S0(n780), .S1(n779), .Q(
        \u_inFIFO/n260 ) );
  IMUX21 \u_cordic/mycordic/U541  ( .A(\u_cordic/mycordic/n574 ), .B(n378), 
        .S(n782), .Q(\u_cordic/mycordic/n573 ) );
  MUX22 \u_cordic/mycordic/U542  ( .A(
        \u_cordic/mycordic/present_ANGLE_table[6][9] ), .B(
        \u_cordic/mycordic/n573 ), .S(n153), .Q(
        \u_cordic/mycordic/next_ANGLE_table[6][9] ) );
  IMUX21 \u_cordic/mycordic/U537  ( .A(\u_cordic/mycordic/n570 ), .B(n376), 
        .S(n781), .Q(\u_cordic/mycordic/n569 ) );
  MUX22 \u_cordic/mycordic/U538  ( .A(
        \u_cordic/mycordic/present_ANGLE_table[6][7] ), .B(
        \u_cordic/mycordic/n569 ), .S(n153), .Q(
        \u_cordic/mycordic/next_ANGLE_table[6][7] ) );
  XOR31 \u_cordic/mycordic/sub_182/U2_7  ( .A(
        \u_cordic/mycordic/present_I_table[1][7] ), .B(n277), .C(
        \u_cordic/mycordic/sub_182/carry [7]), .Q(\u_cordic/mycordic/N291 ) );
  XOR31 \u_cordic/mycordic/sub_178/U2_7  ( .A(
        \u_cordic/mycordic/present_Q_table[1][7] ), .B(n280), .C(
        \u_cordic/mycordic/sub_178/carry [7]), .Q(\u_cordic/mycordic/N267 ) );
  NAND22 \u_cordic/mycordic/U565  ( .A(\u_cordic/mycordic/N623 ), .B(n750), 
        .Q(\u_cordic/mycordic/n572 ) );
  IMUX21 \u_cordic/mycordic/U539  ( .A(\u_cordic/mycordic/n572 ), .B(n379), 
        .S(n783), .Q(\u_cordic/mycordic/n571 ) );
  MUX22 \u_cordic/mycordic/U540  ( .A(
        \u_cordic/mycordic/present_ANGLE_table[6][8] ), .B(
        \u_cordic/mycordic/n571 ), .S(n153), .Q(
        \u_cordic/mycordic/next_ANGLE_table[6][8] ) );
  NAND22 \u_cordic/mycordic/U566  ( .A(\u_cordic/mycordic/N624 ), .B(n750), 
        .Q(\u_cordic/mycordic/n574 ) );
  NAND22 \u_cordic/mycordic/U567  ( .A(\u_cordic/mycordic/N625 ), .B(n750), 
        .Q(\u_cordic/mycordic/n576 ) );
  IMUX21 \u_cordic/mycordic/U545  ( .A(\u_cordic/mycordic/n578 ), .B(n374), 
        .S(n783), .Q(\u_cordic/mycordic/n577 ) );
  MUX22 \u_cordic/mycordic/U546  ( .A(
        \u_cordic/mycordic/present_ANGLE_table[6][11] ), .B(
        \u_cordic/mycordic/n577 ), .S(n153), .Q(
        \u_cordic/mycordic/next_ANGLE_table[6][11] ) );
  IMUX21 \u_cordic/mycordic/U543  ( .A(\u_cordic/mycordic/n576 ), .B(n373), 
        .S(n781), .Q(\u_cordic/mycordic/n575 ) );
  MUX22 \u_cordic/mycordic/U544  ( .A(
        \u_cordic/mycordic/present_ANGLE_table[6][10] ), .B(
        \u_cordic/mycordic/n575 ), .S(n153), .Q(
        \u_cordic/mycordic/next_ANGLE_table[6][10] ) );
  NAND22 \u_cordic/mycordic/U569  ( .A(\u_cordic/mycordic/N627 ), .B(n750), 
        .Q(\u_cordic/mycordic/n580 ) );
  NAND22 \u_cordic/mycordic/U568  ( .A(\u_cordic/mycordic/N626 ), .B(n750), 
        .Q(\u_cordic/mycordic/n578 ) );
  IMUX21 \u_cordic/mycordic/U551  ( .A(\u_cordic/mycordic/n584 ), .B(n372), 
        .S(n783), .Q(\u_cordic/mycordic/n583 ) );
  MUX22 \u_cordic/mycordic/U552  ( .A(
        \u_cordic/mycordic/present_ANGLE_table[6][14] ), .B(
        \u_cordic/mycordic/n583 ), .S(n153), .Q(
        \u_cordic/mycordic/next_ANGLE_table[6][14] ) );
  IMUX21 \u_cordic/mycordic/U549  ( .A(\u_cordic/mycordic/n582 ), .B(n371), 
        .S(n781), .Q(\u_cordic/mycordic/n581 ) );
  MUX22 \u_cordic/mycordic/U550  ( .A(
        \u_cordic/mycordic/present_ANGLE_table[6][13] ), .B(
        \u_cordic/mycordic/n581 ), .S(n153), .Q(
        \u_cordic/mycordic/next_ANGLE_table[6][13] ) );
  IMUX21 \u_cordic/mycordic/U547  ( .A(\u_cordic/mycordic/n580 ), .B(n370), 
        .S(n782), .Q(\u_cordic/mycordic/n579 ) );
  MUX22 \u_cordic/mycordic/U548  ( .A(
        \u_cordic/mycordic/present_ANGLE_table[6][12] ), .B(
        \u_cordic/mycordic/n579 ), .S(n153), .Q(
        \u_cordic/mycordic/next_ANGLE_table[6][12] ) );
  XOR31 \u_cordic/mycordic/sub_223/U2_7  ( .A(
        \u_cordic/mycordic/present_Q_table[5][7] ), .B(n182), .C(
        \u_cordic/mycordic/sub_223/carry[7] ), .Q(\u_cordic/mycordic/N500 ) );
  XOR31 \u_cordic/mycordic/add_228/U1_7  ( .A(
        \u_cordic/mycordic/present_Q_table[5][7] ), .B(
        \u_cordic/mycordic/present_I_table[5][7] ), .C(
        \u_cordic/mycordic/add_228/carry[7] ), .Q(\u_cordic/mycordic/N517 ) );
  XOR31 \u_cordic/mycordic/sub_212/U2_7  ( .A(n749), .B(n214), .C(
        \u_cordic/mycordic/sub_212/carry [7]), .Q(\u_cordic/mycordic/N455 ) );
  XOR31 \u_cordic/mycordic/add_217/U1_7  ( .A(n749), .B(
        \u_cordic/mycordic/present_I_table[4][7] ), .C(
        \u_cordic/mycordic/add_217/carry [7]), .Q(\u_cordic/mycordic/N483 ) );
  XOR31 \u_cordic/mycordic/add_211/U1_7  ( .A(
        \u_cordic/mycordic/present_I_table[4][7] ), .B(n749), .C(
        \u_cordic/mycordic/add_211/carry [7]), .Q(\u_cordic/mycordic/N447 ) );
  XOR31 \u_cordic/mycordic/sub_216/U2_7  ( .A(
        \u_cordic/mycordic/present_I_table[4][7] ), .B(n180), .C(
        \u_cordic/mycordic/sub_216/carry [7]), .Q(\u_cordic/mycordic/N475 ) );
  XOR31 \u_cordic/mycordic/sub_190/U2_7  ( .A(
        \u_cordic/mycordic/present_Q_table[2][7] ), .B(n270), .C(
        \u_cordic/mycordic/sub_190/carry [7]), .Q(\u_cordic/mycordic/N331 ) );
  XOR31 \u_cordic/mycordic/add_195/U1_7  ( .A(
        \u_cordic/mycordic/present_Q_table[2][7] ), .B(
        \u_cordic/mycordic/present_I_table[2][7] ), .C(
        \u_cordic/mycordic/add_195/carry [7]), .Q(\u_cordic/mycordic/N363 ) );
  XOR31 \u_cordic/mycordic/sub_194/U2_7  ( .A(
        \u_cordic/mycordic/present_I_table[2][7] ), .B(n268), .C(
        \u_cordic/mycordic/sub_194/carry [7]), .Q(\u_cordic/mycordic/N355 ) );
  XOR31 \u_cordic/mycordic/add_189/U1_7  ( .A(
        \u_cordic/mycordic/present_I_table[2][7] ), .B(
        \u_cordic/mycordic/present_Q_table[2][7] ), .C(
        \u_cordic/mycordic/add_189/carry [7]), .Q(\u_cordic/mycordic/N323 ) );
  XOR31 \u_cordic/mycordic/sub_201/U2_7  ( .A(
        \u_cordic/mycordic/present_Q_table[3][7] ), .B(n243), .C(
        \u_cordic/mycordic/sub_201/carry [7]), .Q(\u_cordic/mycordic/N395 ) );
  XOR31 \u_cordic/mycordic/add_206/U1_7  ( .A(
        \u_cordic/mycordic/present_Q_table[3][7] ), .B(
        \u_cordic/mycordic/present_I_table[3][7] ), .C(
        \u_cordic/mycordic/add_206/carry [7]), .Q(\u_cordic/mycordic/N427 ) );
  XOR31 \u_cordic/mycordic/sub_205/U2_7  ( .A(
        \u_cordic/mycordic/present_I_table[3][7] ), .B(n242), .C(
        \u_cordic/mycordic/sub_205/carry [7]), .Q(\u_cordic/mycordic/N419 ) );
  XOR31 \u_cordic/mycordic/add_200/U1_7  ( .A(
        \u_cordic/mycordic/present_I_table[3][7] ), .B(
        \u_cordic/mycordic/present_Q_table[3][7] ), .C(
        \u_cordic/mycordic/add_200/carry [7]), .Q(\u_cordic/mycordic/N387 ) );
  NAND22 \u_cordic/mycordic/U571  ( .A(\u_cordic/mycordic/N629 ), .B(n750), 
        .Q(\u_cordic/mycordic/n584 ) );
  NAND22 \u_cordic/mycordic/U570  ( .A(\u_cordic/mycordic/N628 ), .B(n750), 
        .Q(\u_cordic/mycordic/n582 ) );
  NAND22 \u_cordic/mycordic/U572  ( .A(\u_cordic/mycordic/N630 ), .B(n750), 
        .Q(\u_cordic/mycordic/n586 ) );
  IMUX21 \u_cordic/mycordic/U553  ( .A(\u_cordic/mycordic/n586 ), .B(n76), .S(
        n782), .Q(\u_cordic/mycordic/n585 ) );
  MUX22 \u_cordic/mycordic/U554  ( .A(
        \u_cordic/mycordic/present_ANGLE_table[6][15] ), .B(
        \u_cordic/mycordic/n585 ), .S(n153), .Q(
        \u_cordic/mycordic/next_ANGLE_table[6][15] ) );
  XOR31 \u_decoder/fir_filter/add_294/U1_14  ( .A(
        \u_decoder/fir_filter/I_data_mult_0_buff [14]), .B(
        \u_decoder/fir_filter/I_data_add_1_buff [14]), .C(
        \u_decoder/fir_filter/add_294/carry [14]), .Q(
        \u_decoder/fir_filter/I_data_add_0 [14]) );
  XOR31 \u_decoder/fir_filter/add_295/U1_14  ( .A(
        \u_decoder/fir_filter/I_data_mult_1_buff [14]), .B(
        \u_decoder/fir_filter/I_data_add_2_buff [14]), .C(
        \u_decoder/fir_filter/add_295/carry [14]), .Q(
        \u_decoder/fir_filter/I_data_add_1 [14]) );
  XOR31 \u_decoder/fir_filter/add_296/U1_14  ( .A(
        \u_decoder/fir_filter/I_data_mult_2_buff [14]), .B(
        \u_decoder/fir_filter/I_data_add_3_buff [14]), .C(
        \u_decoder/fir_filter/add_296/carry [14]), .Q(
        \u_decoder/fir_filter/I_data_add_2 [14]) );
  XOR31 \u_decoder/fir_filter/add_297/U1_14  ( .A(
        \u_decoder/fir_filter/I_data_mult_3_buff [14]), .B(
        \u_decoder/fir_filter/I_data_add_4_buff [14]), .C(
        \u_decoder/fir_filter/add_297/carry [14]), .Q(
        \u_decoder/fir_filter/I_data_add_3 [14]) );
  XOR31 \u_decoder/fir_filter/add_326/U1_14  ( .A(
        \u_decoder/fir_filter/Q_data_mult_0_buff [14]), .B(
        \u_decoder/fir_filter/Q_data_add_1_buff [14]), .C(
        \u_decoder/fir_filter/add_326/carry [14]), .Q(
        \u_decoder/fir_filter/Q_data_add_0 [14]) );
  XOR31 \u_decoder/fir_filter/add_327/U1_14  ( .A(
        \u_decoder/fir_filter/Q_data_mult_1_buff [14]), .B(
        \u_decoder/fir_filter/Q_data_add_2_buff [14]), .C(
        \u_decoder/fir_filter/add_327/carry [14]), .Q(
        \u_decoder/fir_filter/Q_data_add_1 [14]) );
  XOR31 \u_decoder/fir_filter/add_328/U1_14  ( .A(
        \u_decoder/fir_filter/Q_data_mult_2_buff [14]), .B(
        \u_decoder/fir_filter/Q_data_add_3_buff [14]), .C(
        \u_decoder/fir_filter/add_328/carry [14]), .Q(
        \u_decoder/fir_filter/Q_data_add_2 [14]) );
  XOR31 \u_decoder/fir_filter/add_329/U1_14  ( .A(
        \u_decoder/fir_filter/Q_data_mult_3_buff [14]), .B(
        \u_decoder/fir_filter/Q_data_add_4_buff [14]), .C(
        \u_decoder/fir_filter/add_329/carry [14]), .Q(
        \u_decoder/fir_filter/Q_data_add_3 [14]) );
  XOR31 \u_decoder/fir_filter/add_330/U1_14  ( .A(
        \u_decoder/fir_filter/Q_data_mult_4_buff [14]), .B(
        \u_decoder/fir_filter/Q_data_add_5_buff [14]), .C(
        \u_decoder/fir_filter/add_330/carry [14]), .Q(
        \u_decoder/fir_filter/Q_data_add_4 [14]) );
  XOR31 \u_decoder/fir_filter/add_331/U1_14  ( .A(
        \u_decoder/fir_filter/Q_data_mult_5_buff [14]), .B(
        \u_decoder/fir_filter/Q_data_add_6_buff [14]), .C(
        \u_decoder/fir_filter/add_331/carry [14]), .Q(
        \u_decoder/fir_filter/Q_data_add_5 [14]) );
  XOR31 \u_decoder/fir_filter/add_332/U1_14  ( .A(
        \u_decoder/fir_filter/Q_data_mult_6_buff [14]), .B(
        \u_decoder/fir_filter/Q_data_add_7_buff [14]), .C(
        \u_decoder/fir_filter/add_332/carry [14]), .Q(
        \u_decoder/fir_filter/Q_data_add_6 [14]) );
  XOR31 \u_decoder/fir_filter/add_333/U1_14  ( .A(
        \u_decoder/fir_filter/Q_data_mult_7_buff [14]), .B(
        \u_decoder/fir_filter/Q_data_mult_8_buff [14]), .C(
        \u_decoder/fir_filter/add_333/carry [14]), .Q(
        \u_decoder/fir_filter/Q_data_add_7 [14]) );
  XOR31 \u_decoder/fir_filter/add_298/U1_14  ( .A(
        \u_decoder/fir_filter/I_data_mult_4_buff [14]), .B(
        \u_decoder/fir_filter/I_data_add_5_buff [14]), .C(
        \u_decoder/fir_filter/add_298/carry [14]), .Q(
        \u_decoder/fir_filter/I_data_add_4 [14]) );
  XOR31 \u_decoder/fir_filter/add_299/U1_14  ( .A(
        \u_decoder/fir_filter/I_data_mult_5_buff [14]), .B(
        \u_decoder/fir_filter/I_data_add_6_buff [14]), .C(
        \u_decoder/fir_filter/add_299/carry [14]), .Q(
        \u_decoder/fir_filter/I_data_add_5 [14]) );
  XOR31 \u_decoder/fir_filter/add_300/U1_14  ( .A(
        \u_decoder/fir_filter/I_data_mult_6_buff [14]), .B(
        \u_decoder/fir_filter/I_data_add_7_buff [14]), .C(
        \u_decoder/fir_filter/add_300/carry [14]), .Q(
        \u_decoder/fir_filter/I_data_add_6 [14]) );
  XOR31 \u_decoder/fir_filter/add_301/U1_14  ( .A(
        \u_decoder/fir_filter/I_data_mult_7_buff [14]), .B(
        \u_decoder/fir_filter/I_data_mult_8_buff [14]), .C(
        \u_decoder/fir_filter/add_301/carry [14]), .Q(
        \u_decoder/fir_filter/I_data_add_7 [14]) );
  XOR31 \u_cordic/my_rotation/sub_40/U2_15  ( .A(
        \u_cordic/my_rotation/present_angle[0][15] ), .B(n309), .C(
        \u_cordic/my_rotation/sub_40/carry [15]), .Q(
        \u_cordic/my_rotation/next_delta [15]) );
  XOR31 \u_decoder/iq_demod/dp_cluster_0/sub_153/U2_7  ( .A(
        \u_decoder/iq_demod/dp_cluster_0/mult_I_cos_out [7]), .B(n342), .C(
        \u_decoder/iq_demod/dp_cluster_0/sub_153/carry [7]), .Q(
        \u_decoder/iq_demod/add_I_out [7]) );
  XOR31 \u_decoder/iq_demod/dp_cluster_1/add_154/U1_7  ( .A(
        \u_decoder/iq_demod/dp_cluster_1/mult_I_sin_out [7]), .B(
        \u_decoder/iq_demod/dp_cluster_1/mult_Q_cos_out [7]), .C(
        \u_decoder/iq_demod/dp_cluster_1/add_154/carry [7]), .Q(
        \u_decoder/iq_demod/add_Q_out [7]) );
  ADD32 \u_cordic/mycordic/r144/U1_3  ( .A(
        \u_cordic/mycordic/present_I_table[1][3] ), .B(
        \u_cordic/mycordic/present_Q_table[1][3] ), .CI(n2), .CO(
        \u_cordic/mycordic/r144/carry [4]), .S(\u_cordic/mycordic/N255 ) );
  ADD32 \u_cordic/mycordic/sub_182/U2_3  ( .A(
        \u_cordic/mycordic/present_I_table[1][3] ), .B(n224), .CI(n1), .CO(
        \u_cordic/mycordic/sub_182/carry [4]), .S(\u_cordic/mycordic/N287 ) );
  ADD32 \u_cordic/mycordic/sub_178/U2_3  ( .A(
        \u_cordic/mycordic/present_Q_table[1][3] ), .B(n223), .CI(n1), .CO(
        \u_cordic/mycordic/sub_178/carry [4]), .S(\u_cordic/mycordic/N263 ) );
  LOGIC1 U2 ( .Q(n1) );
  LOGIC0 U3 ( .Q(n2) );
  XOR21 U4 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_276/SUMB[7][3] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[7][2] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/A1[8] ) );
  XOR21 U5 ( .A(\u_decoder/fir_filter/dp_cluster_0/r167/SUMB[7][3] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[7][2] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r167/A1[8] ) );
  XOR21 U6 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_308/SUMB[7][3] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[7][2] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/A1[8] ) );
  XOR21 U7 ( .A(\u_decoder/fir_filter/dp_cluster_0/r180/SUMB[7][3] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[7][2] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r180/A1[8] ) );
  NAND31 U8 ( .A(\u_inFIFO/j_FIFO [1]), .B(\u_inFIFO/j_FIFO [0]), .C(
        \u_inFIFO/j_FIFO [2]), .Q(\u_inFIFO/n142 ) );
  NAND31 U9 ( .A(\u_inFIFO/j_FIFO [0]), .B(\u_inFIFO/n100 ), .C(
        \u_inFIFO/j_FIFO [2]), .Q(\u_inFIFO/n136 ) );
  NAND31 U10 ( .A(\u_inFIFO/n101 ), .B(\u_inFIFO/n100 ), .C(
        \u_inFIFO/j_FIFO [2]), .Q(\u_inFIFO/n133 ) );
  NAND31 U11 ( .A(\u_inFIFO/j_FIFO [0]), .B(\u_inFIFO/n99 ), .C(
        \u_inFIFO/j_FIFO [1]), .Q(\u_inFIFO/n130 ) );
  NAND31 U12 ( .A(\u_inFIFO/n100 ), .B(\u_inFIFO/n99 ), .C(
        \u_inFIFO/j_FIFO [0]), .Q(\u_inFIFO/n124 ) );
  NAND31 U13 ( .A(\u_inFIFO/n100 ), .B(\u_inFIFO/n99 ), .C(\u_inFIFO/n101 ), 
        .Q(\u_inFIFO/n120 ) );
  NAND31 U14 ( .A(\u_inFIFO/j_FIFO [1]), .B(\u_inFIFO/n101 ), .C(
        \u_inFIFO/j_FIFO [2]), .Q(\u_inFIFO/n139 ) );
  NAND31 U15 ( .A(\u_inFIFO/n101 ), .B(\u_inFIFO/n99 ), .C(
        \u_inFIFO/j_FIFO [1]), .Q(\u_inFIFO/n127 ) );
  NOR21 U16 ( .A(n678), .B(n679), .Q(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/A2[5] ) );
  INV3 U17 ( .A(\u_cordic/mycordic/n353 ), .Q(n1178) );
  INV3 U18 ( .A(\u_decoder/fir_filter/n1084 ), .Q(n1822) );
  INV3 U19 ( .A(\u_decoder/fir_filter/n787 ), .Q(n1893) );
  NOR21 U20 ( .A(\u_coder/n315 ), .B(n369), .Q(\u_coder/N522 ) );
  BUF2 U21 ( .A(\u_decoder/I_prefilter [7]), .Q(n961) );
  BUF2 U22 ( .A(\u_decoder/Q_prefilter [7]), .Q(n963) );
  BUF2 U23 ( .A(\u_decoder/I_prefilter [7]), .Q(n960) );
  BUF2 U24 ( .A(\u_decoder/Q_prefilter [7]), .Q(n962) );
  BUF2 U25 ( .A(\u_decoder/I_prefilter [6]), .Q(n764) );
  BUF2 U26 ( .A(\u_decoder/Q_prefilter [6]), .Q(n754) );
  BUF2 U27 ( .A(\u_decoder/I_prefilter [5]), .Q(n765) );
  BUF2 U28 ( .A(\u_decoder/Q_prefilter [5]), .Q(n755) );
  BUF2 U29 ( .A(\u_decoder/Q_prefilter [3]), .Q(n759) );
  BUF2 U30 ( .A(\u_decoder/I_prefilter [3]), .Q(n769) );
  BUF2 U31 ( .A(\u_decoder/Q_prefilter [4]), .Q(n757) );
  BUF2 U32 ( .A(\u_decoder/I_prefilter [4]), .Q(n767) );
  BUF2 U33 ( .A(\u_decoder/Q_prefilter [3]), .Q(n758) );
  BUF2 U34 ( .A(\u_decoder/I_prefilter [3]), .Q(n768) );
  XNR21 U35 ( .A(n305), .B(\u_cordic/mycordic/sub_add_150_b0/carry [7]), .Q(
        n39) );
  XNR21 U36 ( .A(n963), .B(n1910), .Q(n47) );
  XNR21 U37 ( .A(n961), .B(n1839), .Q(n48) );
  XNR21 U38 ( .A(n2406), .B(n2407), .Q(n49) );
  XNR21 U39 ( .A(n2493), .B(n2494), .Q(n50) );
  XOR21 U40 ( .A(n2387), .B(n2388), .Q(n55) );
  XOR21 U41 ( .A(n2474), .B(n2475), .Q(n56) );
  XNR31 U42 ( .A(\u_decoder/fir_filter/dp_cluster_0/r177/A2[7] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r177/A1[7] ), .C(n2346), .Q(n57) );
  XNR31 U43 ( .A(\u_decoder/fir_filter/dp_cluster_0/r164/A2[7] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r164/A1[7] ), .C(n2433), .Q(n58) );
  XNR21 U44 ( .A(n2366), .B(n2367), .Q(n65) );
  XNR21 U45 ( .A(n2453), .B(n2454), .Q(n66) );
  XOR21 U46 ( .A(\u_decoder/iq_demod/dp_cluster_0/mult_151/A1[2] ), .B(n1949), 
        .Q(n67) );
  XNR21 U47 ( .A(\u_cordic/mycordic/present_ANGLE_table[6][15] ), .B(
        \u_cordic/mycordic/r173/carry [15]), .Q(n76) );
  XOR21 U48 ( .A(\u_decoder/fir_filter/dp_cluster_0/r177/A1[5] ), .B(n2353), 
        .Q(n107) );
  XOR21 U49 ( .A(\u_decoder/fir_filter/dp_cluster_0/r164/A1[5] ), .B(n2440), 
        .Q(n108) );
  XOR21 U50 ( .A(n2342), .B(n2343), .Q(n109) );
  XNR21 U51 ( .A(\u_decoder/iq_demod/dp_cluster_0/mult_151/ab[0][1] ), .B(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/ab[1][0] ), .Q(n139) );
  MUX22 U52 ( .A(\u_cordic/mycordic/present_C_table[7][1] ), .B(n751), .S(n781), .Q(n153) );
  XNR21 U53 ( .A(\u_cordic/mycordic/n110 ), .B(
        \u_cordic/mycordic/present_C_table[7][0] ), .Q(n166) );
  IMUX40 U54 ( .A(\u_inFIFO/N183 ), .B(\u_inFIFO/N181 ), .C(\u_inFIFO/N182 ), 
        .D(\u_inFIFO/N180 ), .S0(\u_inFIFO/N39 ), .S1(\u_inFIFO/N38 ), .Q(n233) );
  BUF2 U55 ( .A(\u_decoder/fir_filter/n721 ), .Q(n933) );
  BUF2 U56 ( .A(\u_decoder/fir_filter/n721 ), .Q(n938) );
  BUF2 U57 ( .A(\u_decoder/fir_filter/n721 ), .Q(n936) );
  BUF2 U58 ( .A(\u_decoder/fir_filter/n721 ), .Q(n937) );
  BUF2 U59 ( .A(\u_decoder/fir_filter/n721 ), .Q(n935) );
  BUF2 U60 ( .A(\u_decoder/fir_filter/n721 ), .Q(n934) );
  NAND22 U61 ( .A(n978), .B(\u_coder/n314 ), .Q(\u_coder/n315 ) );
  NAND22 U62 ( .A(n978), .B(\u_coder/n314 ), .Q(n814) );
  BUF2 U63 ( .A(\u_decoder/fir_filter/I_data_mult_0 [0]), .Q(n772) );
  BUF2 U64 ( .A(\u_decoder/fir_filter/Q_data_mult_0 [0]), .Q(n762) );
  BUF2 U65 ( .A(\u_decoder/I_prefilter [2]), .Q(n770) );
  BUF2 U66 ( .A(\u_decoder/Q_prefilter [2]), .Q(n760) );
  BUF2 U67 ( .A(\u_decoder/fir_filter/I_data_mult_0 [0]), .Q(n773) );
  BUF2 U68 ( .A(\u_decoder/fir_filter/Q_data_mult_0 [0]), .Q(n763) );
  BUF2 U69 ( .A(\u_decoder/I_prefilter [2]), .Q(n771) );
  BUF2 U70 ( .A(\u_decoder/Q_prefilter [2]), .Q(n761) );
  AOI221 U71 ( .A(\u_decoder/fir_filter/I_data_mult_4 [14]), .B(n837), .C(
        \u_decoder/fir_filter/I_data_mult_4_buff [14]), .D(n927), .Q(
        \u_decoder/fir_filter/n1084 ) );
  AOI221 U72 ( .A(\u_decoder/fir_filter/Q_data_mult_4 [14]), .B(n837), .C(
        \u_decoder/fir_filter/Q_data_mult_4_buff [14]), .D(n932), .Q(
        \u_decoder/fir_filter/n787 ) );
  BUF2 U73 ( .A(\u_cordic/mycordic/present_Q_table[4][7] ), .Q(n749) );
  NOR21 U74 ( .A(\u_outFIFO/n197 ), .B(n983), .Q(\u_outFIFO/n514 ) );
  NOR21 U75 ( .A(n981), .B(\u_inFIFO/sigEnableCounter ), .Q(\u_inFIFO/n202 )
         );
  BUF2 U76 ( .A(\u_inFIFO/N36 ), .Q(n780) );
  AOI221 U77 ( .A(n1575), .B(\u_cordic/mycordic/N247 ), .C(n784), .D(
        \u_cordic/mycordic/present_Q_table[0][7] ), .Q(
        \u_cordic/mycordic/n353 ) );
  INV3 U78 ( .A(\u_cordic/mycordic/n537 ), .Q(n1579) );
  BUF2 U79 ( .A(\u_cordic/mycordic/n345 ), .Q(n787) );
  BUF2 U80 ( .A(\u_outFIFO/N38 ), .Q(n775) );
  INV3 U81 ( .A(in_MUX_inSEL6[0]), .Q(n1689) );
  INV3 U82 ( .A(n857), .Q(n837) );
  INV3 U83 ( .A(n856), .Q(n838) );
  INV3 U84 ( .A(n856), .Q(n839) );
  INV3 U85 ( .A(n856), .Q(n840) );
  BUF2 U86 ( .A(n909), .Q(n856) );
  BUF2 U87 ( .A(n909), .Q(n857) );
  INV3 U88 ( .A(n854), .Q(n845) );
  INV3 U89 ( .A(n854), .Q(n846) );
  INV3 U90 ( .A(n853), .Q(n847) );
  INV3 U91 ( .A(n853), .Q(n848) );
  INV3 U92 ( .A(n853), .Q(n849) );
  INV3 U93 ( .A(n855), .Q(n841) );
  INV3 U94 ( .A(n855), .Q(n842) );
  INV3 U95 ( .A(n855), .Q(n843) );
  INV3 U96 ( .A(n854), .Q(n844) );
  INV3 U97 ( .A(n852), .Q(n850) );
  INV3 U98 ( .A(n852), .Q(n851) );
  BUF2 U99 ( .A(n908), .Q(n859) );
  BUF2 U100 ( .A(n908), .Q(n858) );
  BUF2 U101 ( .A(n907), .Q(n860) );
  BUF2 U102 ( .A(n899), .Q(n876) );
  BUF2 U103 ( .A(n899), .Q(n877) );
  BUF2 U104 ( .A(n898), .Q(n878) );
  BUF2 U105 ( .A(n898), .Q(n879) );
  BUF2 U106 ( .A(n897), .Q(n880) );
  BUF2 U107 ( .A(n897), .Q(n881) );
  BUF2 U108 ( .A(n896), .Q(n882) );
  BUF2 U109 ( .A(n896), .Q(n883) );
  BUF2 U110 ( .A(n895), .Q(n884) );
  BUF2 U111 ( .A(n895), .Q(n885) );
  BUF2 U112 ( .A(n894), .Q(n886) );
  BUF2 U113 ( .A(n894), .Q(n887) );
  BUF2 U114 ( .A(n893), .Q(n888) );
  BUF2 U115 ( .A(n893), .Q(n889) );
  BUF2 U116 ( .A(n892), .Q(n890) );
  BUF2 U117 ( .A(n907), .Q(n861) );
  BUF2 U118 ( .A(n906), .Q(n862) );
  BUF2 U119 ( .A(n906), .Q(n863) );
  BUF2 U120 ( .A(n905), .Q(n864) );
  BUF2 U121 ( .A(n905), .Q(n865) );
  BUF2 U122 ( .A(n904), .Q(n866) );
  BUF2 U123 ( .A(n904), .Q(n867) );
  BUF2 U124 ( .A(n903), .Q(n868) );
  BUF2 U125 ( .A(n903), .Q(n869) );
  BUF2 U126 ( .A(n902), .Q(n870) );
  BUF2 U127 ( .A(n902), .Q(n871) );
  BUF2 U128 ( .A(n901), .Q(n872) );
  BUF2 U129 ( .A(n901), .Q(n873) );
  BUF2 U130 ( .A(n900), .Q(n874) );
  BUF2 U131 ( .A(n900), .Q(n875) );
  BUF2 U132 ( .A(n892), .Q(n891) );
  AOI211 U133 ( .A(n2474), .B(n1841), .C(n1843), .Q(n2493) );
  INV3 U134 ( .A(n2476), .Q(n1843) );
  AOI211 U135 ( .A(n2387), .B(n1912), .C(n1914), .Q(n2406) );
  INV3 U136 ( .A(n2389), .Q(n1914) );
  INV3 U137 ( .A(n2513), .Q(n1826) );
  INV3 U138 ( .A(n2426), .Q(n1897) );
  NAND22 U139 ( .A(n1838), .B(n2490), .Q(n2494) );
  INV3 U140 ( .A(n2487), .Q(n1838) );
  NAND22 U141 ( .A(n1909), .B(n2403), .Q(n2407) );
  INV3 U142 ( .A(n2400), .Q(n1909) );
  AOI211 U143 ( .A(n2496), .B(n1825), .C(n1827), .Q(n2515) );
  INV3 U144 ( .A(n2498), .Q(n1827) );
  AOI211 U145 ( .A(n2409), .B(n1896), .C(n1898), .Q(n2428) );
  INV3 U146 ( .A(n2411), .Q(n1898) );
  INV3 U147 ( .A(n2477), .Q(n1845) );
  INV3 U148 ( .A(n2390), .Q(n1916) );
  INV3 U149 ( .A(n2508), .Q(n1825) );
  INV3 U150 ( .A(n2421), .Q(n1896) );
  NAND22 U151 ( .A(n1841), .B(n2476), .Q(n2475) );
  NAND22 U152 ( .A(n1912), .B(n2389), .Q(n2388) );
  INV3 U153 ( .A(n2491), .Q(n1842) );
  INV3 U154 ( .A(n2404), .Q(n1913) );
  INV3 U155 ( .A(n2509), .Q(n1820) );
  INV3 U156 ( .A(n2422), .Q(n1891) );
  INV3 U157 ( .A(n2486), .Q(n1841) );
  INV3 U158 ( .A(n2399), .Q(n1912) );
  BUF2 U159 ( .A(n912), .Q(n909) );
  BUF2 U160 ( .A(n911), .Q(n853) );
  BUF2 U161 ( .A(n910), .Q(n855) );
  BUF2 U162 ( .A(n910), .Q(n854) );
  BUF2 U163 ( .A(n911), .Q(n852) );
  BUF2 U164 ( .A(n1460), .Q(n815) );
  BUF2 U165 ( .A(n1460), .Q(n830) );
  BUF2 U166 ( .A(n1460), .Q(n829) );
  BUF2 U167 ( .A(n1460), .Q(n828) );
  BUF2 U168 ( .A(n1460), .Q(n827) );
  BUF2 U169 ( .A(n1460), .Q(n826) );
  BUF2 U170 ( .A(n1460), .Q(n825) );
  BUF2 U171 ( .A(n1460), .Q(n824) );
  BUF2 U172 ( .A(n1460), .Q(n823) );
  BUF2 U173 ( .A(n1460), .Q(n822) );
  BUF2 U174 ( .A(n1460), .Q(n821) );
  BUF2 U175 ( .A(n1460), .Q(n820) );
  BUF2 U176 ( .A(n1460), .Q(n819) );
  BUF2 U177 ( .A(n1460), .Q(n818) );
  BUF2 U178 ( .A(n1460), .Q(n817) );
  BUF2 U179 ( .A(n1460), .Q(n816) );
  BUF2 U180 ( .A(n904), .Q(n899) );
  BUF2 U181 ( .A(n908), .Q(n898) );
  BUF2 U182 ( .A(n906), .Q(n897) );
  BUF2 U183 ( .A(n908), .Q(n896) );
  BUF2 U184 ( .A(n907), .Q(n895) );
  BUF2 U185 ( .A(n908), .Q(n894) );
  BUF2 U186 ( .A(n856), .Q(n893) );
  BUF2 U187 ( .A(n893), .Q(n892) );
  BUF2 U188 ( .A(n856), .Q(n907) );
  BUF2 U189 ( .A(n856), .Q(n906) );
  BUF2 U190 ( .A(n856), .Q(n905) );
  BUF2 U191 ( .A(n856), .Q(n904) );
  BUF2 U192 ( .A(n908), .Q(n903) );
  BUF2 U193 ( .A(n908), .Q(n902) );
  BUF2 U194 ( .A(n912), .Q(n908) );
  BUF2 U195 ( .A(n905), .Q(n901) );
  BUF2 U196 ( .A(n908), .Q(n900) );
  INV3 U197 ( .A(n955), .Q(n948) );
  INV3 U198 ( .A(n955), .Q(n949) );
  INV3 U199 ( .A(n955), .Q(n950) );
  INV3 U200 ( .A(n956), .Q(n951) );
  INV3 U201 ( .A(n956), .Q(n952) );
  INV3 U202 ( .A(n957), .Q(n953) );
  INV3 U203 ( .A(n958), .Q(n954) );
  NOR21 U204 ( .A(\u_decoder/fir_filter/dp_cluster_0/r167/A1[8] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r167/A2[8] ), .Q(n2495) );
  NOR21 U205 ( .A(\u_decoder/fir_filter/dp_cluster_0/r180/A1[8] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r180/A2[8] ), .Q(n2408) );
  AOI211 U206 ( .A(n2452), .B(\u_decoder/fir_filter/dp_cluster_0/r165/A1[7] ), 
        .C(n1805), .Q(n2451) );
  INV3 U207 ( .A(n2463), .Q(n1805) );
  AOI211 U208 ( .A(n2365), .B(\u_decoder/fir_filter/dp_cluster_0/r178/A1[7] ), 
        .C(n1876), .Q(n2364) );
  INV3 U209 ( .A(n2376), .Q(n1876) );
  INV3 U210 ( .A(\u_decoder/fir_filter/dp_cluster_0/r165/A1[9] ), .Q(n1801) );
  INV3 U211 ( .A(n2450), .Q(n1802) );
  INV3 U212 ( .A(\u_decoder/fir_filter/dp_cluster_0/r178/A1[9] ), .Q(n1872) );
  INV3 U213 ( .A(n2363), .Q(n1873) );
  INV3 U214 ( .A(\u_decoder/fir_filter/dp_cluster_0/r164/A1[6] ), .Q(n1855) );
  INV3 U215 ( .A(\u_decoder/fir_filter/dp_cluster_0/r177/A1[6] ), .Q(n1926) );
  NOR21 U216 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_276/A2[9] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/A1[9] ), .Q(n2508) );
  NOR21 U217 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_308/A2[9] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/A1[9] ), .Q(n2421) );
  INV3 U218 ( .A(\u_decoder/fir_filter/dp_cluster_0/r164/A1[8] ), .Q(n1860) );
  INV3 U219 ( .A(n2432), .Q(n1853) );
  INV3 U220 ( .A(\u_decoder/fir_filter/dp_cluster_0/r177/A1[8] ), .Q(n1931) );
  INV3 U221 ( .A(n2345), .Q(n1924) );
  XNR21 U222 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_276/A1[8] ), .B(
        n2499), .Q(n2502) );
  XNR21 U223 ( .A(\u_decoder/fir_filter/dp_cluster_0/r167/A1[8] ), .B(n2477), 
        .Q(n2480) );
  XNR21 U224 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_308/A1[8] ), .B(
        n2412), .Q(n2415) );
  XNR21 U225 ( .A(\u_decoder/fir_filter/dp_cluster_0/r180/A1[8] ), .B(n2390), 
        .Q(n2393) );
  INV3 U226 ( .A(n2466), .Q(n1811) );
  INV3 U227 ( .A(n2451), .Q(n1804) );
  INV3 U228 ( .A(n2379), .Q(n1882) );
  INV3 U229 ( .A(n2364), .Q(n1875) );
  INV3 U230 ( .A(\u_decoder/fir_filter/I_data_mult_3 [10]), .Q(n1844) );
  IMUX21 U231 ( .A(n2480), .B(n2481), .S(
        \u_decoder/fir_filter/dp_cluster_0/r167/A2[8] ), .Q(n2479) );
  NOR21 U232 ( .A(\u_decoder/fir_filter/dp_cluster_0/r167/A1[8] ), .B(n1845), 
        .Q(n2481) );
  INV3 U233 ( .A(\u_decoder/fir_filter/Q_data_mult_3 [10]), .Q(n1915) );
  IMUX21 U234 ( .A(n2393), .B(n2394), .S(
        \u_decoder/fir_filter/dp_cluster_0/r180/A2[8] ), .Q(n2392) );
  NOR21 U235 ( .A(\u_decoder/fir_filter/dp_cluster_0/r180/A1[8] ), .B(n1916), 
        .Q(n2394) );
  NOR21 U236 ( .A(n570), .B(n571), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r167/A2[7] ) );
  INV3 U237 ( .A(\u_decoder/fir_filter/dp_cluster_0/r167/SUMB[7][1] ), .Q(n571) );
  INV3 U238 ( .A(\u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[7][0] ), .Q(
        n570) );
  NOR21 U239 ( .A(n632), .B(n633), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r180/A2[7] ) );
  INV3 U240 ( .A(\u_decoder/fir_filter/dp_cluster_0/r180/SUMB[7][1] ), .Q(n633) );
  INV3 U241 ( .A(\u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[7][0] ), .Q(
        n632) );
  XNR31 U242 ( .A(\u_decoder/fir_filter/dp_cluster_0/r165/A2[10] ), .B(n1868), 
        .C(n2459), .Q(n316) );
  XNR31 U243 ( .A(\u_decoder/fir_filter/dp_cluster_0/r178/A2[10] ), .B(n1939), 
        .C(n2372), .Q(n317) );
  XNR31 U244 ( .A(\u_decoder/fir_filter/dp_cluster_0/r164/A2[9] ), .B(n1868), 
        .C(n2431), .Q(n318) );
  XNR31 U245 ( .A(\u_decoder/fir_filter/dp_cluster_0/r177/A2[9] ), .B(n1939), 
        .C(n2344), .Q(n319) );
  NOR21 U246 ( .A(n1855), .B(n1857), .Q(n2448) );
  NOR21 U247 ( .A(n1926), .B(n1928), .Q(n2361) );
  XNR21 U248 ( .A(\u_decoder/fir_filter/dp_cluster_0/r167/SUMB[7][1] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[7][0] ), .Q(n320) );
  XNR21 U249 ( .A(\u_decoder/fir_filter/dp_cluster_0/r180/SUMB[7][1] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[7][0] ), .Q(n321) );
  AOI211 U250 ( .A(n1814), .B(\u_decoder/fir_filter/dp_cluster_0/r166/A1[7] ), 
        .C(n1812), .Q(n2466) );
  INV3 U251 ( .A(n2472), .Q(n1812) );
  AOI211 U252 ( .A(n1885), .B(\u_decoder/fir_filter/dp_cluster_0/r179/A1[7] ), 
        .C(n1883), .Q(n2379) );
  INV3 U253 ( .A(n2385), .Q(n1883) );
  NOR21 U254 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_276/A1[8] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/A2[8] ), .Q(n2517) );
  NOR21 U255 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_308/A1[8] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/A2[8] ), .Q(n2430) );
  NOR21 U256 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_276/A1[8] ), .B(
        n1829), .Q(n2503) );
  INV3 U257 ( .A(n2499), .Q(n1829) );
  NOR21 U258 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_308/A1[8] ), .B(
        n1900), .Q(n2416) );
  INV3 U259 ( .A(n2412), .Q(n1900) );
  NOR21 U260 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_276/A2[10] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/A1[10] ), .Q(n2509) );
  NOR21 U261 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_308/A2[10] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/A1[10] ), .Q(n2422) );
  NAND22 U262 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_276/A2[8] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/A1[8] ), .Q(n2500) );
  NAND22 U263 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_308/A2[8] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/A1[8] ), .Q(n2413) );
  NAND22 U264 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_276/A2[9] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/A1[9] ), .Q(n2498) );
  NAND22 U265 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_308/A2[9] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/A1[9] ), .Q(n2411) );
  NAND22 U266 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_276/A2[10] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/A1[10] ), .Q(n2512) );
  NAND22 U267 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_308/A2[10] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/A1[10] ), .Q(n2425) );
  XNR31 U268 ( .A(\u_decoder/fir_filter/dp_cluster_0/r165/A2[9] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r165/A1[9] ), .C(n2450), .Q(n322)
         );
  XNR31 U269 ( .A(\u_decoder/fir_filter/dp_cluster_0/r178/A2[9] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r178/A1[9] ), .C(n2363), .Q(n323)
         );
  XOR31 U270 ( .A(\u_decoder/fir_filter/dp_cluster_0/r164/A2[8] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r164/A1[8] ), .C(n2432), .Q(n324)
         );
  XOR31 U271 ( .A(\u_decoder/fir_filter/dp_cluster_0/r177/A2[8] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r177/A1[8] ), .C(n2345), .Q(n325)
         );
  INV3 U272 ( .A(\u_decoder/fir_filter/dp_cluster_0/r166/A1[8] ), .Q(n1810) );
  INV3 U273 ( .A(\u_decoder/fir_filter/dp_cluster_0/r179/A1[8] ), .Q(n1881) );
  NAND31 U274 ( .A(n1122), .B(n1041), .C(n1123), .Q(n1044) );
  NAND22 U275 ( .A(\u_decoder/fir_filter/dp_cluster_0/r167/A2[8] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r167/A1[8] ), .Q(n2478) );
  NAND22 U276 ( .A(\u_decoder/fir_filter/dp_cluster_0/r180/A2[8] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r180/A1[8] ), .Q(n2391) );
  XNR31 U277 ( .A(\u_decoder/fir_filter/dp_cluster_0/r166/A2[8] ), .B(n1810), 
        .C(n2466), .Q(n326) );
  XNR31 U278 ( .A(\u_decoder/fir_filter/dp_cluster_0/r166/A2[7] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r166/A1[7] ), .C(n1814), .Q(n327)
         );
  XNR31 U279 ( .A(\u_decoder/fir_filter/dp_cluster_0/r165/A2[8] ), .B(n1803), 
        .C(n2451), .Q(n328) );
  XNR31 U280 ( .A(\u_decoder/fir_filter/dp_cluster_0/r179/A2[8] ), .B(n1881), 
        .C(n2379), .Q(n329) );
  XNR31 U281 ( .A(\u_decoder/fir_filter/dp_cluster_0/r179/A2[7] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r179/A1[7] ), .C(n1885), .Q(n330)
         );
  XNR31 U282 ( .A(\u_decoder/fir_filter/dp_cluster_0/r178/A2[8] ), .B(n1874), 
        .C(n2364), .Q(n331) );
  INV3 U283 ( .A(\u_decoder/fir_filter/dp_cluster_0/r165/A1[8] ), .Q(n1803) );
  INV3 U284 ( .A(\u_decoder/fir_filter/dp_cluster_0/r178/A1[8] ), .Q(n1874) );
  NOR21 U285 ( .A(\u_decoder/fir_filter/dp_cluster_0/r167/A2[10] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r167/A1[10] ), .Q(n2487) );
  NOR21 U286 ( .A(\u_decoder/fir_filter/dp_cluster_0/r180/A2[10] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r180/A1[10] ), .Q(n2400) );
  NOR21 U287 ( .A(\u_decoder/fir_filter/dp_cluster_0/r164/A1[6] ), .B(n1857), 
        .Q(n2439) );
  NOR21 U288 ( .A(\u_decoder/fir_filter/dp_cluster_0/r177/A1[6] ), .B(n1928), 
        .Q(n2352) );
  NOR21 U289 ( .A(\u_decoder/fir_filter/dp_cluster_0/r167/A2[9] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r167/A1[9] ), .Q(n2486) );
  NOR21 U290 ( .A(\u_decoder/fir_filter/dp_cluster_0/r180/A2[9] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r180/A1[9] ), .Q(n2399) );
  NAND22 U291 ( .A(\u_decoder/fir_filter/dp_cluster_0/r167/A2[9] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r167/A1[9] ), .Q(n2476) );
  NAND22 U292 ( .A(\u_decoder/fir_filter/dp_cluster_0/r180/A2[9] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r180/A1[9] ), .Q(n2389) );
  XNR31 U293 ( .A(\u_decoder/fir_filter/dp_cluster_0/r167/A1[7] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r167/A2[7] ), .C(n2482), .Q(n332)
         );
  XNR31 U294 ( .A(\u_decoder/fir_filter/dp_cluster_0/r180/A1[7] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r180/A2[7] ), .C(n2395), .Q(n333)
         );
  XNR31 U295 ( .A(\u_decoder/fir_filter/dp_cluster_0/r165/A2[7] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r165/A1[7] ), .C(n2452), .Q(n334)
         );
  XNR31 U296 ( .A(\u_decoder/fir_filter/dp_cluster_0/r178/A2[7] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r178/A1[7] ), .C(n2365), .Q(n335)
         );
  INV3 U297 ( .A(n2436), .Q(n1856) );
  INV3 U298 ( .A(n2349), .Q(n1927) );
  NAND22 U299 ( .A(\u_decoder/fir_filter/dp_cluster_0/r167/A2[10] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r167/A1[10] ), .Q(n2490) );
  NAND22 U300 ( .A(\u_decoder/fir_filter/dp_cluster_0/r180/A2[10] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r180/A1[10] ), .Q(n2403) );
  INV3 U301 ( .A(n2441), .Q(n1858) );
  INV3 U302 ( .A(n2354), .Q(n1929) );
  INV3 U303 ( .A(n933), .Q(n913) );
  INV3 U304 ( .A(\u_coder/n230 ), .Q(n1748) );
  INV3 U305 ( .A(\u_coder/n167 ), .Q(n1709) );
  INV3 U306 ( .A(\u_decoder/fir_filter/n554 ), .Q(n912) );
  BUF6 U307 ( .A(\u_inFIFO/n118 ), .Q(n966) );
  INV3 U308 ( .A(n968), .Q(n967) );
  INV3 U309 ( .A(\u_outFIFO/n502 ), .Q(n1460) );
  BUF2 U310 ( .A(n959), .Q(n958) );
  BUF2 U311 ( .A(n908), .Q(n911) );
  BUF2 U312 ( .A(n908), .Q(n910) );
  BUF2 U313 ( .A(n957), .Q(n955) );
  BUF2 U314 ( .A(n959), .Q(n957) );
  BUF2 U315 ( .A(n957), .Q(n956) );
  INV3 U316 ( .A(n936), .Q(n924) );
  INV3 U317 ( .A(n934), .Q(n919) );
  INV3 U318 ( .A(n934), .Q(n918) );
  INV3 U319 ( .A(n934), .Q(n917) );
  INV3 U320 ( .A(n934), .Q(n916) );
  INV3 U321 ( .A(n937), .Q(n930) );
  INV3 U322 ( .A(n937), .Q(n931) );
  INV3 U323 ( .A(n937), .Q(n928) );
  INV3 U324 ( .A(n936), .Q(n926) );
  INV3 U325 ( .A(n936), .Q(n925) );
  INV3 U326 ( .A(n936), .Q(n927) );
  INV3 U327 ( .A(n937), .Q(n929) );
  INV3 U328 ( .A(n933), .Q(n915) );
  INV3 U329 ( .A(n933), .Q(n914) );
  INV3 U330 ( .A(n935), .Q(n923) );
  INV3 U331 ( .A(n935), .Q(n921) );
  INV3 U332 ( .A(n935), .Q(n920) );
  INV3 U333 ( .A(n935), .Q(n922) );
  INV3 U334 ( .A(n938), .Q(n932) );
  XOR21 U335 ( .A(\u_decoder/fir_filter/dp_cluster_0/r164/SUMB[7][1] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r164/CARRYB[7][0] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r164/A1[6] ) );
  XOR21 U336 ( .A(\u_decoder/fir_filter/dp_cluster_0/r177/SUMB[7][1] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r177/CARRYB[7][0] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r177/A1[6] ) );
  NOR40 U337 ( .A(n2486), .B(n2477), .C(n2487), .D(n2488), .Q(n2485) );
  NOR40 U338 ( .A(n2399), .B(n2390), .C(n2400), .D(n2401), .Q(n2398) );
  AOI311 U339 ( .A(n2446), .B(\u_decoder/fir_filter/dp_cluster_0/r164/A1[4] ), 
        .C(\u_decoder/fir_filter/dp_cluster_0/r164/A1[5] ), .D(n2447), .Q(
        n2432) );
  NOR21 U340 ( .A(n2449), .B(n2441), .Q(n2446) );
  MAJ31 U341 ( .A(\u_decoder/fir_filter/dp_cluster_0/r164/A2[7] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r164/A1[7] ), .C(n2448), .Q(n2447)
         );
  AOI311 U342 ( .A(n2359), .B(\u_decoder/fir_filter/dp_cluster_0/r177/A1[4] ), 
        .C(\u_decoder/fir_filter/dp_cluster_0/r177/A1[5] ), .D(n2360), .Q(
        n2345) );
  NOR21 U343 ( .A(n2362), .B(n2354), .Q(n2359) );
  MAJ31 U344 ( .A(\u_decoder/fir_filter/dp_cluster_0/r177/A2[7] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r177/A1[7] ), .C(n2361), .Q(n2360)
         );
  XOR21 U345 ( .A(\u_decoder/fir_filter/dp_cluster_0/r166/SUMB[7][1] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r166/CARRYB[7][0] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r166/A1[6] ) );
  XOR21 U346 ( .A(\u_decoder/fir_filter/dp_cluster_0/r179/SUMB[7][1] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r179/CARRYB[7][0] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r179/A1[6] ) );
  XOR21 U347 ( .A(\u_decoder/fir_filter/dp_cluster_0/r165/SUMB[7][1] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r165/CARRYB[7][0] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r165/A1[6] ) );
  XOR21 U348 ( .A(\u_decoder/fir_filter/dp_cluster_0/r178/SUMB[7][1] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r178/CARRYB[7][0] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r178/A1[6] ) );
  OAI311 U349 ( .A(n1806), .B(n2456), .C(n2455), .D(n2464), .Q(n2452) );
  NAND22 U350 ( .A(\u_decoder/fir_filter/dp_cluster_0/r165/A2[6] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r165/A1[6] ), .Q(n2464) );
  OAI311 U351 ( .A(n1877), .B(n2369), .C(n2368), .D(n2377), .Q(n2365) );
  NAND22 U352 ( .A(\u_decoder/fir_filter/dp_cluster_0/r178/A2[6] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r178/A1[6] ), .Q(n2377) );
  XOR21 U353 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_276/SUMB[7][4] ), 
        .B(\u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[7][3] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/A1[9] ) );
  XOR21 U354 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_308/SUMB[7][4] ), 
        .B(\u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[7][3] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/A1[9] ) );
  XOR21 U355 ( .A(\u_decoder/fir_filter/dp_cluster_0/r164/SUMB[7][2] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r164/CARRYB[7][1] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r164/A1[7] ) );
  XOR21 U356 ( .A(\u_decoder/fir_filter/dp_cluster_0/r177/SUMB[7][2] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r177/CARRYB[7][1] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r177/A1[7] ) );
  XOR21 U357 ( .A(\u_decoder/fir_filter/dp_cluster_0/r167/SUMB[6][1] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[6][0] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r167/SUMB[7][0] ) );
  XOR21 U358 ( .A(\u_decoder/fir_filter/dp_cluster_0/r180/SUMB[6][1] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[6][0] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r180/SUMB[7][0] ) );
  XOR21 U359 ( .A(\u_decoder/fir_filter/dp_cluster_0/r165/SUMB[4][3] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r165/CARRYB[6][0] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r165/SUMB[7][0] ) );
  XOR21 U360 ( .A(\u_decoder/fir_filter/dp_cluster_0/r178/SUMB[4][3] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r178/CARRYB[6][0] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r178/SUMB[7][0] ) );
  XOR21 U361 ( .A(\u_decoder/fir_filter/dp_cluster_0/r166/SUMB[7][2] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r166/CARRYB[7][1] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r166/A1[7] ) );
  XOR21 U362 ( .A(\u_decoder/fir_filter/dp_cluster_0/r165/SUMB[7][2] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r165/CARRYB[7][1] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r165/A1[7] ) );
  XOR21 U363 ( .A(\u_decoder/fir_filter/dp_cluster_0/r179/SUMB[7][2] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r179/CARRYB[7][1] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r179/A1[7] ) );
  XOR21 U364 ( .A(\u_decoder/fir_filter/dp_cluster_0/r178/SUMB[7][2] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r178/CARRYB[7][1] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r178/A1[7] ) );
  XOR21 U365 ( .A(\u_decoder/fir_filter/dp_cluster_0/r166/SUMB[5][3] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r166/CARRYB[6][1] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r166/SUMB[7][1] ) );
  XOR21 U366 ( .A(\u_decoder/fir_filter/dp_cluster_0/r179/SUMB[5][3] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r179/CARRYB[6][1] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r179/SUMB[7][1] ) );
  XOR21 U367 ( .A(\u_decoder/fir_filter/dp_cluster_0/r167/SUMB[5][3] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[6][1] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r167/SUMB[7][1] ) );
  XOR21 U368 ( .A(\u_decoder/fir_filter/dp_cluster_0/r180/SUMB[5][3] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[6][1] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r180/SUMB[7][1] ) );
  XOR21 U369 ( .A(n30), .B(
        \u_decoder/fir_filter/dp_cluster_0/r164/CARRYB[6][2] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r164/SUMB[7][2] ) );
  XOR21 U370 ( .A(n31), .B(
        \u_decoder/fir_filter/dp_cluster_0/r177/CARRYB[6][2] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r177/SUMB[7][2] ) );
  AOI2111 U371 ( .A(n2506), .B(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[7][5] ), .C(n1823), 
        .D(n2507), .Q(n2505) );
  INV3 U372 ( .A(n2511), .Q(n1823) );
  NOR40 U373 ( .A(n2508), .B(n2499), .C(n2509), .D(n2510), .Q(n2507) );
  AOI2111 U374 ( .A(n2419), .B(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[7][5] ), .C(n1894), 
        .D(n2420), .Q(n2418) );
  INV3 U375 ( .A(n2424), .Q(n1894) );
  NOR40 U376 ( .A(n2421), .B(n2412), .C(n2422), .D(n2423), .Q(n2420) );
  XNR31 U377 ( .A(\u_decoder/fir_filter/dp_cluster_0/r167/A2[11] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[7][5] ), .C(n2492), .Q(
        n336) );
  XNR31 U378 ( .A(\u_decoder/fir_filter/dp_cluster_0/r180/A2[11] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[7][5] ), .C(n2405), .Q(
        n337) );
  XOR21 U379 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_276/SUMB[7][2] ), 
        .B(\u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[7][1] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/A1[7] ) );
  XOR21 U380 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_308/SUMB[7][2] ), 
        .B(\u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[7][1] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/A1[7] ) );
  INV3 U381 ( .A(\u_decoder/fir_filter/dp_cluster_0/r166/CARRYB[7][3] ), .Q(
        n1808) );
  INV3 U382 ( .A(n2465), .Q(n1809) );
  INV3 U383 ( .A(\u_decoder/fir_filter/dp_cluster_0/r179/CARRYB[7][3] ), .Q(
        n1879) );
  INV3 U384 ( .A(n2378), .Q(n1880) );
  NOR21 U385 ( .A(n350), .B(n320), .Q(n2482) );
  NOR21 U386 ( .A(n351), .B(n321), .Q(n2395) );
  NOR21 U387 ( .A(n352), .B(n338), .Q(n2504) );
  NOR21 U388 ( .A(n353), .B(n339), .Q(n2417) );
  NOR21 U389 ( .A(n607), .B(n608), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r164/A2[7] ) );
  INV3 U390 ( .A(\u_decoder/fir_filter/dp_cluster_0/r164/CARRYB[7][0] ), .Q(
        n607) );
  INV3 U391 ( .A(\u_decoder/fir_filter/dp_cluster_0/r164/SUMB[7][1] ), .Q(n608) );
  NOR21 U392 ( .A(n669), .B(n670), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r177/A2[7] ) );
  INV3 U393 ( .A(\u_decoder/fir_filter/dp_cluster_0/r177/CARRYB[7][0] ), .Q(
        n669) );
  INV3 U394 ( .A(\u_decoder/fir_filter/dp_cluster_0/r177/SUMB[7][1] ), .Q(n670) );
  NOR21 U395 ( .A(\u_decoder/fir_filter/dp_cluster_0/r165/A2[6] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r165/A1[6] ), .Q(n2456) );
  NOR21 U396 ( .A(\u_decoder/fir_filter/dp_cluster_0/r178/A2[6] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r178/A1[6] ), .Q(n2369) );
  NOR21 U397 ( .A(n565), .B(n566), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[7][0] ) );
  INV3 U398 ( .A(\u_decoder/fir_filter/dp_cluster_0/r167/SUMB[6][1] ), .Q(n565) );
  INV3 U399 ( .A(\u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[6][0] ), .Q(
        n566) );
  NOR21 U400 ( .A(n627), .B(n628), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[7][0] ) );
  INV3 U401 ( .A(\u_decoder/fir_filter/dp_cluster_0/r180/SUMB[6][1] ), .Q(n627) );
  INV3 U402 ( .A(\u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[6][0] ), .Q(
        n628) );
  NOR21 U403 ( .A(n603), .B(n604), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r164/CARRYB[7][0] ) );
  INV3 U404 ( .A(\u_decoder/fir_filter/dp_cluster_0/r164/SUMB[5][2] ), .Q(n603) );
  INV3 U405 ( .A(\u_decoder/fir_filter/dp_cluster_0/r164/CARRYB[6][0] ), .Q(
        n604) );
  NOR21 U406 ( .A(n665), .B(n666), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r177/CARRYB[7][0] ) );
  INV3 U407 ( .A(\u_decoder/fir_filter/dp_cluster_0/r177/SUMB[5][2] ), .Q(n665) );
  INV3 U408 ( .A(\u_decoder/fir_filter/dp_cluster_0/r177/CARRYB[6][0] ), .Q(
        n666) );
  NAND22 U409 ( .A(\u_decoder/fir_filter/I_data_mult_1_15 ), .B(n837), .Q(
        \u_decoder/fir_filter/n1033 ) );
  XOR21 U410 ( .A(n2458), .B(
        \u_decoder/fir_filter/dp_cluster_0/r165/CARRYB[7][4] ), .Q(
        \u_decoder/fir_filter/I_data_mult_1_15 ) );
  AOI211 U411 ( .A(n2459), .B(n1868), .C(n1800), .Q(n2458) );
  INV3 U412 ( .A(n2460), .Q(n1800) );
  NAND22 U413 ( .A(\u_decoder/fir_filter/I_data_mult_0_15 ), .B(n837), .Q(
        \u_decoder/fir_filter/n1019 ) );
  XOR21 U414 ( .A(n2443), .B(
        \u_decoder/fir_filter/dp_cluster_0/r164/CARRYB[7][3] ), .Q(
        \u_decoder/fir_filter/I_data_mult_0_15 ) );
  AOI211 U415 ( .A(n2431), .B(n1868), .C(n1852), .Q(n2443) );
  INV3 U416 ( .A(n2444), .Q(n1852) );
  NAND22 U417 ( .A(\u_decoder/fir_filter/Q_data_mult_1_15 ), .B(n837), .Q(
        \u_decoder/fir_filter/n736 ) );
  XOR21 U418 ( .A(n2371), .B(
        \u_decoder/fir_filter/dp_cluster_0/r178/CARRYB[7][4] ), .Q(
        \u_decoder/fir_filter/Q_data_mult_1_15 ) );
  AOI211 U419 ( .A(n2372), .B(n1939), .C(n1871), .Q(n2371) );
  INV3 U420 ( .A(n2373), .Q(n1871) );
  NAND22 U421 ( .A(\u_decoder/fir_filter/Q_data_mult_0_15 ), .B(n837), .Q(
        \u_decoder/fir_filter/n722 ) );
  XOR21 U422 ( .A(n2356), .B(
        \u_decoder/fir_filter/dp_cluster_0/r177/CARRYB[7][3] ), .Q(
        \u_decoder/fir_filter/Q_data_mult_0_15 ) );
  AOI211 U423 ( .A(n2344), .B(n1939), .C(n1923), .Q(n2356) );
  INV3 U424 ( .A(n2357), .Q(n1923) );
  INV3 U425 ( .A(\u_decoder/fir_filter/dp_cluster_0/r165/A1[5] ), .Q(n1806) );
  INV3 U426 ( .A(\u_decoder/fir_filter/dp_cluster_0/r178/A1[5] ), .Q(n1877) );
  INV3 U427 ( .A(n2473), .Q(n1814) );
  NAND22 U428 ( .A(\u_decoder/fir_filter/dp_cluster_0/r166/A2[6] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r166/A1[6] ), .Q(n2473) );
  INV3 U429 ( .A(n2386), .Q(n1885) );
  NAND22 U430 ( .A(\u_decoder/fir_filter/dp_cluster_0/r179/A2[6] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r179/A1[6] ), .Q(n2386) );
  XNR21 U431 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_276/SUMB[7][1] ), 
        .B(\u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[7][0] ), .Q(n338) );
  XNR21 U432 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_308/SUMB[7][1] ), 
        .B(\u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[7][0] ), .Q(n339) );
  XOR21 U433 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_276/SUMB[7][5] ), 
        .B(\u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[7][4] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/A1[10] ) );
  XOR21 U434 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_308/SUMB[7][5] ), 
        .B(\u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[7][4] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/A1[10] ) );
  XOR21 U435 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_276/SUMB[4][3] ), 
        .B(\u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[6][0] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/SUMB[7][0] ) );
  XOR21 U436 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_308/SUMB[4][3] ), 
        .B(\u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[6][0] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/SUMB[7][0] ) );
  XOR21 U437 ( .A(\u_decoder/fir_filter/dp_cluster_0/r164/SUMB[5][2] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r164/CARRYB[6][0] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r164/SUMB[7][0] ) );
  XOR21 U438 ( .A(\u_decoder/fir_filter/dp_cluster_0/r177/SUMB[5][2] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r177/CARRYB[6][0] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r177/SUMB[7][0] ) );
  XOR21 U439 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_276/SUMB[5][5] ), 
        .B(\u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[6][3] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/SUMB[7][3] ) );
  XOR21 U440 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_308/SUMB[5][5] ), 
        .B(\u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[6][3] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/SUMB[7][3] ) );
  XOR21 U441 ( .A(n30), .B(
        \u_decoder/fir_filter/dp_cluster_0/r165/CARRYB[6][3] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r165/SUMB[7][3] ) );
  XOR21 U442 ( .A(n31), .B(
        \u_decoder/fir_filter/dp_cluster_0/r178/CARRYB[6][3] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r178/SUMB[7][3] ) );
  XOR21 U443 ( .A(\u_decoder/fir_filter/dp_cluster_0/r166/SUMB[7][3] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r166/CARRYB[7][2] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r166/A1[8] ) );
  XOR21 U444 ( .A(\u_decoder/fir_filter/dp_cluster_0/r165/SUMB[7][3] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r165/CARRYB[7][2] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r165/A1[8] ) );
  XOR21 U445 ( .A(\u_decoder/fir_filter/dp_cluster_0/r179/SUMB[7][3] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r179/CARRYB[7][2] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r179/A1[8] ) );
  XOR21 U446 ( .A(\u_decoder/fir_filter/dp_cluster_0/r178/SUMB[7][3] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r178/CARRYB[7][2] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r178/A1[8] ) );
  XOR21 U447 ( .A(\u_decoder/fir_filter/dp_cluster_0/r167/SUMB[7][2] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[7][1] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r167/A1[7] ) );
  XOR21 U448 ( .A(\u_decoder/fir_filter/dp_cluster_0/r180/SUMB[7][2] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[7][1] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r180/A1[7] ) );
  NOR21 U449 ( .A(n590), .B(n591), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r165/CARRYB[7][0] ) );
  INV3 U450 ( .A(\u_decoder/fir_filter/dp_cluster_0/r165/SUMB[4][3] ), .Q(n590) );
  INV3 U451 ( .A(\u_decoder/fir_filter/dp_cluster_0/r165/CARRYB[6][0] ), .Q(
        n591) );
  NOR21 U452 ( .A(n652), .B(n653), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r178/CARRYB[7][0] ) );
  INV3 U453 ( .A(\u_decoder/fir_filter/dp_cluster_0/r178/SUMB[4][3] ), .Q(n652) );
  INV3 U454 ( .A(\u_decoder/fir_filter/dp_cluster_0/r178/CARRYB[6][0] ), .Q(
        n653) );
  NOR21 U455 ( .A(n580), .B(n581), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r166/CARRYB[7][1] ) );
  INV3 U456 ( .A(\u_decoder/fir_filter/dp_cluster_0/r166/CARRYB[6][1] ), .Q(
        n581) );
  INV3 U457 ( .A(\u_decoder/fir_filter/dp_cluster_0/r166/SUMB[5][3] ), .Q(n580) );
  NOR21 U458 ( .A(n642), .B(n643), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r179/CARRYB[7][1] ) );
  INV3 U459 ( .A(\u_decoder/fir_filter/dp_cluster_0/r179/CARRYB[6][1] ), .Q(
        n643) );
  INV3 U460 ( .A(\u_decoder/fir_filter/dp_cluster_0/r179/SUMB[5][3] ), .Q(n642) );
  NOR21 U461 ( .A(n567), .B(n568), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[7][1] ) );
  INV3 U462 ( .A(\u_decoder/fir_filter/dp_cluster_0/r167/SUMB[5][3] ), .Q(n567) );
  INV3 U463 ( .A(\u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[6][1] ), .Q(
        n568) );
  NOR21 U464 ( .A(n629), .B(n630), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[7][1] ) );
  INV3 U465 ( .A(\u_decoder/fir_filter/dp_cluster_0/r180/SUMB[5][3] ), .Q(n629) );
  INV3 U466 ( .A(\u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[6][1] ), .Q(
        n630) );
  NOR21 U467 ( .A(n550), .B(n551), .Q(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[7][0] ) );
  INV3 U468 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_276/SUMB[4][3] ), .Q(
        n550) );
  INV3 U469 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[6][0] ), 
        .Q(n551) );
  NOR21 U470 ( .A(n612), .B(n613), .Q(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[7][0] ) );
  INV3 U471 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_308/SUMB[4][3] ), .Q(
        n612) );
  INV3 U472 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[6][0] ), 
        .Q(n613) );
  NOR21 U473 ( .A(n561), .B(n562), .Q(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/A2[10] ) );
  INV3 U474 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[7][3] ), 
        .Q(n561) );
  INV3 U475 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_276/SUMB[7][4] ), .Q(
        n562) );
  NOR21 U476 ( .A(n623), .B(n624), .Q(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/A2[10] ) );
  INV3 U477 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[7][3] ), 
        .Q(n623) );
  INV3 U478 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_308/SUMB[7][4] ), .Q(
        n624) );
  XNR21 U479 ( .A(\u_decoder/iq_demod/dp_cluster_1/mult_149/A1[2] ), .B(n1955), 
        .Q(\u_decoder/iq_demod/dp_cluster_1/mult_I_sin_out [4]) );
  XNR21 U480 ( .A(\u_decoder/iq_demod/dp_cluster_1/mult_150/A1[2] ), .B(n1945), 
        .Q(\u_decoder/iq_demod/dp_cluster_1/mult_Q_cos_out [4]) );
  INV3 U481 ( .A(\u_decoder/fir_filter/dp_cluster_0/r164/A2[6] ), .Q(n1857) );
  INV3 U482 ( .A(\u_decoder/fir_filter/dp_cluster_0/r177/A2[6] ), .Q(n1928) );
  NOR21 U483 ( .A(n555), .B(n556), .Q(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/A2[7] ) );
  INV3 U484 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[7][0] ), 
        .Q(n555) );
  INV3 U485 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_276/SUMB[7][1] ), .Q(
        n556) );
  NOR21 U486 ( .A(n617), .B(n618), .Q(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/A2[7] ) );
  INV3 U487 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[7][0] ), 
        .Q(n617) );
  INV3 U488 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_308/SUMB[7][1] ), .Q(
        n618) );
  XNR31 U489 ( .A(\u_decoder/fir_filter/dp_cluster_0/r166/A2[9] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r166/CARRYB[7][3] ), .C(n2465), .Q(
        n340) );
  XNR31 U490 ( .A(\u_decoder/fir_filter/dp_cluster_0/r179/A2[9] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r179/CARRYB[7][3] ), .C(n2378), .Q(
        n341) );
  NOR21 U491 ( .A(n586), .B(n587), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r166/A2[8] ) );
  INV3 U492 ( .A(\u_decoder/fir_filter/dp_cluster_0/r166/CARRYB[7][1] ), .Q(
        n586) );
  INV3 U493 ( .A(\u_decoder/fir_filter/dp_cluster_0/r166/SUMB[7][2] ), .Q(n587) );
  NOR21 U494 ( .A(n648), .B(n649), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r179/A2[8] ) );
  INV3 U495 ( .A(\u_decoder/fir_filter/dp_cluster_0/r179/CARRYB[7][1] ), .Q(
        n648) );
  INV3 U496 ( .A(\u_decoder/fir_filter/dp_cluster_0/r179/SUMB[7][2] ), .Q(n649) );
  NOR21 U497 ( .A(n595), .B(n596), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r165/A2[7] ) );
  INV3 U498 ( .A(\u_decoder/fir_filter/dp_cluster_0/r165/CARRYB[7][0] ), .Q(
        n595) );
  INV3 U499 ( .A(\u_decoder/fir_filter/dp_cluster_0/r165/SUMB[7][1] ), .Q(n596) );
  NOR21 U500 ( .A(n657), .B(n658), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r178/A2[7] ) );
  INV3 U501 ( .A(\u_decoder/fir_filter/dp_cluster_0/r178/CARRYB[7][0] ), .Q(
        n657) );
  INV3 U502 ( .A(\u_decoder/fir_filter/dp_cluster_0/r178/SUMB[7][1] ), .Q(n658) );
  NOR21 U503 ( .A(n584), .B(n585), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r166/A2[7] ) );
  INV3 U504 ( .A(\u_decoder/fir_filter/dp_cluster_0/r166/CARRYB[7][0] ), .Q(
        n584) );
  INV3 U505 ( .A(\u_decoder/fir_filter/dp_cluster_0/r166/SUMB[7][1] ), .Q(n585) );
  NOR21 U506 ( .A(n646), .B(n647), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r179/A2[7] ) );
  INV3 U507 ( .A(\u_decoder/fir_filter/dp_cluster_0/r179/CARRYB[7][0] ), .Q(
        n646) );
  INV3 U508 ( .A(\u_decoder/fir_filter/dp_cluster_0/r179/SUMB[7][1] ), .Q(n647) );
  NOR21 U509 ( .A(n557), .B(n558), .Q(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/A2[8] ) );
  INV3 U510 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[7][1] ), 
        .Q(n557) );
  INV3 U511 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_276/SUMB[7][2] ), .Q(
        n558) );
  NOR21 U512 ( .A(n619), .B(n620), .Q(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/A2[8] ) );
  INV3 U513 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[7][1] ), 
        .Q(n619) );
  INV3 U514 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_308/SUMB[7][2] ), .Q(
        n620) );
  NOR21 U515 ( .A(n597), .B(n598), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r165/A2[8] ) );
  INV3 U516 ( .A(\u_decoder/fir_filter/dp_cluster_0/r165/CARRYB[7][1] ), .Q(
        n597) );
  INV3 U517 ( .A(\u_decoder/fir_filter/dp_cluster_0/r165/SUMB[7][2] ), .Q(n598) );
  NOR21 U518 ( .A(n659), .B(n660), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r178/A2[8] ) );
  INV3 U519 ( .A(\u_decoder/fir_filter/dp_cluster_0/r178/CARRYB[7][1] ), .Q(
        n659) );
  INV3 U520 ( .A(\u_decoder/fir_filter/dp_cluster_0/r178/SUMB[7][2] ), .Q(n660) );
  NAND31 U521 ( .A(\u_decoder/fir_filter/dp_cluster_0/r164/A1[4] ), .B(n1858), 
        .C(\u_decoder/fir_filter/dp_cluster_0/r164/A1[5] ), .Q(n2435) );
  NAND31 U522 ( .A(\u_decoder/fir_filter/dp_cluster_0/r177/A1[4] ), .B(n1929), 
        .C(\u_decoder/fir_filter/dp_cluster_0/r177/A1[5] ), .Q(n2348) );
  OAI311 U523 ( .A(n1949), .B(n2340), .C(n1948), .D(n2341), .Q(n2338) );
  NAND22 U524 ( .A(\u_decoder/iq_demod/dp_cluster_0/mult_151/A2[3] ), .B(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/A1[3] ), .Q(n2341) );
  INV3 U525 ( .A(\u_decoder/iq_demod/dp_cluster_0/mult_151/A1[2] ), .Q(n1948)
         );
  OAI311 U526 ( .A(n1945), .B(n2326), .C(n1944), .D(n2327), .Q(n2324) );
  NAND22 U527 ( .A(\u_decoder/iq_demod/dp_cluster_1/mult_150/A2[3] ), .B(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/A1[3] ), .Q(n2327) );
  INV3 U528 ( .A(\u_decoder/iq_demod/dp_cluster_1/mult_150/A1[2] ), .Q(n1944)
         );
  OAI311 U529 ( .A(n1955), .B(n2319), .C(n1954), .D(n2320), .Q(n2317) );
  NAND22 U530 ( .A(\u_decoder/iq_demod/dp_cluster_1/mult_149/A2[3] ), .B(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/A1[3] ), .Q(n2320) );
  INV3 U531 ( .A(\u_decoder/iq_demod/dp_cluster_1/mult_149/A1[2] ), .Q(n1954)
         );
  OAI311 U532 ( .A(n1958), .B(n2333), .C(n1957), .D(n2334), .Q(n2331) );
  NAND22 U533 ( .A(\u_decoder/iq_demod/dp_cluster_0/mult_148/A2[3] ), .B(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/A1[3] ), .Q(n2334) );
  INV3 U534 ( .A(\u_decoder/iq_demod/dp_cluster_0/mult_148/A1[2] ), .Q(n1957)
         );
  XOR21 U535 ( .A(\u_decoder/fir_filter/dp_cluster_0/r165/SUMB[7][4] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r165/CARRYB[7][3] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r165/A1[9] ) );
  XOR21 U536 ( .A(\u_decoder/fir_filter/dp_cluster_0/r164/SUMB[7][3] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r164/CARRYB[7][2] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r164/A1[8] ) );
  XOR21 U537 ( .A(\u_decoder/fir_filter/dp_cluster_0/r178/SUMB[7][4] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r178/CARRYB[7][3] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r178/A1[9] ) );
  XOR21 U538 ( .A(\u_decoder/fir_filter/dp_cluster_0/r177/SUMB[7][3] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r177/CARRYB[7][2] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r177/A1[8] ) );
  XNR31 U539 ( .A(\u_decoder/iq_demod/dp_cluster_0/mult_151/A2[5] ), .B(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/CARRYB[3][3] ), .C(n2337), 
        .Q(n342) );
  NAND22 U540 ( .A(\u_decoder/fir_filter/dp_cluster_0/r165/PROD1[5] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r165/A1[4] ), .Q(n2455) );
  NAND22 U541 ( .A(\u_decoder/fir_filter/dp_cluster_0/r178/PROD1[5] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r178/A1[4] ), .Q(n2368) );
  NOR21 U542 ( .A(n572), .B(n573), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r167/A2[8] ) );
  INV3 U543 ( .A(\u_decoder/fir_filter/dp_cluster_0/r167/SUMB[7][2] ), .Q(n573) );
  INV3 U544 ( .A(\u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[7][1] ), .Q(
        n572) );
  NOR21 U545 ( .A(n634), .B(n635), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r180/A2[8] ) );
  INV3 U546 ( .A(\u_decoder/fir_filter/dp_cluster_0/r180/SUMB[7][2] ), .Q(n635) );
  INV3 U547 ( .A(\u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[7][1] ), .Q(
        n634) );
  NAND22 U548 ( .A(\u_decoder/fir_filter/dp_cluster_0/r164/A2[6] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r164/A1[6] ), .Q(n2436) );
  NAND22 U549 ( .A(\u_decoder/fir_filter/dp_cluster_0/r177/A2[6] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r177/A1[6] ), .Q(n2349) );
  AOI211 U550 ( .A(\u_decoder/iq_demod/dp_cluster_0/mult_151/A2[3] ), .B(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/A1[3] ), .C(n2340), .Q(n2343) );
  AOI211 U551 ( .A(\u_decoder/iq_demod/dp_cluster_1/mult_150/A2[3] ), .B(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/A1[3] ), .C(n2326), .Q(n2329) );
  AOI211 U552 ( .A(\u_decoder/iq_demod/dp_cluster_1/mult_149/A2[3] ), .B(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/A1[3] ), .C(n2319), .Q(n2322) );
  AOI211 U553 ( .A(\u_decoder/iq_demod/dp_cluster_0/mult_148/A2[3] ), .B(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/A1[3] ), .C(n2333), .Q(n2336) );
  NOR21 U554 ( .A(\u_decoder/fir_filter/dp_cluster_0/r164/A1[6] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r164/A2[6] ), .Q(n2434) );
  NOR21 U555 ( .A(\u_decoder/fir_filter/dp_cluster_0/r177/A1[6] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r177/A2[6] ), .Q(n2347) );
  AOI211 U556 ( .A(n2338), .B(\u_decoder/iq_demod/dp_cluster_0/mult_151/A1[4] ), .C(n1947), .Q(n2337) );
  INV3 U557 ( .A(n2339), .Q(n1947) );
  AOI211 U558 ( .A(n2317), .B(\u_decoder/iq_demod/dp_cluster_1/mult_149/A1[4] ), .C(n1953), .Q(n2316) );
  INV3 U559 ( .A(n2318), .Q(n1953) );
  AOI211 U560 ( .A(n2331), .B(\u_decoder/iq_demod/dp_cluster_0/mult_148/A1[4] ), .C(n1956), .Q(n2330) );
  INV3 U561 ( .A(n2332), .Q(n1956) );
  INV3 U562 ( .A(\u_decoder/iq_demod/dp_cluster_1/mult_150/CARRYB[3][3] ), .Q(
        n1952) );
  NOR21 U563 ( .A(n702), .B(n703), .Q(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/A2[5] ) );
  AOI211 U564 ( .A(n2324), .B(\u_decoder/iq_demod/dp_cluster_1/mult_150/A1[4] ), .C(n1943), .Q(n2323) );
  NOR21 U565 ( .A(\u_decoder/iq_demod/dp_cluster_0/mult_151/A2[3] ), .B(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/A1[3] ), .Q(n2340) );
  NOR21 U566 ( .A(\u_decoder/iq_demod/dp_cluster_1/mult_150/A2[3] ), .B(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/A1[3] ), .Q(n2326) );
  NOR21 U567 ( .A(\u_decoder/iq_demod/dp_cluster_1/mult_149/A2[3] ), .B(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/A1[3] ), .Q(n2319) );
  NOR21 U568 ( .A(\u_decoder/iq_demod/dp_cluster_0/mult_148/A2[3] ), .B(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/A1[3] ), .Q(n2333) );
  NOR21 U569 ( .A(n552), .B(n553), .Q(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[7][3] ) );
  INV3 U570 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[6][3] ), 
        .Q(n553) );
  INV3 U571 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_276/SUMB[5][5] ), .Q(
        n552) );
  NOR21 U572 ( .A(n614), .B(n615), .Q(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[7][3] ) );
  INV3 U573 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[6][3] ), 
        .Q(n615) );
  INV3 U574 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_308/SUMB[5][5] ), .Q(
        n614) );
  NOR21 U575 ( .A(n559), .B(n560), .Q(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/A2[9] ) );
  INV3 U576 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[7][2] ), 
        .Q(n559) );
  INV3 U577 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_276/SUMB[7][3] ), .Q(
        n560) );
  NOR21 U578 ( .A(n621), .B(n622), .Q(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/A2[9] ) );
  INV3 U579 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[7][2] ), 
        .Q(n621) );
  INV3 U580 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_308/SUMB[7][3] ), .Q(
        n622) );
  XNR31 U581 ( .A(\u_decoder/iq_demod/dp_cluster_0/mult_151/A2[4] ), .B(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/A1[4] ), .C(n2338), .Q(n343)
         );
  XNR21 U582 ( .A(n2335), .B(n2336), .Q(
        \u_decoder/iq_demod/dp_cluster_0/mult_I_cos_out [5]) );
  XNR21 U583 ( .A(\u_decoder/iq_demod/dp_cluster_0/mult_148/A1[2] ), .B(n1958), 
        .Q(\u_decoder/iq_demod/dp_cluster_0/mult_I_cos_out [4]) );
  NOR21 U584 ( .A(n563), .B(n564), .Q(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/A2[11] ) );
  INV3 U585 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[7][4] ), 
        .Q(n563) );
  INV3 U586 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_276/SUMB[7][5] ), .Q(
        n564) );
  NOR21 U587 ( .A(n625), .B(n626), .Q(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/A2[11] ) );
  INV3 U588 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[7][4] ), 
        .Q(n625) );
  INV3 U589 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_308/SUMB[7][5] ), .Q(
        n626) );
  NOR21 U590 ( .A(n609), .B(n610), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r164/A2[8] ) );
  INV3 U591 ( .A(\u_decoder/fir_filter/dp_cluster_0/r164/CARRYB[7][1] ), .Q(
        n609) );
  INV3 U592 ( .A(\u_decoder/fir_filter/dp_cluster_0/r164/SUMB[7][2] ), .Q(n610) );
  NOR21 U593 ( .A(n671), .B(n672), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r177/A2[8] ) );
  INV3 U594 ( .A(\u_decoder/fir_filter/dp_cluster_0/r177/CARRYB[7][1] ), .Q(
        n671) );
  INV3 U595 ( .A(\u_decoder/fir_filter/dp_cluster_0/r177/SUMB[7][2] ), .Q(n672) );
  INV3 U596 ( .A(\u_decoder/fir_filter/I_data_mult_0 [8]), .Q(n1854) );
  IMUX21 U597 ( .A(n1856), .B(n2439), .S(n2435), .Q(n2438) );
  XNR21 U598 ( .A(n1855), .B(n2435), .Q(n2437) );
  INV3 U599 ( .A(\u_decoder/fir_filter/Q_data_mult_0 [8]), .Q(n1925) );
  IMUX21 U600 ( .A(n1927), .B(n2352), .S(n2348), .Q(n2351) );
  XNR21 U601 ( .A(n1926), .B(n2348), .Q(n2350) );
  NOR21 U602 ( .A(\u_decoder/I_prefilter [5]), .B(n592), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r165/CARRYB[7][3] ) );
  INV3 U603 ( .A(\u_decoder/fir_filter/dp_cluster_0/r165/CARRYB[6][3] ), .Q(
        n592) );
  NOR21 U604 ( .A(\u_decoder/I_prefilter [5]), .B(n605), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r164/CARRYB[7][2] ) );
  INV3 U605 ( .A(\u_decoder/fir_filter/dp_cluster_0/r164/CARRYB[6][2] ), .Q(
        n605) );
  NOR21 U606 ( .A(\u_decoder/Q_prefilter [5]), .B(n654), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r178/CARRYB[7][3] ) );
  INV3 U607 ( .A(\u_decoder/fir_filter/dp_cluster_0/r178/CARRYB[6][3] ), .Q(
        n654) );
  NOR21 U608 ( .A(\u_decoder/Q_prefilter [5]), .B(n667), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r177/CARRYB[7][2] ) );
  INV3 U609 ( .A(\u_decoder/fir_filter/dp_cluster_0/r177/CARRYB[6][2] ), .Q(
        n667) );
  INV3 U610 ( .A(\u_decoder/iq_demod/dp_cluster_1/mult_150/ab[0][2] ), .Q(n706) );
  INV3 U611 ( .A(\u_decoder/iq_demod/dp_cluster_1/mult_150/ab[0][1] ), .Q(n704) );
  INV3 U612 ( .A(\u_decoder/iq_demod/dp_cluster_0/mult_148/ab[0][2] ), .Q(n694) );
  INV3 U613 ( .A(\u_decoder/iq_demod/dp_cluster_0/mult_148/ab[0][1] ), .Q(n692) );
  INV3 U614 ( .A(\u_decoder/iq_demod/dp_cluster_0/mult_151/ab[0][2] ), .Q(n682) );
  INV3 U615 ( .A(\u_decoder/iq_demod/dp_cluster_0/mult_151/ab[0][1] ), .Q(n680) );
  INV3 U616 ( .A(\u_decoder/iq_demod/dp_cluster_1/mult_149/ab[0][2] ), .Q(n718) );
  INV3 U617 ( .A(\u_decoder/iq_demod/dp_cluster_1/mult_149/ab[0][1] ), .Q(n716) );
  INV3 U618 ( .A(\u_decoder/iq_demod/dp_cluster_0/mult_151/ab[1][0] ), .Q(n681) );
  INV3 U619 ( .A(\u_decoder/iq_demod/dp_cluster_1/mult_150/ab[1][1] ), .Q(n707) );
  INV3 U620 ( .A(\u_decoder/iq_demod/dp_cluster_1/mult_149/ab[1][0] ), .Q(n717) );
  INV3 U621 ( .A(\u_decoder/iq_demod/dp_cluster_0/mult_148/ab[1][1] ), .Q(n695) );
  INV3 U622 ( .A(\u_decoder/iq_demod/dp_cluster_1/mult_150/ab[1][2] ), .Q(n709) );
  INV3 U623 ( .A(\u_decoder/iq_demod/dp_cluster_0/mult_148/ab[1][2] ), .Q(n697) );
  INV3 U624 ( .A(\u_decoder/iq_demod/dp_cluster_1/mult_150/ab[1][0] ), .Q(n705) );
  INV3 U625 ( .A(\u_decoder/iq_demod/dp_cluster_0/mult_148/ab[1][0] ), .Q(n693) );
  INV3 U626 ( .A(\u_decoder/iq_demod/dp_cluster_0/mult_151/ab[1][1] ), .Q(n683) );
  INV3 U627 ( .A(\u_decoder/iq_demod/dp_cluster_1/mult_149/ab[1][1] ), .Q(n719) );
  INV3 U628 ( .A(\u_decoder/iq_demod/dp_cluster_0/mult_151/ab[1][2] ), .Q(n685) );
  INV3 U629 ( .A(\u_decoder/iq_demod/dp_cluster_1/mult_149/ab[1][2] ), .Q(n721) );
  INV3 U630 ( .A(n2325), .Q(n1943) );
  INV3 U631 ( .A(n2489), .Q(n1840) );
  INV3 U632 ( .A(n2402), .Q(n1911) );
  OAI2111 U633 ( .A(n1125), .B(n1045), .C(n1042), .D(n1090), .Q(
        \u_cdr/phd1/cnt_phd/N12 ) );
  XOR21 U634 ( .A(\u_decoder/fir_filter/dp_cluster_0/r167/SUMB[7][4] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[7][3] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r167/A1[9] ) );
  XOR21 U635 ( .A(\u_decoder/fir_filter/dp_cluster_0/r180/SUMB[7][4] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[7][3] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r180/A1[9] ) );
  NAND31 U636 ( .A(n1125), .B(n1124), .C(n1045), .Q(n1042) );
  NAND22 U637 ( .A(\u_decoder/fir_filter/dp_cluster_0/r164/PROD1[4] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r164/A1[3] ), .Q(n2441) );
  NAND22 U638 ( .A(\u_decoder/fir_filter/dp_cluster_0/r177/PROD1[4] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r177/A1[3] ), .Q(n2354) );
  NAND22 U639 ( .A(n977), .B(n1660), .Q(\u_coder/n274 ) );
  NOR21 U640 ( .A(n576), .B(n577), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r167/A2[10] ) );
  INV3 U641 ( .A(\u_decoder/fir_filter/dp_cluster_0/r167/SUMB[7][4] ), .Q(n577) );
  INV3 U642 ( .A(\u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[7][3] ), .Q(
        n576) );
  NOR21 U643 ( .A(n638), .B(n639), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r180/A2[10] ) );
  INV3 U644 ( .A(\u_decoder/fir_filter/dp_cluster_0/r180/SUMB[7][4] ), .Q(n639) );
  INV3 U645 ( .A(\u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[7][3] ), .Q(
        n638) );
  NOR21 U646 ( .A(n574), .B(n575), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r167/A2[9] ) );
  INV3 U647 ( .A(\u_decoder/fir_filter/dp_cluster_0/r167/SUMB[7][3] ), .Q(n575) );
  INV3 U648 ( .A(\u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[7][2] ), .Q(
        n574) );
  NOR21 U649 ( .A(n636), .B(n637), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r180/A2[9] ) );
  INV3 U650 ( .A(\u_decoder/fir_filter/dp_cluster_0/r180/SUMB[7][3] ), .Q(n637) );
  INV3 U651 ( .A(\u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[7][2] ), .Q(
        n636) );
  NOR21 U652 ( .A(n722), .B(n723), .Q(
        \u_decoder/iq_demod/dp_cluster_1/add_154/carry [1]) );
  XOR21 U653 ( .A(\u_decoder/iq_demod/dp_cluster_1/mult_149/ab[0][1] ), .B(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/ab[1][0] ), .Q(
        \u_decoder/iq_demod/dp_cluster_1/mult_I_sin_out [1]) );
  XOR21 U654 ( .A(\u_decoder/iq_demod/dp_cluster_1/mult_150/ab[0][1] ), .B(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/ab[1][0] ), .Q(
        \u_decoder/iq_demod/dp_cluster_1/mult_Q_cos_out [1]) );
  INV3 U655 ( .A(\u_decoder/iq_demod/dp_cluster_0/mult_Q_sin_out [2]), .Q(
        n1951) );
  INV3 U656 ( .A(n470), .Q(\u_decoder/iq_demod/dp_cluster_0/sub_153/carry [1])
         );
  XOR21 U657 ( .A(\u_decoder/iq_demod/dp_cluster_0/mult_148/ab[0][1] ), .B(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/ab[1][0] ), .Q(
        \u_decoder/iq_demod/dp_cluster_0/mult_I_cos_out [1]) );
  BUF2 U658 ( .A(n812), .Q(n813) );
  AOI211 U659 ( .A(n1724), .B(n1716), .C(\u_coder/n274 ), .Q(n812) );
  INV3 U660 ( .A(\u_decoder/fir_filter/I_data_mult_2[8] ), .Q(n1813) );
  AOI211 U661 ( .A(\u_decoder/fir_filter/dp_cluster_0/r166/A1[6] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r166/A2[6] ), .C(n2467), .Q(
        \u_decoder/fir_filter/I_data_mult_2[8] ) );
  NOR21 U662 ( .A(\u_decoder/fir_filter/dp_cluster_0/r166/A2[6] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r166/A1[6] ), .Q(n2467) );
  INV3 U663 ( .A(\u_decoder/fir_filter/Q_data_mult_2[8] ), .Q(n1884) );
  AOI211 U664 ( .A(\u_decoder/fir_filter/dp_cluster_0/r179/A1[6] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r179/A2[6] ), .C(n2380), .Q(
        \u_decoder/fir_filter/Q_data_mult_2[8] ) );
  NOR21 U665 ( .A(\u_decoder/fir_filter/dp_cluster_0/r179/A2[6] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r179/A1[6] ), .Q(n2380) );
  NOR21 U666 ( .A(n611), .B(n602), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r164/A2[9] ) );
  INV3 U667 ( .A(\u_decoder/fir_filter/dp_cluster_0/r164/CARRYB[7][2] ), .Q(
        n611) );
  NOR21 U668 ( .A(n673), .B(n664), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r177/A2[9] ) );
  INV3 U669 ( .A(\u_decoder/fir_filter/dp_cluster_0/r177/CARRYB[7][2] ), .Q(
        n673) );
  NOR21 U670 ( .A(n599), .B(n600), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r165/A2[9] ) );
  INV3 U671 ( .A(\u_decoder/fir_filter/dp_cluster_0/r165/CARRYB[7][2] ), .Q(
        n599) );
  INV3 U672 ( .A(\u_decoder/fir_filter/dp_cluster_0/r165/SUMB[7][3] ), .Q(n600) );
  NOR21 U673 ( .A(n661), .B(n662), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r178/A2[9] ) );
  INV3 U674 ( .A(\u_decoder/fir_filter/dp_cluster_0/r178/CARRYB[7][2] ), .Q(
        n661) );
  INV3 U675 ( .A(\u_decoder/fir_filter/dp_cluster_0/r178/SUMB[7][3] ), .Q(n662) );
  NOR21 U676 ( .A(n588), .B(n589), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r166/A2[9] ) );
  INV3 U677 ( .A(\u_decoder/fir_filter/dp_cluster_0/r166/CARRYB[7][2] ), .Q(
        n588) );
  INV3 U678 ( .A(\u_decoder/fir_filter/dp_cluster_0/r166/SUMB[7][3] ), .Q(n589) );
  NOR21 U679 ( .A(n650), .B(n651), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r179/A2[9] ) );
  INV3 U680 ( .A(\u_decoder/fir_filter/dp_cluster_0/r179/CARRYB[7][2] ), .Q(
        n650) );
  INV3 U681 ( .A(\u_decoder/fir_filter/dp_cluster_0/r179/SUMB[7][3] ), .Q(n651) );
  INV3 U682 ( .A(\u_decoder/fir_filter/I_data_mult_3 [8]), .Q(n1846) );
  AOI211 U683 ( .A(n350), .B(n320), .C(n2482), .Q(
        \u_decoder/fir_filter/I_data_mult_3 [8]) );
  INV3 U684 ( .A(\u_decoder/fir_filter/Q_data_mult_3 [8]), .Q(n1917) );
  AOI211 U685 ( .A(n351), .B(n321), .C(n2395), .Q(
        \u_decoder/fir_filter/Q_data_mult_3 [8]) );
  NOR21 U686 ( .A(n2455), .B(n1806), .Q(n2454) );
  AOI211 U687 ( .A(\u_decoder/fir_filter/dp_cluster_0/r165/A1[6] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r165/A2[6] ), .C(n2456), .Q(n2453)
         );
  NOR21 U688 ( .A(n2368), .B(n1877), .Q(n2367) );
  AOI211 U689 ( .A(\u_decoder/fir_filter/dp_cluster_0/r178/A1[6] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r178/A2[6] ), .C(n2369), .Q(n2366)
         );
  NAND22 U690 ( .A(n1858), .B(\u_decoder/fir_filter/dp_cluster_0/r164/A1[4] ), 
        .Q(n2440) );
  NAND22 U691 ( .A(n1929), .B(\u_decoder/fir_filter/dp_cluster_0/r177/A1[4] ), 
        .Q(n2353) );
  INV3 U692 ( .A(\u_inFIFO/N249 ), .Q(n1699) );
  INV3 U693 ( .A(\u_coder/n152 ), .Q(n1589) );
  NOR21 U694 ( .A(n1946), .B(
        \u_decoder/iq_demod/dp_cluster_0/mult_I_cos_out [0]), .Q(n470) );
  NOR21 U695 ( .A(n601), .B(n602), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r165/A2[10] ) );
  INV3 U696 ( .A(\u_decoder/fir_filter/dp_cluster_0/r165/SUMB[7][4] ), .Q(n602) );
  INV3 U697 ( .A(\u_decoder/fir_filter/dp_cluster_0/r165/CARRYB[7][3] ), .Q(
        n601) );
  NOR21 U698 ( .A(n663), .B(n664), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r178/A2[10] ) );
  INV3 U699 ( .A(\u_decoder/fir_filter/dp_cluster_0/r178/SUMB[7][4] ), .Q(n664) );
  INV3 U700 ( .A(\u_decoder/fir_filter/dp_cluster_0/r178/CARRYB[7][3] ), .Q(
        n663) );
  INV3 U701 ( .A(\u_decoder/iq_demod/dp_cluster_1/mult_Q_cos_out [0]), .Q(n722) );
  INV3 U702 ( .A(\u_decoder/iq_demod/dp_cluster_1/mult_I_sin_out [0]), .Q(n723) );
  XOR21 U703 ( .A(\u_decoder/fir_filter/dp_cluster_0/r167/SUMB[7][5] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[7][4] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r167/A1[10] ) );
  XOR21 U704 ( .A(\u_decoder/fir_filter/dp_cluster_0/r180/SUMB[7][5] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[7][4] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r180/A1[10] ) );
  NAND22 U705 ( .A(\u_coder/n188 ), .B(\u_coder/n196 ), .Q(\u_coder/n167 ) );
  NAND22 U706 ( .A(n1756), .B(n1749), .Q(\u_coder/n230 ) );
  XOR21 U707 ( .A(n2441), .B(\u_decoder/fir_filter/dp_cluster_0/r164/A1[4] ), 
        .Q(n344) );
  XOR21 U708 ( .A(n2354), .B(\u_decoder/fir_filter/dp_cluster_0/r177/A1[4] ), 
        .Q(n345) );
  XOR21 U709 ( .A(n2455), .B(\u_decoder/fir_filter/dp_cluster_0/r165/A1[5] ), 
        .Q(n346) );
  XOR21 U710 ( .A(n2368), .B(\u_decoder/fir_filter/dp_cluster_0/r178/A1[5] ), 
        .Q(n347) );
  INV3 U711 ( .A(\u_coder/n241 ), .Q(n1749) );
  INV3 U712 ( .A(\u_decoder/iq_demod/dp_cluster_0/mult_151/SUMB[3][3] ), .Q(
        n679) );
  INV3 U713 ( .A(\u_decoder/iq_demod/dp_cluster_1/mult_150/SUMB[3][3] ), .Q(
        n703) );
  INV3 U714 ( .A(\u_decoder/fir_filter/I_data_mult_3 [6]), .Q(n1847) );
  INV3 U715 ( .A(\u_decoder/fir_filter/Q_data_mult_3 [6]), .Q(n1918) );
  INV3 U716 ( .A(\u_coder/n254 ), .Q(n1473) );
  NOR21 U717 ( .A(n966), .B(n1702), .Q(\u_inFIFO/n195 ) );
  NAND22 U718 ( .A(n1724), .B(\u_coder/n196 ), .Q(\u_coder/n186 ) );
  NAND22 U719 ( .A(n977), .B(n958), .Q(\u_outFIFO/n502 ) );
  NOR21 U720 ( .A(\u_coder/n233 ), .B(\u_coder/n241 ), .Q(\u_coder/n211 ) );
  NAND22 U721 ( .A(\u_outFIFO/n511 ), .B(n969), .Q(\u_outFIFO/n544 ) );
  NAND22 U722 ( .A(n978), .B(n967), .Q(\u_inFIFO/n118 ) );
  INV3 U723 ( .A(\u_inFIFO/n119 ), .Q(n968) );
  NAND22 U724 ( .A(n978), .B(\u_coder/n186 ), .Q(\u_coder/n273 ) );
  NOR21 U725 ( .A(n578), .B(n579), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r167/A2[11] ) );
  INV3 U726 ( .A(\u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[7][4] ), .Q(
        n578) );
  INV3 U727 ( .A(\u_decoder/fir_filter/dp_cluster_0/r167/SUMB[7][5] ), .Q(n579) );
  NOR21 U728 ( .A(n640), .B(n641), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r180/A2[11] ) );
  INV3 U729 ( .A(\u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[7][4] ), .Q(
        n640) );
  INV3 U730 ( .A(\u_decoder/fir_filter/dp_cluster_0/r180/SUMB[7][5] ), .Q(n641) );
  INV3 U731 ( .A(\u_coder/n310 ), .Q(n1714) );
  INV3 U732 ( .A(\u_coder/n309 ), .Q(n1726) );
  INV3 U733 ( .A(\u_decoder/fir_filter/I_data_mult_3 [5]), .Q(n1848) );
  INV3 U734 ( .A(\u_decoder/fir_filter/I_data_mult_3 [4]), .Q(n1849) );
  INV3 U735 ( .A(\u_decoder/fir_filter/dp_cluster_0/r166/SUMB[5][1] ), .Q(
        n1815) );
  INV3 U736 ( .A(\u_decoder/fir_filter/Q_data_mult_3 [5]), .Q(n1919) );
  INV3 U737 ( .A(\u_decoder/fir_filter/Q_data_mult_3 [4]), .Q(n1920) );
  INV3 U738 ( .A(\u_decoder/fir_filter/dp_cluster_0/r179/SUMB[5][1] ), .Q(
        n1886) );
  INV3 U739 ( .A(\u_outFIFO/n215 ), .Q(n959) );
  INV3 U740 ( .A(\u_decoder/iq_demod/dp_cluster_1/mult_149/CARRYB[3][3] ), .Q(
        n1959) );
  INV3 U741 ( .A(\u_decoder/iq_demod/dp_cluster_0/mult_148/CARRYB[3][3] ), .Q(
        n1960) );
  NOR31 U742 ( .A(\u_inFIFO/n225 ), .B(n1702), .C(\u_inFIFO/n223 ), .Q(
        \u_inFIFO/n211 ) );
  NAND22 U743 ( .A(n1746), .B(n1756), .Q(n808) );
  NAND22 U744 ( .A(n1746), .B(n1756), .Q(\u_coder/n283 ) );
  NOR21 U745 ( .A(\u_outFIFO/n525 ), .B(n1466), .Q(\u_outFIFO/n520 ) );
  NAND22 U746 ( .A(n977), .B(\u_cdr/n43 ), .Q(\u_cdr/n46 ) );
  NAND22 U747 ( .A(n977), .B(n1656), .Q(\u_cdr/n23 ) );
  INV3 U748 ( .A(\u_cdr/n38 ), .Q(n1656) );
  BUF2 U749 ( .A(\u_coder/n286 ), .Q(n810) );
  BUF2 U750 ( .A(\u_coder/n286 ), .Q(n811) );
  INV3 U751 ( .A(\u_decoder/fir_filter/dp_cluster_0/r164/CARRYB[7][3] ), .Q(
        n1868) );
  INV3 U752 ( .A(\u_decoder/fir_filter/dp_cluster_0/r177/CARRYB[7][3] ), .Q(
        n1939) );
  INV3 U753 ( .A(\u_decoder/fir_filter/I_data_mult_3 [3]), .Q(n1850) );
  INV3 U754 ( .A(\u_decoder/fir_filter/dp_cluster_0/r166/SUMB[4][1] ), .Q(
        n1816) );
  INV3 U755 ( .A(\u_decoder/fir_filter/Q_data_mult_3 [3]), .Q(n1921) );
  INV3 U756 ( .A(\u_decoder/fir_filter/dp_cluster_0/r179/SUMB[4][1] ), .Q(
        n1887) );
  NAND22 U757 ( .A(n978), .B(\u_inFIFO/n209 ), .Q(\u_inFIFO/n111 ) );
  INV3 U758 ( .A(\u_inFIFO/n223 ), .Q(n1485) );
  NAND22 U759 ( .A(n977), .B(\u_inFIFO/n111 ), .Q(\u_inFIFO/n110 ) );
  NAND22 U760 ( .A(\u_decoder/iq_demod/cossin_dig/n41 ), .B(
        \u_decoder/iq_demod/cossin_dig/n40 ), .Q(
        \u_decoder/iq_demod/cossin_dig/n39 ) );
  NAND22 U761 ( .A(n976), .B(\u_decoder/iq_demod/cossin_dig/n42 ), .Q(
        \u_decoder/iq_demod/cossin_dig/n41 ) );
  INV3 U762 ( .A(\u_decoder/fir_filter/I_data_mult_3 [2]), .Q(n1851) );
  INV3 U763 ( .A(\u_decoder/fir_filter/dp_cluster_0/r166/SUMB[3][1] ), .Q(
        n1817) );
  INV3 U764 ( .A(\u_decoder/fir_filter/Q_data_mult_3 [2]), .Q(n1922) );
  INV3 U765 ( .A(\u_decoder/fir_filter/I_data_mult_1[4] ), .Q(n1807) );
  INV3 U766 ( .A(\u_decoder/fir_filter/dp_cluster_0/r179/SUMB[3][1] ), .Q(
        n1888) );
  INV3 U767 ( .A(\u_decoder/fir_filter/Q_data_mult_1[4] ), .Q(n1878) );
  INV3 U768 ( .A(\u_decoder/fir_filter/I_data_mult_0 [3]), .Q(n1859) );
  INV3 U769 ( .A(\u_decoder/fir_filter/Q_data_mult_0 [3]), .Q(n1930) );
  NAND22 U770 ( .A(n977), .B(n1468), .Q(\u_outFIFO/n533 ) );
  BUF2 U771 ( .A(\u_cordic/mycordic/n363 ), .Q(n835) );
  BUF2 U772 ( .A(\u_decoder/fir_filter/n721 ), .Q(n940) );
  BUF2 U773 ( .A(\u_decoder/fir_filter/n721 ), .Q(n939) );
  BUF2 U774 ( .A(\u_decoder/fir_filter/n721 ), .Q(n941) );
  BUF2 U775 ( .A(\u_cordic/mycordic/n363 ), .Q(n836) );
  INV3 U776 ( .A(\u_decoder/iq_demod/n69 ), .Q(n1584) );
  NOR21 U777 ( .A(n814), .B(n1758), .Q(\u_coder/N521 ) );
  INV3 U778 ( .A(\u_coder/N476 ), .Q(n1758) );
  NOR21 U779 ( .A(\u_coder/n315 ), .B(n1759), .Q(\u_coder/N520 ) );
  INV3 U780 ( .A(\u_coder/N475 ), .Q(n1759) );
  XOR21 U781 ( .A(n960), .B(
        \u_decoder/fir_filter/dp_cluster_0/r166/SUMB[6][1] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r166/SUMB[7][0] ) );
  XOR21 U782 ( .A(n962), .B(
        \u_decoder/fir_filter/dp_cluster_0/r179/SUMB[6][1] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r179/SUMB[7][0] ) );
  XOR21 U783 ( .A(n961), .B(
        \u_decoder/fir_filter/dp_cluster_0/r165/SUMB[7][0] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r165/A1[5] ) );
  XOR21 U784 ( .A(n963), .B(
        \u_decoder/fir_filter/dp_cluster_0/r178/SUMB[7][0] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r178/A1[5] ) );
  XOR21 U785 ( .A(n960), .B(
        \u_decoder/fir_filter/dp_cluster_0/r166/SUMB[6][3] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r166/SUMB[7][2] ) );
  XOR21 U786 ( .A(n962), .B(
        \u_decoder/fir_filter/dp_cluster_0/r179/SUMB[6][3] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r179/SUMB[7][2] ) );
  XOR21 U787 ( .A(n960), .B(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/SUMB[6][5] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/SUMB[7][4] ) );
  XOR21 U788 ( .A(n962), .B(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/SUMB[6][5] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/SUMB[7][4] ) );
  XOR21 U789 ( .A(n960), .B(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/SUMB[5][3] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/SUMB[7][1] ) );
  XOR21 U790 ( .A(n962), .B(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/SUMB[5][3] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/SUMB[7][1] ) );
  XOR21 U791 ( .A(n960), .B(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/SUMB[6][3] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/SUMB[7][2] ) );
  XOR21 U792 ( .A(n962), .B(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/SUMB[6][3] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/SUMB[7][2] ) );
  XOR21 U793 ( .A(n961), .B(
        \u_decoder/fir_filter/dp_cluster_0/r165/SUMB[5][3] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r165/SUMB[7][1] ) );
  XOR21 U794 ( .A(n963), .B(
        \u_decoder/fir_filter/dp_cluster_0/r178/SUMB[5][3] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r178/SUMB[7][1] ) );
  XOR21 U795 ( .A(n961), .B(
        \u_decoder/fir_filter/dp_cluster_0/r165/SUMB[6][3] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r165/SUMB[7][2] ) );
  XOR21 U796 ( .A(n963), .B(
        \u_decoder/fir_filter/dp_cluster_0/r178/SUMB[6][3] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r178/SUMB[7][2] ) );
  XOR21 U797 ( .A(n961), .B(
        \u_decoder/fir_filter/dp_cluster_0/r164/SUMB[6][2] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r164/SUMB[7][1] ) );
  XOR21 U798 ( .A(n963), .B(
        \u_decoder/fir_filter/dp_cluster_0/r177/SUMB[6][2] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r177/SUMB[7][1] ) );
  NAND22 U799 ( .A(\u_decoder/fir_filter/I_data_mult_2_15 ), .B(n837), .Q(
        \u_decoder/fir_filter/n1050 ) );
  XNR21 U800 ( .A(n961), .B(n2468), .Q(\u_decoder/fir_filter/I_data_mult_2_15 ) );
  NAND22 U801 ( .A(n2469), .B(n961), .Q(n2468) );
  NAND22 U802 ( .A(\u_decoder/fir_filter/Q_data_mult_2_15 ), .B(n837), .Q(
        \u_decoder/fir_filter/n753 ) );
  XNR21 U803 ( .A(n963), .B(n2381), .Q(\u_decoder/fir_filter/Q_data_mult_2_15 ) );
  NAND22 U804 ( .A(n2382), .B(n963), .Q(n2381) );
  NOR21 U805 ( .A(n583), .B(n229), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r166/A2[6] ) );
  INV3 U806 ( .A(\u_decoder/fir_filter/dp_cluster_0/r166/SUMB[7][0] ), .Q(n583) );
  NOR21 U807 ( .A(n645), .B(n230), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r179/A2[6] ) );
  INV3 U808 ( .A(\u_decoder/fir_filter/dp_cluster_0/r179/SUMB[7][0] ), .Q(n645) );
  XOR21 U809 ( .A(n771), .B(n773), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r167/SUMB[2][1] ) );
  XOR21 U810 ( .A(n770), .B(n51), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r165/SUMB[2][3] ) );
  XOR21 U811 ( .A(n761), .B(n763), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r180/SUMB[2][1] ) );
  XOR21 U812 ( .A(n760), .B(n52), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r178/SUMB[2][3] ) );
  XOR21 U813 ( .A(n768), .B(n773), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r167/SUMB[3][3] ) );
  XOR21 U814 ( .A(n770), .B(n51), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r164/SUMB[2][2] ) );
  XOR21 U815 ( .A(n758), .B(n763), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r180/SUMB[3][3] ) );
  XOR21 U816 ( .A(n760), .B(n52), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r177/SUMB[2][2] ) );
  NOR21 U817 ( .A(n51), .B(n59), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r166/CARRYB[1][3] ) );
  NOR21 U818 ( .A(n52), .B(n60), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r179/CARRYB[1][3] ) );
  NOR21 U819 ( .A(n59), .B(n51), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[1][0] ) );
  NOR21 U820 ( .A(n60), .B(n52), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[1][0] ) );
  NOR21 U821 ( .A(n51), .B(n59), .Q(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[1][5] ) );
  NOR21 U822 ( .A(n52), .B(n60), .Q(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[1][5] ) );
  NOR21 U823 ( .A(n53), .B(n51), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r166/CARRYB[2][1] ) );
  XOR21 U824 ( .A(n772), .B(\u_decoder/I_prefilter [1]), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r166/SUMB[1][3] ) );
  NOR21 U825 ( .A(n54), .B(n52), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r179/CARRYB[2][1] ) );
  XOR21 U826 ( .A(n762), .B(\u_decoder/Q_prefilter [1]), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r179/SUMB[1][3] ) );
  NOR21 U827 ( .A(n53), .B(n51), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[2][1] ) );
  NOR21 U828 ( .A(n54), .B(n52), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[2][1] ) );
  NOR21 U829 ( .A(n51), .B(n53), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r164/CARRYB[2][0] ) );
  NOR21 U830 ( .A(n52), .B(n54), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r177/CARRYB[2][0] ) );
  NOR21 U831 ( .A(n53), .B(n51), .Q(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[2][3] ) );
  XOR21 U832 ( .A(n772), .B(\u_decoder/I_prefilter [1]), .Q(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/SUMB[1][5] ) );
  NOR21 U833 ( .A(n54), .B(n52), .Q(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[2][3] ) );
  XOR21 U834 ( .A(n762), .B(\u_decoder/Q_prefilter [1]), .Q(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/SUMB[1][5] ) );
  NOR21 U835 ( .A(n51), .B(n69), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r165/CARRYB[3][0] ) );
  NOR21 U836 ( .A(n52), .B(n70), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r178/CARRYB[3][0] ) );
  NOR21 U837 ( .A(n53), .B(n772), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r165/CARRYB[2][3] ) );
  NOR21 U838 ( .A(n54), .B(n762), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r178/CARRYB[2][3] ) );
  NOR21 U839 ( .A(n53), .B(n773), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r164/CARRYB[2][2] ) );
  NOR21 U840 ( .A(n54), .B(n763), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r177/CARRYB[2][2] ) );
  NOR21 U841 ( .A(n741), .B(n742), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r166/CARRYB[7][0] ) );
  INV3 U842 ( .A(n960), .Q(n741) );
  INV3 U843 ( .A(\u_decoder/fir_filter/dp_cluster_0/r166/SUMB[6][1] ), .Q(n742) );
  NOR21 U844 ( .A(n730), .B(n731), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r179/CARRYB[7][0] ) );
  INV3 U845 ( .A(n962), .Q(n730) );
  INV3 U846 ( .A(\u_decoder/fir_filter/dp_cluster_0/r179/SUMB[6][1] ), .Q(n731) );
  NOR21 U847 ( .A(n735), .B(n736), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r164/CARRYB[7][1] ) );
  INV3 U848 ( .A(n961), .Q(n735) );
  INV3 U849 ( .A(\u_decoder/fir_filter/dp_cluster_0/r164/SUMB[6][2] ), .Q(n736) );
  NOR21 U850 ( .A(n724), .B(n725), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r177/CARRYB[7][1] ) );
  INV3 U851 ( .A(n963), .Q(n724) );
  INV3 U852 ( .A(\u_decoder/fir_filter/dp_cluster_0/r177/SUMB[6][2] ), .Q(n725) );
  INV3 U853 ( .A(n2555), .Q(n2091) );
  INV3 U854 ( .A(n2536), .Q(n1971) );
  INV3 U855 ( .A(n2546), .Q(n2099) );
  INV3 U856 ( .A(n2527), .Q(n1979) );
  INV3 U857 ( .A(n2483), .Q(n1839) );
  AOI2111 U858 ( .A(n2484), .B(
        \u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[7][5] ), .C(n1840), .D(
        n2485), .Q(n2483) );
  XNR21 U859 ( .A(n961), .B(n2469), .Q(n348) );
  INV3 U860 ( .A(n2396), .Q(n1910) );
  AOI2111 U861 ( .A(n2397), .B(
        \u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[7][5] ), .C(n1911), .D(
        n2398), .Q(n2396) );
  XNR21 U862 ( .A(n963), .B(n2382), .Q(n349) );
  NAND22 U863 ( .A(\u_decoder/fir_filter/dp_cluster_0/r167/SUMB[7][0] ), .B(
        n960), .Q(n350) );
  NAND22 U864 ( .A(\u_decoder/fir_filter/dp_cluster_0/r180/SUMB[7][0] ), .B(
        n962), .Q(n351) );
  NOR21 U865 ( .A(\u_coder/n315 ), .B(n1761), .Q(\u_coder/N518 ) );
  INV3 U866 ( .A(\u_coder/N473 ), .Q(n1761) );
  NOR21 U867 ( .A(n814), .B(n1760), .Q(\u_coder/N519 ) );
  INV3 U868 ( .A(\u_coder/N474 ), .Q(n1760) );
  INV3 U869 ( .A(\u_cordic/my_rotation/n70 ), .Q(n1514) );
  NAND22 U870 ( .A(\u_cordic/my_rotation/next_delta [14]), .B(n975), .Q(
        \u_cordic/my_rotation/n70 ) );
  XOR21 U871 ( .A(\u_decoder/iq_demod/dp_cluster_1/mult_150/SUMB[3][1] ), .B(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/CARRYB[3][0] ), .Q(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/A1[2] ) );
  NAND31 U872 ( .A(n1135), .B(n1136), .C(n976), .Q(n1134) );
  NAND31 U873 ( .A(n978), .B(n1137), .C(n1136), .Q(n1138) );
  XOR21 U874 ( .A(n961), .B(
        \u_decoder/fir_filter/dp_cluster_0/r164/SUMB[7][0] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r164/A1[5] ) );
  XOR21 U875 ( .A(n963), .B(
        \u_decoder/fir_filter/dp_cluster_0/r177/SUMB[7][0] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r177/A1[5] ) );
  XOR21 U876 ( .A(n960), .B(
        \u_decoder/fir_filter/dp_cluster_0/r167/SUMB[6][3] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r167/SUMB[7][2] ) );
  XOR21 U877 ( .A(n962), .B(
        \u_decoder/fir_filter/dp_cluster_0/r180/SUMB[6][3] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r180/SUMB[7][2] ) );
  XOR21 U878 ( .A(\u_decoder/I_prefilter [6]), .B(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[6][5] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/SUMB[7][5] ) );
  XOR21 U879 ( .A(\u_decoder/I_prefilter [6]), .B(
        \u_decoder/fir_filter/dp_cluster_0/r166/CARRYB[6][3] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r166/SUMB[7][3] ) );
  XOR21 U880 ( .A(\u_decoder/Q_prefilter [6]), .B(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[6][5] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/SUMB[7][5] ) );
  XOR21 U881 ( .A(\u_decoder/Q_prefilter [6]), .B(
        \u_decoder/fir_filter/dp_cluster_0/r179/CARRYB[6][3] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r179/SUMB[7][3] ) );
  NOR21 U882 ( .A(n593), .B(n594), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r165/A2[6] ) );
  INV3 U883 ( .A(n961), .Q(n594) );
  INV3 U884 ( .A(\u_decoder/fir_filter/dp_cluster_0/r165/SUMB[7][0] ), .Q(n593) );
  NOR21 U885 ( .A(n655), .B(n656), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r178/A2[6] ) );
  INV3 U886 ( .A(n963), .Q(n656) );
  INV3 U887 ( .A(\u_decoder/fir_filter/dp_cluster_0/r178/SUMB[7][0] ), .Q(n655) );
  XOR21 U888 ( .A(n771), .B(n773), .Q(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/SUMB[2][3] ) );
  XOR21 U889 ( .A(n761), .B(n763), .Q(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/SUMB[2][3] ) );
  NOR21 U890 ( .A(n69), .B(n51), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[3][3] ) );
  NOR21 U891 ( .A(n70), .B(n52), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[3][3] ) );
  NOR21 U892 ( .A(n52), .B(n70), .Q(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[3][0] ) );
  NOR21 U893 ( .A(n229), .B(n739), .Q(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[7][2] ) );
  INV3 U894 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_276/SUMB[6][3] ), .Q(
        n739) );
  NOR21 U895 ( .A(n230), .B(n728), .Q(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[7][2] ) );
  INV3 U896 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_308/SUMB[6][3] ), .Q(
        n728) );
  NOR21 U897 ( .A(n229), .B(n738), .Q(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[7][1] ) );
  INV3 U898 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_276/SUMB[5][3] ), .Q(
        n738) );
  NOR21 U899 ( .A(n230), .B(n727), .Q(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[7][1] ) );
  INV3 U900 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_308/SUMB[5][3] ), .Q(
        n727) );
  NOR21 U901 ( .A(n229), .B(n744), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r165/CARRYB[7][1] ) );
  INV3 U902 ( .A(\u_decoder/fir_filter/dp_cluster_0/r165/SUMB[5][3] ), .Q(n744) );
  NOR21 U903 ( .A(n230), .B(n733), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r178/CARRYB[7][1] ) );
  INV3 U904 ( .A(\u_decoder/fir_filter/dp_cluster_0/r178/SUMB[5][3] ), .Q(n733) );
  NOR21 U905 ( .A(n229), .B(n745), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r165/CARRYB[7][2] ) );
  INV3 U906 ( .A(\u_decoder/fir_filter/dp_cluster_0/r165/SUMB[6][3] ), .Q(n745) );
  NOR21 U907 ( .A(n230), .B(n734), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r178/CARRYB[7][2] ) );
  INV3 U908 ( .A(\u_decoder/fir_filter/dp_cluster_0/r178/SUMB[6][3] ), .Q(n734) );
  XNR21 U909 ( .A(n2321), .B(n2322), .Q(
        \u_decoder/iq_demod/dp_cluster_1/mult_I_sin_out [5]) );
  XNR21 U910 ( .A(n2328), .B(n2329), .Q(
        \u_decoder/iq_demod/dp_cluster_1/mult_Q_cos_out [5]) );
  NAND22 U911 ( .A(\u_decoder/iq_demod/dp_cluster_1/mult_149/A2[2] ), .B(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/A1[2] ), .Q(n2321) );
  NOR21 U912 ( .A(n606), .B(n229), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r164/A2[6] ) );
  INV3 U913 ( .A(\u_decoder/fir_filter/dp_cluster_0/r164/SUMB[7][0] ), .Q(n606) );
  NOR21 U914 ( .A(n668), .B(n230), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r177/A2[6] ) );
  INV3 U915 ( .A(\u_decoder/fir_filter/dp_cluster_0/r177/SUMB[7][0] ), .Q(n668) );
  NOR31 U916 ( .A(n1781), .B(n2242), .C(n986), .Q(n2622) );
  INV3 U917 ( .A(\u_cdr/phd1/cnt_phd/N76 ), .Q(n2242) );
  INV3 U918 ( .A(n2629), .Q(n1781) );
  NOR31 U919 ( .A(n1782), .B(n2238), .C(n986), .Q(n2635) );
  INV3 U920 ( .A(\u_cdr/dec1/cnt_dec/N76 ), .Q(n2238) );
  INV3 U921 ( .A(n2642), .Q(n1782) );
  NOR31 U922 ( .A(n1783), .B(n2237), .C(n985), .Q(\u_cdr/div1/cnt_div/n41 ) );
  INV3 U923 ( .A(\u_cdr/div1/cnt_div/N76 ), .Q(n2237) );
  INV3 U924 ( .A(\u_cdr/div1/cnt_div/n48 ), .Q(n1783) );
  NOR21 U925 ( .A(n229), .B(n740), .Q(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[7][4] ) );
  INV3 U926 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_276/SUMB[6][5] ), .Q(
        n740) );
  NOR21 U927 ( .A(n229), .B(n743), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r166/CARRYB[7][2] ) );
  INV3 U928 ( .A(\u_decoder/fir_filter/dp_cluster_0/r166/SUMB[6][3] ), .Q(n743) );
  NOR21 U929 ( .A(n230), .B(n729), .Q(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[7][4] ) );
  INV3 U930 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_308/SUMB[6][5] ), .Q(
        n729) );
  NOR21 U931 ( .A(n230), .B(n732), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r179/CARRYB[7][2] ) );
  INV3 U932 ( .A(\u_decoder/fir_filter/dp_cluster_0/r179/SUMB[6][3] ), .Q(n732) );
  INV3 U933 ( .A(\u_decoder/iq_demod/dp_cluster_1/mult_150/ab[0][3] ), .Q(n708) );
  NOR21 U934 ( .A(n51), .B(n69), .Q(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[3][0] ) );
  NAND22 U935 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_276/SUMB[7][0] ), 
        .B(n960), .Q(n352) );
  NAND22 U936 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_308/SUMB[7][0] ), 
        .B(n962), .Q(n353) );
  NOR21 U937 ( .A(n814), .B(n1762), .Q(\u_coder/N517 ) );
  INV3 U938 ( .A(\u_coder/N472 ), .Q(n1762) );
  INV3 U939 ( .A(\u_decoder/iq_demod/n57 ), .Q(n1941) );
  AOI221 U940 ( .A(\u_decoder/iq_demod/add_Q_out [7]), .B(n790), .C(n963), .D(
        n752), .Q(\u_decoder/iq_demod/n57 ) );
  INV3 U941 ( .A(\u_cordic/my_rotation/n72 ), .Q(n1516) );
  NAND22 U942 ( .A(\u_cordic/my_rotation/next_delta [12]), .B(n975), .Q(
        \u_cordic/my_rotation/n72 ) );
  INV3 U943 ( .A(\u_cordic/my_rotation/n71 ), .Q(n1515) );
  NAND22 U944 ( .A(\u_cordic/my_rotation/next_delta [13]), .B(n975), .Q(
        \u_cordic/my_rotation/n71 ) );
  XOR21 U945 ( .A(\u_decoder/iq_demod/dp_cluster_0/mult_151/SUMB[3][1] ), .B(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/CARRYB[3][0] ), .Q(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/A1[2] ) );
  XOR21 U946 ( .A(\u_decoder/iq_demod/dp_cluster_1/mult_149/SUMB[3][1] ), .B(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/CARRYB[3][0] ), .Q(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/A1[2] ) );
  XOR21 U947 ( .A(\u_decoder/iq_demod/dp_cluster_0/mult_148/SUMB[3][1] ), .B(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/CARRYB[3][0] ), .Q(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/A1[2] ) );
  XOR21 U948 ( .A(\u_decoder/iq_demod/dp_cluster_0/mult_151/SUMB[3][2] ), .B(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/CARRYB[3][1] ), .Q(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/A1[3] ) );
  XOR21 U949 ( .A(\u_decoder/iq_demod/dp_cluster_1/mult_150/SUMB[3][2] ), .B(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/CARRYB[3][1] ), .Q(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/A1[3] ) );
  XOR21 U950 ( .A(\u_decoder/iq_demod/dp_cluster_1/mult_149/SUMB[3][2] ), .B(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/CARRYB[3][1] ), .Q(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/A1[3] ) );
  XOR21 U951 ( .A(\u_decoder/iq_demod/dp_cluster_0/mult_148/SUMB[3][2] ), .B(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/CARRYB[3][1] ), .Q(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/A1[3] ) );
  XOR21 U952 ( .A(n767), .B(
        \u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[6][3] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r167/SUMB[7][3] ) );
  XOR21 U953 ( .A(n757), .B(
        \u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[6][3] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r180/SUMB[7][3] ) );
  NOR21 U954 ( .A(n982), .B(n2629), .Q(n2623) );
  NOR21 U955 ( .A(n980), .B(n2642), .Q(n2636) );
  NOR21 U956 ( .A(n980), .B(\u_cdr/div1/cnt_div/n48 ), .Q(
        \u_cdr/div1/cnt_div/n42 ) );
  NOR21 U957 ( .A(n24), .B(n101), .Q(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/ab[1][0] ) );
  NOR21 U958 ( .A(n28), .B(n101), .Q(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/ab[1][2] ) );
  NOR21 U959 ( .A(n26), .B(n101), .Q(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/ab[1][1] ) );
  NOR21 U960 ( .A(n25), .B(n101), .Q(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/ab[1][2] ) );
  NOR21 U961 ( .A(n23), .B(n101), .Q(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/ab[1][1] ) );
  NOR21 U962 ( .A(n28), .B(n102), .Q(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/ab[1][2] ) );
  NOR21 U963 ( .A(n26), .B(n102), .Q(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/ab[1][1] ) );
  NOR21 U964 ( .A(n25), .B(n102), .Q(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/ab[1][2] ) );
  NOR21 U965 ( .A(n23), .B(n102), .Q(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/ab[1][1] ) );
  NOR21 U966 ( .A(n27), .B(n101), .Q(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/ab[1][0] ) );
  NOR21 U967 ( .A(n24), .B(n102), .Q(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/ab[1][0] ) );
  NOR21 U968 ( .A(n27), .B(n102), .Q(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/ab[1][0] ) );
  NOR21 U969 ( .A(n26), .B(n104), .Q(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/ab[0][1] ) );
  NOR21 U970 ( .A(n28), .B(n104), .Q(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/ab[0][2] ) );
  NOR21 U971 ( .A(n25), .B(n104), .Q(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/ab[0][2] ) );
  NOR21 U972 ( .A(n28), .B(n103), .Q(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/ab[0][2] ) );
  NOR21 U973 ( .A(n25), .B(n103), .Q(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/ab[0][2] ) );
  NOR21 U974 ( .A(n23), .B(n104), .Q(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/ab[0][1] ) );
  NOR21 U975 ( .A(n26), .B(n103), .Q(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/ab[0][1] ) );
  NOR21 U976 ( .A(n23), .B(n103), .Q(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/ab[0][1] ) );
  NOR21 U977 ( .A(n698), .B(n699), .Q(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/A2[3] ) );
  INV3 U978 ( .A(\u_decoder/iq_demod/dp_cluster_1/mult_150/CARRYB[3][0] ), .Q(
        n698) );
  INV3 U979 ( .A(\u_decoder/iq_demod/dp_cluster_1/mult_150/SUMB[3][1] ), .Q(
        n699) );
  NOR21 U980 ( .A(n686), .B(n687), .Q(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/A2[3] ) );
  INV3 U981 ( .A(\u_decoder/iq_demod/dp_cluster_0/mult_148/CARRYB[3][0] ), .Q(
        n686) );
  INV3 U982 ( .A(\u_decoder/iq_demod/dp_cluster_0/mult_148/SUMB[3][1] ), .Q(
        n687) );
  NOR21 U983 ( .A(n674), .B(n675), .Q(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/A2[3] ) );
  INV3 U984 ( .A(\u_decoder/iq_demod/dp_cluster_0/mult_151/CARRYB[3][0] ), .Q(
        n674) );
  INV3 U985 ( .A(\u_decoder/iq_demod/dp_cluster_0/mult_151/SUMB[3][1] ), .Q(
        n675) );
  NOR21 U986 ( .A(n710), .B(n711), .Q(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/A2[3] ) );
  INV3 U987 ( .A(\u_decoder/iq_demod/dp_cluster_1/mult_149/CARRYB[3][0] ), .Q(
        n710) );
  INV3 U988 ( .A(\u_decoder/iq_demod/dp_cluster_1/mult_149/SUMB[3][1] ), .Q(
        n711) );
  NOR21 U989 ( .A(n125), .B(n24), .Q(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/ab[2][0] ) );
  NOR21 U990 ( .A(n680), .B(n681), .Q(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/CARRYB[1][0] ) );
  XOR21 U991 ( .A(\u_decoder/iq_demod/dp_cluster_0/mult_151/ab[0][2] ), .B(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/ab[1][1] ), .Q(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/SUMB[1][1] ) );
  NOR21 U992 ( .A(n125), .B(n23), .Q(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/ab[2][1] ) );
  NOR21 U993 ( .A(n706), .B(n707), .Q(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/CARRYB[1][1] ) );
  XOR21 U994 ( .A(\u_decoder/iq_demod/dp_cluster_1/mult_150/ab[0][3] ), .B(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/ab[1][2] ), .Q(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/SUMB[1][2] ) );
  NOR21 U995 ( .A(n125), .B(n27), .Q(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/ab[2][0] ) );
  NOR21 U996 ( .A(n704), .B(n705), .Q(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/CARRYB[1][0] ) );
  XOR21 U997 ( .A(\u_decoder/iq_demod/dp_cluster_1/mult_150/ab[0][2] ), .B(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/ab[1][1] ), .Q(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/SUMB[1][1] ) );
  NOR21 U998 ( .A(n126), .B(n26), .Q(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/ab[2][1] ) );
  NOR21 U999 ( .A(n718), .B(n719), .Q(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/CARRYB[1][1] ) );
  XOR21 U1000 ( .A(\u_decoder/iq_demod/dp_cluster_1/mult_149/ab[0][3] ), .B(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/ab[1][2] ), .Q(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/SUMB[1][2] ) );
  NOR21 U1001 ( .A(n126), .B(n24), .Q(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/ab[2][0] ) );
  NOR21 U1002 ( .A(n716), .B(n717), .Q(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/CARRYB[1][0] ) );
  XOR21 U1003 ( .A(\u_decoder/iq_demod/dp_cluster_1/mult_149/ab[0][2] ), .B(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/ab[1][1] ), .Q(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/SUMB[1][1] ) );
  NOR21 U1004 ( .A(n126), .B(n23), .Q(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/ab[2][1] ) );
  NOR21 U1005 ( .A(n694), .B(n695), .Q(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/CARRYB[1][1] ) );
  XOR21 U1006 ( .A(\u_decoder/iq_demod/dp_cluster_0/mult_148/ab[0][3] ), .B(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/ab[1][2] ), .Q(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/SUMB[1][2] ) );
  NOR21 U1007 ( .A(n126), .B(n27), .Q(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/ab[2][0] ) );
  NOR21 U1008 ( .A(n692), .B(n693), .Q(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/CARRYB[1][0] ) );
  XOR21 U1009 ( .A(\u_decoder/iq_demod/dp_cluster_0/mult_148/ab[0][2] ), .B(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/ab[1][1] ), .Q(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/SUMB[1][1] ) );
  NOR21 U1010 ( .A(n814), .B(n1764), .Q(\u_coder/N515 ) );
  INV3 U1011 ( .A(\u_coder/N470 ), .Q(n1764) );
  NOR21 U1012 ( .A(n229), .B(n737), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[7][2] ) );
  INV3 U1013 ( .A(\u_decoder/fir_filter/dp_cluster_0/r167/SUMB[6][3] ), .Q(
        n737) );
  NOR21 U1014 ( .A(n230), .B(n726), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[7][2] ) );
  INV3 U1015 ( .A(\u_decoder/fir_filter/dp_cluster_0/r180/SUMB[6][3] ), .Q(
        n726) );
  INV3 U1016 ( .A(\u_decoder/iq_demod/dp_cluster_0/mult_Q_sin_out [3]), .Q(
        n1950) );
  NAND22 U1017 ( .A(\u_decoder/iq_demod/dp_cluster_0/mult_151/A2[2] ), .B(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/A1[2] ), .Q(n2342) );
  NAND22 U1018 ( .A(\u_decoder/iq_demod/dp_cluster_1/mult_150/A2[2] ), .B(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/A1[2] ), .Q(n2328) );
  NAND22 U1019 ( .A(\u_decoder/iq_demod/dp_cluster_0/mult_148/A2[2] ), .B(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/A1[2] ), .Q(n2335) );
  NOR21 U1020 ( .A(n125), .B(n26), .Q(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/ab[2][1] ) );
  NOR21 U1021 ( .A(n682), .B(n683), .Q(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/CARRYB[1][1] ) );
  XOR21 U1022 ( .A(\u_decoder/iq_demod/dp_cluster_0/mult_151/ab[0][3] ), .B(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/ab[1][2] ), .Q(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/SUMB[1][2] ) );
  INV3 U1023 ( .A(\u_decoder/iq_demod/dp_cluster_0/mult_151/A2[2] ), .Q(n1949)
         );
  INV3 U1024 ( .A(\u_decoder/iq_demod/dp_cluster_1/mult_150/A2[2] ), .Q(n1945)
         );
  INV3 U1025 ( .A(\u_decoder/iq_demod/dp_cluster_1/mult_149/A2[2] ), .Q(n1955)
         );
  INV3 U1026 ( .A(\u_decoder/iq_demod/dp_cluster_0/mult_148/A2[2] ), .Q(n1958)
         );
  INV3 U1027 ( .A(\u_decoder/iq_demod/dp_cluster_0/mult_151/ab[0][3] ), .Q(
        n684) );
  INV3 U1028 ( .A(\u_decoder/iq_demod/dp_cluster_1/mult_149/ab[0][3] ), .Q(
        n720) );
  INV3 U1029 ( .A(\u_decoder/iq_demod/dp_cluster_0/mult_148/ab[0][3] ), .Q(
        n696) );
  NOR21 U1030 ( .A(\u_coder/n315 ), .B(n1763), .Q(\u_coder/N516 ) );
  INV3 U1031 ( .A(\u_coder/N471 ), .Q(n1763) );
  INV3 U1032 ( .A(\u_decoder/iq_demod/n56 ), .Q(n1940) );
  AOI221 U1033 ( .A(\u_decoder/iq_demod/add_Q_out [6]), .B(n790), .C(
        \u_decoder/Q_prefilter [6]), .D(n752), .Q(\u_decoder/iq_demod/n56 ) );
  INV3 U1034 ( .A(\u_decoder/iq_demod/n49 ), .Q(n1870) );
  AOI221 U1035 ( .A(\u_decoder/iq_demod/add_I_out [7]), .B(n790), .C(n961), 
        .D(n753), .Q(\u_decoder/iq_demod/n49 ) );
  INV3 U1036 ( .A(\u_decoder/iq_demod/n48 ), .Q(n1869) );
  AOI221 U1037 ( .A(\u_decoder/iq_demod/add_I_out [6]), .B(n790), .C(
        \u_decoder/I_prefilter [6]), .D(n753), .Q(\u_decoder/iq_demod/n48 ) );
  INV3 U1038 ( .A(n2632), .Q(n1493) );
  NAND22 U1039 ( .A(\u_cdr/phd1/cnt_phd/N42 ), .B(n975), .Q(n2632) );
  NOR40 U1040 ( .A(n2612), .B(n2611), .C(n2239), .D(\u_cdr/phd1/cnt_phd/N41 ), 
        .Q(\u_cdr/phd1/cnt_phd/N42 ) );
  NAND22 U1041 ( .A(n2241), .B(n2610), .Q(n2611) );
  INV3 U1042 ( .A(\u_cordic/my_rotation/n73 ), .Q(n1517) );
  NAND22 U1043 ( .A(\u_cordic/my_rotation/next_delta [11]), .B(n975), .Q(
        \u_cordic/my_rotation/n73 ) );
  XOR21 U1044 ( .A(\u_decoder/iq_demod/dp_cluster_0/mult_151/SUMB[3][3] ), .B(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/CARRYB[3][2] ), .Q(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/A1[4] ) );
  XOR21 U1045 ( .A(\u_decoder/iq_demod/dp_cluster_1/mult_150/SUMB[3][3] ), .B(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/CARRYB[3][2] ), .Q(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/A1[4] ) );
  XOR21 U1046 ( .A(\u_decoder/iq_demod/dp_cluster_1/mult_149/SUMB[3][3] ), .B(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/CARRYB[3][2] ), .Q(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/A1[4] ) );
  XOR21 U1047 ( .A(\u_decoder/iq_demod/dp_cluster_0/mult_148/SUMB[3][3] ), .B(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/CARRYB[3][2] ), .Q(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/A1[4] ) );
  NOR40 U1048 ( .A(n2268), .B(n1705), .C(n2267), .D(n1701), .Q(
        \sig_MUX_inMUX5[0] ) );
  INV3 U1049 ( .A(n2266), .Q(n1701) );
  INV3 U1050 ( .A(n2265), .Q(n1705) );
  NAND22 U1051 ( .A(n1700), .B(n2264), .Q(n2268) );
  AOI211 U1052 ( .A(n2594), .B(n2593), .C(n2223), .Q(n2595) );
  NOR40 U1053 ( .A(n2236), .B(n2235), .C(n2234), .D(n2592), .Q(n2594) );
  NOR40 U1054 ( .A(n2224), .B(n2225), .C(n2231), .D(n2230), .Q(n2593) );
  AOI211 U1055 ( .A(\u_cordic/my_rotation/n64 ), .B(n2591), .C(
        \u_cordic/my_rotation/n63 ), .Q(n2592) );
  NOR21 U1056 ( .A(n37), .B(n554), .Q(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[7][5] ) );
  INV3 U1057 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[6][5] ), 
        .Q(n554) );
  NOR21 U1058 ( .A(n38), .B(n616), .Q(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[7][5] ) );
  INV3 U1059 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[6][5] ), 
        .Q(n616) );
  INV3 U1060 ( .A(\u_cordic/my_rotation/n100 ), .Q(n2223) );
  AOI221 U1061 ( .A(n748), .B(n33), .C(\u_cordic/my_rotation/N56 ), .D(n747), 
        .Q(\u_cordic/my_rotation/n100 ) );
  XOR21 U1062 ( .A(\u_cordic/my_rotation/add_43/carry [15]), .B(n747), .Q(
        \u_cordic/my_rotation/N56 ) );
  NOR21 U1063 ( .A(n477), .B(n267), .Q(\u_cordic/my_rotation/add_43/carry [15]) );
  INV3 U1064 ( .A(\u_cordic/my_rotation/n85 ), .Q(n1529) );
  NAND31 U1065 ( .A(n978), .B(\u_cordic/my_rotation/n86 ), .C(n2222), .Q(
        \u_cordic/my_rotation/n85 ) );
  INV3 U1066 ( .A(n2595), .Q(n2222) );
  NAND41 U1067 ( .A(\u_cordic/my_rotation/n87 ), .B(\u_cordic/my_rotation/n88 ), .C(\u_cordic/my_rotation/n89 ), .D(\u_cordic/my_rotation/n90 ), .Q(
        \u_cordic/my_rotation/n86 ) );
  NOR21 U1068 ( .A(n37), .B(n582), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r166/CARRYB[7][3] ) );
  INV3 U1069 ( .A(\u_decoder/fir_filter/dp_cluster_0/r166/CARRYB[6][3] ), .Q(
        n582) );
  NOR21 U1070 ( .A(n38), .B(n644), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r179/CARRYB[7][3] ) );
  INV3 U1071 ( .A(\u_decoder/fir_filter/dp_cluster_0/r179/CARRYB[6][3] ), .Q(
        n644) );
  NOR21 U1072 ( .A(\u_coder/n315 ), .B(n1765), .Q(\u_coder/N514 ) );
  INV3 U1073 ( .A(\u_coder/N469 ), .Q(n1765) );
  INV3 U1074 ( .A(\u_coder/n155 ), .Q(n1660) );
  NOR21 U1075 ( .A(n164), .B(n569), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[7][3] ) );
  INV3 U1076 ( .A(\u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[6][3] ), .Q(
        n569) );
  NOR21 U1077 ( .A(n165), .B(n631), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[7][3] ) );
  INV3 U1078 ( .A(\u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[6][3] ), .Q(
        n631) );
  INV3 U1079 ( .A(n2262), .Q(n1700) );
  NOR21 U1080 ( .A(n700), .B(n701), .Q(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/A2[4] ) );
  INV3 U1081 ( .A(\u_decoder/iq_demod/dp_cluster_1/mult_150/CARRYB[3][1] ), 
        .Q(n700) );
  INV3 U1082 ( .A(\u_decoder/iq_demod/dp_cluster_1/mult_150/SUMB[3][2] ), .Q(
        n701) );
  NOR21 U1083 ( .A(n712), .B(n713), .Q(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/A2[4] ) );
  INV3 U1084 ( .A(\u_decoder/iq_demod/dp_cluster_1/mult_149/CARRYB[3][1] ), 
        .Q(n712) );
  INV3 U1085 ( .A(\u_decoder/iq_demod/dp_cluster_1/mult_149/SUMB[3][2] ), .Q(
        n713) );
  NOR21 U1086 ( .A(n688), .B(n689), .Q(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/A2[4] ) );
  INV3 U1087 ( .A(\u_decoder/iq_demod/dp_cluster_0/mult_148/CARRYB[3][1] ), 
        .Q(n688) );
  INV3 U1088 ( .A(\u_decoder/iq_demod/dp_cluster_0/mult_148/SUMB[3][2] ), .Q(
        n689) );
  NOR21 U1089 ( .A(n676), .B(n677), .Q(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/A2[4] ) );
  INV3 U1090 ( .A(\u_decoder/iq_demod/dp_cluster_0/mult_151/CARRYB[3][1] ), 
        .Q(n676) );
  INV3 U1091 ( .A(\u_decoder/iq_demod/dp_cluster_0/mult_151/SUMB[3][2] ), .Q(
        n677) );
  INV3 U1092 ( .A(\u_cordic/my_rotation/add_43/carry [14]), .Q(n477) );
  INV3 U1093 ( .A(\u_cordic/mycordic/r173/carry [14]), .Q(n483) );
  INV3 U1094 ( .A(\u_decoder/iq_demod/n55 ), .Q(n1938) );
  AOI221 U1095 ( .A(\u_decoder/iq_demod/add_Q_out [5]), .B(n790), .C(
        \u_decoder/Q_prefilter [5]), .D(n752), .Q(\u_decoder/iq_demod/n55 ) );
  INV3 U1096 ( .A(\u_decoder/iq_demod/n47 ), .Q(n1867) );
  AOI221 U1097 ( .A(\u_decoder/iq_demod/add_I_out [5]), .B(n790), .C(
        \u_decoder/I_prefilter [5]), .D(n753), .Q(\u_decoder/iq_demod/n47 ) );
  INV3 U1098 ( .A(\u_decoder/iq_demod/n46 ), .Q(n1866) );
  AOI221 U1099 ( .A(\u_decoder/iq_demod/add_I_out [4]), .B(n790), .C(n766), 
        .D(n753), .Q(\u_decoder/iq_demod/n46 ) );
  INV3 U1100 ( .A(\u_coder/n304 ), .Q(n1592) );
  AOI221 U1101 ( .A(n778), .B(n813), .C(n811), .D(\u_coder/n89 ), .Q(
        \u_coder/n304 ) );
  INV3 U1102 ( .A(\u_cordic/my_rotation/n75 ), .Q(n1519) );
  NAND22 U1103 ( .A(\u_cordic/my_rotation/next_delta [9]), .B(n974), .Q(
        \u_cordic/my_rotation/n75 ) );
  INV3 U1104 ( .A(\u_cordic/my_rotation/n74 ), .Q(n1518) );
  NAND22 U1105 ( .A(\u_cordic/my_rotation/next_delta [10]), .B(n975), .Q(
        \u_cordic/my_rotation/n74 ) );
  AOI2111 U1106 ( .A(\u_coder/n234 ), .B(\u_coder/n76 ), .C(n1726), .D(n1473), 
        .Q(\u_coder/n246 ) );
  AOI2111 U1107 ( .A(\u_coder/n189 ), .B(\u_coder/n72 ), .C(n1714), .D(
        \u_coder/n273 ), .Q(\u_coder/n265 ) );
  NOR40 U1108 ( .A(n2255), .B(\u_inFIFO/N125 ), .C(\u_inFIFO/N127 ), .D(
        \u_inFIFO/N126 ), .Q(\u_inFIFO/N249 ) );
  NAND22 U1109 ( .A(n2254), .B(\u_inFIFO/N128 ), .Q(n2255) );
  NOR21 U1110 ( .A(\u_inFIFO/N124 ), .B(\u_inFIFO/N123 ), .Q(n2254) );
  NOR21 U1111 ( .A(n6), .B(\u_decoder/iq_demod/I_if_buff[3] ), .Q(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/ab[3][3] ) );
  NOR21 U1112 ( .A(n6), .B(\u_decoder/iq_demod/Q_if_buff[3] ), .Q(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/ab[3][3] ) );
  NOR21 U1113 ( .A(n5), .B(\u_decoder/iq_demod/I_if_buff[3] ), .Q(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/ab[3][3] ) );
  NOR21 U1114 ( .A(n5), .B(\u_decoder/iq_demod/Q_if_buff[3] ), .Q(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/ab[3][3] ) );
  NAND31 U1115 ( .A(\u_coder/n185 ), .B(\u_coder/n186 ), .C(n1590), .Q(
        \u_coder/n152 ) );
  INV3 U1116 ( .A(\u_coder/n187 ), .Q(n1590) );
  OAI311 U1117 ( .A(\u_coder/n189 ), .B(\u_coder/n154 ), .C(\u_coder/n168 ), 
        .D(\u_coder/n72 ), .Q(\u_coder/n185 ) );
  AOI211 U1118 ( .A(\u_outFIFO/n540 ), .B(n1791), .C(\u_outFIFO/n542 ), .Q(
        \u_outFIFO/n541 ) );
  INV3 U1119 ( .A(\u_outFIFO/N474 ), .Q(n1791) );
  BUF6 U1120 ( .A(\u_coder/n282 ), .Q(n809) );
  NOR21 U1121 ( .A(n27), .B(n103), .Q(
        \u_decoder/iq_demod/dp_cluster_0/mult_I_cos_out [0]) );
  AOI221 U1122 ( .A(\u_inFIFO/n234 ), .B(n1699), .C(\u_inFIFO/n233 ), .D(n2262), .Q(\u_inFIFO/n235 ) );
  NOR21 U1123 ( .A(n27), .B(n104), .Q(
        \u_decoder/iq_demod/dp_cluster_1/mult_Q_cos_out [0]) );
  NOR21 U1124 ( .A(n24), .B(n103), .Q(
        \u_decoder/iq_demod/dp_cluster_1/mult_I_sin_out [0]) );
  NOR21 U1125 ( .A(n814), .B(n1766), .Q(\u_coder/N513 ) );
  INV3 U1126 ( .A(\u_coder/N468 ), .Q(n1766) );
  AOI311 U1127 ( .A(\u_inFIFO/n237 ), .B(\u_inFIFO/n209 ), .C(\u_inFIFO/n242 ), 
        .D(n987), .Q(\u_inFIFO/N41 ) );
  AOI311 U1128 ( .A(n1698), .B(\u_inFIFO/n230 ), .C(\u_inFIFO/sig_fsm_start_R ), .D(\u_inFIFO/n243 ), .Q(\u_inFIFO/n242 ) );
  NOR21 U1129 ( .A(n1699), .B(\u_inFIFO/n236 ), .Q(\u_inFIFO/n243 ) );
  INV3 U1130 ( .A(\u_coder/n229 ), .Q(n1472) );
  NAND31 U1131 ( .A(\u_coder/n230 ), .B(\u_coder/n231 ), .C(\u_coder/n232 ), 
        .Q(\u_coder/n229 ) );
  AOI211 U1132 ( .A(n1756), .B(\u_coder/n233 ), .C(n985), .Q(\u_coder/n232 )
         );
  OAI311 U1133 ( .A(\u_coder/n234 ), .B(\u_coder/n220 ), .C(\u_coder/n218 ), 
        .D(\u_coder/n76 ), .Q(\u_coder/n231 ) );
  NOR21 U1134 ( .A(n981), .B(\u_coder/n205 ), .Q(\u_coder/n256 ) );
  NOR40 U1135 ( .A(n2302), .B(\u_outFIFO/N133 ), .C(\u_outFIFO/N135 ), .D(
        \u_outFIFO/N134 ), .Q(\u_outFIFO/N473 ) );
  NAND22 U1136 ( .A(n2301), .B(\u_outFIFO/N136 ), .Q(n2302) );
  NOR21 U1137 ( .A(\u_outFIFO/N132 ), .B(\u_outFIFO/N131 ), .Q(n2301) );
  INV3 U1138 ( .A(\u_decoder/iq_demod/dp_cluster_0/mult_Q_sin_out [0]), .Q(
        n1946) );
  NOR21 U1139 ( .A(n24), .B(n104), .Q(
        \u_decoder/iq_demod/dp_cluster_0/mult_Q_sin_out [0]) );
  INV3 U1140 ( .A(\u_coder/n205 ), .Q(n1661) );
  INV3 U1141 ( .A(\u_decoder/iq_demod/dp_cluster_0/mult_151/CARRYB[3][2] ), 
        .Q(n678) );
  INV3 U1142 ( .A(\u_decoder/iq_demod/dp_cluster_1/mult_150/CARRYB[3][2] ), 
        .Q(n702) );
  NOR21 U1143 ( .A(n690), .B(n691), .Q(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/A2[5] ) );
  INV3 U1144 ( .A(\u_decoder/iq_demod/dp_cluster_0/mult_148/SUMB[3][3] ), .Q(
        n691) );
  INV3 U1145 ( .A(\u_decoder/iq_demod/dp_cluster_0/mult_148/CARRYB[3][2] ), 
        .Q(n690) );
  XNR21 U1146 ( .A(n960), .B(
        \u_decoder/fir_filter/dp_cluster_0/r167/SUMB[7][0] ), .Q(n354) );
  XNR21 U1147 ( .A(n960), .B(
        \u_decoder/fir_filter/dp_cluster_0/r166/SUMB[7][0] ), .Q(n355) );
  XNR21 U1148 ( .A(n962), .B(
        \u_decoder/fir_filter/dp_cluster_0/r180/SUMB[7][0] ), .Q(n356) );
  XNR21 U1149 ( .A(n962), .B(
        \u_decoder/fir_filter/dp_cluster_0/r179/SUMB[7][0] ), .Q(n357) );
  NOR21 U1150 ( .A(n714), .B(n715), .Q(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/A2[5] ) );
  INV3 U1151 ( .A(\u_decoder/iq_demod/dp_cluster_1/mult_149/SUMB[3][3] ), .Q(
        n715) );
  INV3 U1152 ( .A(\u_decoder/iq_demod/dp_cluster_1/mult_149/CARRYB[3][2] ), 
        .Q(n714) );
  INV3 U1153 ( .A(\u_cordic/mycordic/add_262/carry [14]), .Q(n545) );
  NOR21 U1154 ( .A(\u_coder/n315 ), .B(n1767), .Q(\u_coder/N512 ) );
  INV3 U1155 ( .A(\u_coder/N467 ), .Q(n1767) );
  INV3 U1156 ( .A(\u_decoder/iq_demod/n54 ), .Q(n1937) );
  AOI221 U1157 ( .A(\u_decoder/iq_demod/add_Q_out [4]), .B(n790), .C(n756), 
        .D(n752), .Q(\u_decoder/iq_demod/n54 ) );
  INV3 U1158 ( .A(\u_decoder/iq_demod/n53 ), .Q(n1936) );
  AOI221 U1159 ( .A(\u_decoder/iq_demod/add_Q_out [3]), .B(n790), .C(n758), 
        .D(n752), .Q(\u_decoder/iq_demod/n53 ) );
  INV3 U1160 ( .A(\u_decoder/iq_demod/n45 ), .Q(n1865) );
  AOI221 U1161 ( .A(\u_decoder/iq_demod/add_I_out [3]), .B(n790), .C(n768), 
        .D(n753), .Q(\u_decoder/iq_demod/n45 ) );
  INV3 U1162 ( .A(\u_cordic/my_rotation/n76 ), .Q(n1520) );
  NAND22 U1163 ( .A(\u_cordic/my_rotation/next_delta [8]), .B(n975), .Q(
        \u_cordic/my_rotation/n76 ) );
  XOR21 U1164 ( .A(n960), .B(n765), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r167/SUMB[7][4] ) );
  XOR21 U1165 ( .A(n962), .B(n755), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r180/SUMB[7][4] ) );
  XOR21 U1166 ( .A(n960), .B(n764), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r167/SUMB[7][5] ) );
  XOR21 U1167 ( .A(n962), .B(n754), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r180/SUMB[7][5] ) );
  XOR21 U1168 ( .A(n960), .B(n37), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r165/SUMB[7][4] ) );
  XOR21 U1169 ( .A(n962), .B(n38), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r178/SUMB[7][4] ) );
  XOR21 U1170 ( .A(n961), .B(n37), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r164/SUMB[7][3] ) );
  XOR21 U1171 ( .A(n963), .B(n38), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r177/SUMB[7][3] ) );
  AOI211 U1172 ( .A(\u_coder/n195 ), .B(n1709), .C(\u_coder/n162 ), .Q(
        \u_coder/n156 ) );
  NAND22 U1173 ( .A(n2202), .B(\u_decoder/fir_filter/n1153 ), .Q(
        \u_decoder/fir_filter/n721 ) );
  INV3 U1174 ( .A(\u_decoder/fir_filter/n1149 ), .Q(n2202) );
  NOR31 U1175 ( .A(n1017), .B(\u_cdr/phd1/n9 ), .C(n998), .Q(n1000) );
  NOR31 U1176 ( .A(n1017), .B(\u_cdr/phd1/n9 ), .C(n1051), .Q(n993) );
  NOR21 U1177 ( .A(n913), .B(\u_decoder/fir_filter/n1149 ), .Q(
        \u_decoder/fir_filter/n554 ) );
  INV3 U1178 ( .A(\u_coder/n194 ), .Q(n1719) );
  NAND22 U1179 ( .A(\u_coder/n225 ), .B(n1753), .Q(\u_coder/n241 ) );
  INV3 U1180 ( .A(\u_coder/n262 ), .Q(n1753) );
  NOR21 U1181 ( .A(\u_coder/n162 ), .B(\u_coder/n176 ), .Q(\u_coder/n188 ) );
  NOR21 U1182 ( .A(n982), .B(n1748), .Q(\u_coder/n254 ) );
  NOR21 U1183 ( .A(\u_coder/n315 ), .B(n1769), .Q(\u_coder/N510 ) );
  INV3 U1184 ( .A(\u_coder/N465 ), .Q(n1769) );
  NOR21 U1185 ( .A(n814), .B(n1768), .Q(\u_coder/N511 ) );
  INV3 U1186 ( .A(\u_coder/N466 ), .Q(n1768) );
  INV3 U1187 ( .A(\u_cordic/mycordic/n368 ), .Q(n1310) );
  AOI221 U1188 ( .A(\u_cordic/mycordic/N386 ), .B(n832), .C(
        \u_cordic/mycordic/N418 ), .D(n1582), .Q(\u_cordic/mycordic/n368 ) );
  INV3 U1189 ( .A(\u_cordic/mycordic/n550 ), .Q(n1286) );
  AOI221 U1190 ( .A(\u_cordic/mycordic/N394 ), .B(n831), .C(
        \u_cordic/mycordic/N426 ), .D(n1582), .Q(\u_cordic/mycordic/n550 ) );
  INV3 U1191 ( .A(\u_cordic/mycordic/n551 ), .Q(n1285) );
  AOI221 U1192 ( .A(\u_cordic/mycordic/N393 ), .B(n831), .C(
        \u_cordic/mycordic/N425 ), .D(n1582), .Q(\u_cordic/mycordic/n551 ) );
  INV3 U1193 ( .A(\u_cordic/mycordic/n376 ), .Q(n1217) );
  AOI221 U1194 ( .A(\u_cordic/mycordic/N322 ), .B(n834), .C(
        \u_cordic/mycordic/N354 ), .D(n1578), .Q(\u_cordic/mycordic/n376 ) );
  INV3 U1195 ( .A(\u_cordic/mycordic/n338 ), .Q(n1224) );
  AOI221 U1196 ( .A(\u_cordic/mycordic/N329 ), .B(n834), .C(
        \u_cordic/mycordic/N361 ), .D(n1578), .Q(\u_cordic/mycordic/n338 ) );
  INV3 U1197 ( .A(\u_cordic/mycordic/n337 ), .Q(n1225) );
  AOI221 U1198 ( .A(\u_cordic/mycordic/N330 ), .B(n834), .C(
        \u_cordic/mycordic/N362 ), .D(n1578), .Q(\u_cordic/mycordic/n337 ) );
  INV3 U1199 ( .A(\u_cordic/mycordic/n365 ), .Q(n1280) );
  AOI221 U1200 ( .A(\u_cordic/mycordic/N445 ), .B(n836), .C(
        \u_cordic/mycordic/N473 ), .D(n1581), .Q(\u_cordic/mycordic/n365 ) );
  INV3 U1201 ( .A(\u_cordic/mycordic/n364 ), .Q(n1281) );
  AOI221 U1202 ( .A(\u_cordic/mycordic/N446 ), .B(n836), .C(
        \u_cordic/mycordic/N474 ), .D(n1581), .Q(\u_cordic/mycordic/n364 ) );
  INV3 U1203 ( .A(\u_cordic/mycordic/n542 ), .Q(n1260) );
  AOI221 U1204 ( .A(\u_cordic/mycordic/N453 ), .B(n835), .C(
        \u_cordic/mycordic/N481 ), .D(n1581), .Q(\u_cordic/mycordic/n542 ) );
  INV3 U1205 ( .A(\u_cordic/mycordic/n541 ), .Q(n1261) );
  AOI221 U1206 ( .A(\u_cordic/mycordic/N454 ), .B(n835), .C(
        \u_cordic/mycordic/N482 ), .D(n1581), .Q(\u_cordic/mycordic/n541 ) );
  INV3 U1207 ( .A(\u_cordic/my_rotation/n78 ), .Q(n1522) );
  NAND22 U1208 ( .A(\u_cordic/my_rotation/next_delta [6]), .B(n974), .Q(
        \u_cordic/my_rotation/n78 ) );
  INV3 U1209 ( .A(\u_cordic/my_rotation/n77 ), .Q(n1521) );
  NAND22 U1210 ( .A(\u_cordic/my_rotation/next_delta [7]), .B(n974), .Q(
        \u_cordic/my_rotation/n77 ) );
  NAND22 U1211 ( .A(\u_outFIFO/n495 ), .B(\u_outFIFO/N178 ), .Q(
        \u_outFIFO/n435 ) );
  NAND22 U1212 ( .A(\u_outFIFO/n426 ), .B(\u_outFIFO/N178 ), .Q(
        \u_outFIFO/n366 ) );
  NAND22 U1213 ( .A(\u_outFIFO/n357 ), .B(\u_outFIFO/N178 ), .Q(
        \u_outFIFO/n297 ) );
  NAND22 U1214 ( .A(\u_outFIFO/N178 ), .B(\u_outFIFO/n285 ), .Q(
        \u_outFIFO/n218 ) );
  NOR40 U1215 ( .A(n2315), .B(n1796), .C(n2314), .D(n1793), .Q(
        \u_outFIFO/N474 ) );
  INV3 U1216 ( .A(n2313), .Q(n1793) );
  INV3 U1217 ( .A(n2312), .Q(n1796) );
  NAND22 U1218 ( .A(n1792), .B(n2311), .Q(n2315) );
  NOR21 U1219 ( .A(n983), .B(\u_outFIFO/n511 ), .Q(\u_outFIFO/n215 ) );
  AOI211 U1220 ( .A(\u_coder/n212 ), .B(\u_coder/n211 ), .C(n1710), .Q(
        \u_coder/n201 ) );
  INV3 U1221 ( .A(\u_coder/n209 ), .Q(n1710) );
  NOR21 U1222 ( .A(\u_coder/n178 ), .B(\u_coder/n275 ), .Q(\u_coder/n196 ) );
  NOR31 U1223 ( .A(n777), .B(n776), .C(n1751), .Q(\u_coder/n225 ) );
  NAND22 U1224 ( .A(n978), .B(\u_inFIFO/n200 ), .Q(\u_inFIFO/n119 ) );
  INV3 U1225 ( .A(\u_outFIFO/n529 ), .Q(n1467) );
  NAND22 U1226 ( .A(\u_outFIFO/n512 ), .B(\u_outFIFO/n530 ), .Q(
        \u_outFIFO/n529 ) );
  INV3 U1227 ( .A(\u_coder/n239 ), .Q(n1750) );
  AOI221 U1228 ( .A(\u_coder/n211 ), .B(\u_coder/n212 ), .C(n1711), .D(
        \u_coder/n219 ), .Q(\u_coder/n221 ) );
  AOI221 U1229 ( .A(\u_coder/n211 ), .B(\u_coder/n212 ), .C(n1711), .D(n1751), 
        .Q(\u_coder/n210 ) );
  AOI211 U1230 ( .A(\u_outFIFO/N474 ), .B(\u_outFIFO/n540 ), .C(
        \u_outFIFO/n545 ), .Q(\u_outFIFO/n543 ) );
  OAI311 U1231 ( .A(\u_outFIFO/n546 ), .B(\u_outFIFO/n547 ), .C(
        \u_outFIFO/n534 ), .D(n1789), .Q(\u_outFIFO/n545 ) );
  XNR21 U1232 ( .A(\u_outFIFO/sig_fsm_start_W ), .B(
        \u_outFIFO/sig_fsm_start_R ), .Q(\u_outFIFO/n547 ) );
  AOI211 U1233 ( .A(\u_coder/n162 ), .B(\u_coder/n173 ), .C(\u_coder/n174 ), 
        .Q(\u_coder/n172 ) );
  INV3 U1234 ( .A(\u_coder/n177 ), .Q(n1715) );
  AOI211 U1235 ( .A(\u_coder/n162 ), .B(\u_coder/n163 ), .C(\u_coder/n164 ), 
        .Q(\u_coder/n160 ) );
  NAND22 U1236 ( .A(\u_coder/n209 ), .B(\u_coder/n240 ), .Q(\u_coder/n233 ) );
  NAND22 U1237 ( .A(\u_coder/n266 ), .B(n1724), .Q(\u_coder/n310 ) );
  NOR21 U1238 ( .A(n229), .B(n30), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[7][4] ) );
  NOR21 U1239 ( .A(n230), .B(n31), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[7][4] ) );
  NAND22 U1240 ( .A(\u_coder/n247 ), .B(n1756), .Q(\u_coder/n309 ) );
  NOR21 U1241 ( .A(\u_outFIFO/n205 ), .B(\u_outFIFO/n538 ), .Q(
        \u_outFIFO/n511 ) );
  INV3 U1242 ( .A(\u_coder/n208 ), .Q(n1751) );
  INV3 U1243 ( .A(\u_coder/n176 ), .Q(n1708) );
  NOR21 U1244 ( .A(n814), .B(n1770), .Q(\u_coder/N509 ) );
  INV3 U1245 ( .A(\u_coder/N464 ), .Q(n1770) );
  INV3 U1246 ( .A(\u_cordic/mycordic/n369 ), .Q(n1309) );
  AOI221 U1247 ( .A(\u_cordic/mycordic/N385 ), .B(n832), .C(
        \u_cordic/mycordic/N417 ), .D(n1582), .Q(\u_cordic/mycordic/n369 ) );
  INV3 U1248 ( .A(\u_cordic/mycordic/n370 ), .Q(n1308) );
  AOI221 U1249 ( .A(\u_cordic/mycordic/N384 ), .B(n832), .C(
        \u_cordic/mycordic/N416 ), .D(n1582), .Q(\u_cordic/mycordic/n370 ) );
  INV3 U1250 ( .A(\u_cordic/mycordic/n552 ), .Q(n1284) );
  AOI221 U1251 ( .A(\u_cordic/mycordic/N392 ), .B(n831), .C(
        \u_cordic/mycordic/N424 ), .D(n1582), .Q(\u_cordic/mycordic/n552 ) );
  INV3 U1252 ( .A(\u_cordic/mycordic/n378 ), .Q(n1215) );
  AOI221 U1253 ( .A(\u_cordic/mycordic/N320 ), .B(n834), .C(
        \u_cordic/mycordic/N352 ), .D(n1578), .Q(\u_cordic/mycordic/n378 ) );
  INV3 U1254 ( .A(\u_cordic/mycordic/n377 ), .Q(n1216) );
  AOI221 U1255 ( .A(\u_cordic/mycordic/N321 ), .B(n834), .C(
        \u_cordic/mycordic/N353 ), .D(n1578), .Q(\u_cordic/mycordic/n377 ) );
  INV3 U1256 ( .A(\u_cordic/mycordic/n339 ), .Q(n1223) );
  AOI221 U1257 ( .A(\u_cordic/mycordic/N328 ), .B(n834), .C(
        \u_cordic/mycordic/N360 ), .D(n1578), .Q(\u_cordic/mycordic/n339 ) );
  INV3 U1258 ( .A(\u_decoder/iq_demod/n52 ), .Q(n1935) );
  AOI221 U1259 ( .A(\u_decoder/iq_demod/add_Q_out [2]), .B(n790), .C(n761), 
        .D(n752), .Q(\u_decoder/iq_demod/n52 ) );
  INV3 U1260 ( .A(\u_decoder/iq_demod/n44 ), .Q(n1864) );
  AOI221 U1261 ( .A(\u_decoder/iq_demod/add_I_out [2]), .B(n790), .C(n771), 
        .D(n753), .Q(\u_decoder/iq_demod/n44 ) );
  INV3 U1262 ( .A(\u_cordic/mycordic/n366 ), .Q(n1279) );
  AOI221 U1263 ( .A(\u_cordic/mycordic/N444 ), .B(n836), .C(
        \u_cordic/mycordic/N472 ), .D(n1581), .Q(\u_cordic/mycordic/n366 ) );
  INV3 U1264 ( .A(\u_cordic/mycordic/n543 ), .Q(n1259) );
  AOI221 U1265 ( .A(\u_cordic/mycordic/N452 ), .B(n835), .C(
        \u_cordic/mycordic/N480 ), .D(n1581), .Q(\u_cordic/mycordic/n543 ) );
  INV3 U1266 ( .A(\u_cordic/my_rotation/n79 ), .Q(n1523) );
  NAND22 U1267 ( .A(\u_cordic/my_rotation/next_delta [5]), .B(n974), .Q(
        \u_cordic/my_rotation/n79 ) );
  NOR31 U1268 ( .A(\u_inFIFO/n223 ), .B(n984), .C(\u_inFIFO/n224 ), .Q(
        \u_inFIFO/n212 ) );
  NAND22 U1269 ( .A(\u_cordic/n29 ), .B(n1777), .Q(\u_cordic/n21 ) );
  NAND31 U1270 ( .A(n295), .B(n36), .C(n1657), .Q(\u_cdr/n29 ) );
  NAND22 U1271 ( .A(n978), .B(n2689), .Q(\u_cdr/n43 ) );
  NOR21 U1272 ( .A(n982), .B(\u_outFIFO/n209 ), .Q(\u_outFIFO/n208 ) );
  OAI2111 U1273 ( .A(n2226), .B(n2227), .C(n2228), .D(n2229), .Q(n2591) );
  INV3 U1274 ( .A(\u_coder/n161 ), .Q(n1724) );
  INV3 U1275 ( .A(n216), .Q(n964) );
  INV3 U1276 ( .A(n215), .Q(n942) );
  NAND31 U1277 ( .A(\u_inFIFO/n224 ), .B(\u_inFIFO/n200 ), .C(\u_inFIFO/n202 ), 
        .Q(\u_inFIFO/n226 ) );
  INV3 U1278 ( .A(\u_inFIFO/n224 ), .Q(n1702) );
  INV3 U1279 ( .A(\u_outFIFO/n526 ), .Q(n1466) );
  NOR21 U1280 ( .A(\u_outFIFO/n527 ), .B(\u_outFIFO/n514 ), .Q(
        \u_outFIFO/n526 ) );
  INV3 U1281 ( .A(\u_outFIFO/n530 ), .Q(n1468) );
  NAND22 U1282 ( .A(n1697), .B(n973), .Q(\u_inFIFO/n225 ) );
  INV3 U1283 ( .A(\u_inFIFO/n200 ), .Q(n1697) );
  NAND22 U1284 ( .A(\u_inFIFO/n226 ), .B(\u_inFIFO/n227 ), .Q(\u_inFIFO/n223 )
         );
  NOR21 U1285 ( .A(n229), .B(n37), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[7][5] ) );
  NOR21 U1286 ( .A(n230), .B(n38), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[7][5] ) );
  NOR21 U1287 ( .A(n2282), .B(\u_coder/n161 ), .Q(\u_coder/n286 ) );
  INV3 U1288 ( .A(\u_coder/n200 ), .Q(n1756) );
  XOR21 U1289 ( .A(n1786), .B(\u_cdr/dp_cluster_0/mult_add_59_aco/PROD_not[0] ), .Q(n358) );
  XNR21 U1290 ( .A(\u_cdr/dp_cluster_0/mult_add_59_aco/PROD_not[2] ), .B(
        \u_cdr/n48 ), .Q(n359) );
  XNR21 U1291 ( .A(n1784), .B(\u_cdr/n47 ), .Q(\u_cdr/n45 ) );
  INV3 U1292 ( .A(\u_cdr/dp_cluster_0/mult_add_59_aco/PROD_not[3] ), .Q(n1784)
         );
  NOR21 U1293 ( .A(\u_cdr/n48 ), .B(
        \u_cdr/dp_cluster_0/mult_add_59_aco/PROD_not[2] ), .Q(\u_cdr/n47 ) );
  NAND22 U1294 ( .A(\u_coder/n280 ), .B(n776), .Q(\u_coder/n259 ) );
  NAND22 U1295 ( .A(n1786), .B(n1785), .Q(\u_cdr/n48 ) );
  INV3 U1296 ( .A(n2275), .Q(n1746) );
  OAI311 U1297 ( .A(n294), .B(\u_cdr/n29 ), .C(n3), .D(n978), .Q(\u_cdr/n44 )
         );
  NAND22 U1298 ( .A(n1657), .B(\u_cdr/n42 ), .Q(\u_cdr/n38 ) );
  BUF6 U1299 ( .A(n805), .Q(n944) );
  BUF6 U1300 ( .A(n805), .Q(n945) );
  BUF6 U1301 ( .A(n805), .Q(n946) );
  INV3 U1302 ( .A(n2689), .Q(n1657) );
  INV3 U1303 ( .A(n2282), .Q(n1716) );
  INV3 U1304 ( .A(\u_coder/n165 ), .Q(n1720) );
  BUF2 U1305 ( .A(n805), .Q(n947) );
  BUF2 U1306 ( .A(n166), .Q(n781) );
  INV3 U1307 ( .A(\u_cdr/dp_cluster_0/mult_add_59_aco/PROD_not[0] ), .Q(n1785)
         );
  INV3 U1308 ( .A(\u_coder/n240 ), .Q(n1711) );
  INV3 U1309 ( .A(\u_cordic/n29 ), .Q(n1778) );
  INV3 U1310 ( .A(\u_inFIFO/n192 ), .Q(n1620) );
  NOR21 U1311 ( .A(\u_inFIFO/n142 ), .B(\u_inFIFO/n179 ), .Q(\u_inFIFO/n193 )
         );
  INV3 U1312 ( .A(\u_inFIFO/n190 ), .Q(n1621) );
  NOR21 U1313 ( .A(\u_inFIFO/n139 ), .B(\u_inFIFO/n179 ), .Q(\u_inFIFO/n191 )
         );
  INV3 U1314 ( .A(\u_inFIFO/n188 ), .Q(n1622) );
  NOR21 U1315 ( .A(\u_inFIFO/n136 ), .B(\u_inFIFO/n179 ), .Q(\u_inFIFO/n189 )
         );
  INV3 U1316 ( .A(\u_inFIFO/n186 ), .Q(n1623) );
  NOR21 U1317 ( .A(\u_inFIFO/n133 ), .B(\u_inFIFO/n179 ), .Q(\u_inFIFO/n187 )
         );
  INV3 U1318 ( .A(\u_inFIFO/n184 ), .Q(n1624) );
  NOR21 U1319 ( .A(\u_inFIFO/n130 ), .B(\u_inFIFO/n179 ), .Q(\u_inFIFO/n185 )
         );
  INV3 U1320 ( .A(\u_inFIFO/n182 ), .Q(n1625) );
  NOR21 U1321 ( .A(\u_inFIFO/n127 ), .B(\u_inFIFO/n179 ), .Q(\u_inFIFO/n183 )
         );
  INV3 U1322 ( .A(\u_inFIFO/n180 ), .Q(n1626) );
  NOR21 U1323 ( .A(\u_inFIFO/n124 ), .B(\u_inFIFO/n179 ), .Q(\u_inFIFO/n181 )
         );
  INV3 U1324 ( .A(\u_inFIFO/n177 ), .Q(n1627) );
  NOR21 U1325 ( .A(\u_inFIFO/n120 ), .B(\u_inFIFO/n179 ), .Q(\u_inFIFO/n178 )
         );
  INV3 U1326 ( .A(\u_inFIFO/n175 ), .Q(n1628) );
  NOR21 U1327 ( .A(\u_inFIFO/n142 ), .B(\u_inFIFO/n162 ), .Q(\u_inFIFO/n176 )
         );
  INV3 U1328 ( .A(\u_inFIFO/n173 ), .Q(n1629) );
  NOR21 U1329 ( .A(\u_inFIFO/n139 ), .B(\u_inFIFO/n162 ), .Q(\u_inFIFO/n174 )
         );
  INV3 U1330 ( .A(\u_inFIFO/n171 ), .Q(n1630) );
  NOR21 U1331 ( .A(\u_inFIFO/n136 ), .B(\u_inFIFO/n162 ), .Q(\u_inFIFO/n172 )
         );
  INV3 U1332 ( .A(\u_inFIFO/n169 ), .Q(n1631) );
  NOR21 U1333 ( .A(\u_inFIFO/n133 ), .B(\u_inFIFO/n162 ), .Q(\u_inFIFO/n170 )
         );
  INV3 U1334 ( .A(\u_inFIFO/n167 ), .Q(n1632) );
  NOR21 U1335 ( .A(\u_inFIFO/n130 ), .B(\u_inFIFO/n162 ), .Q(\u_inFIFO/n168 )
         );
  INV3 U1336 ( .A(\u_inFIFO/n165 ), .Q(n1633) );
  NOR21 U1337 ( .A(\u_inFIFO/n127 ), .B(\u_inFIFO/n162 ), .Q(\u_inFIFO/n166 )
         );
  INV3 U1338 ( .A(\u_inFIFO/n163 ), .Q(n1634) );
  NOR21 U1339 ( .A(\u_inFIFO/n124 ), .B(\u_inFIFO/n162 ), .Q(\u_inFIFO/n164 )
         );
  INV3 U1340 ( .A(\u_inFIFO/n160 ), .Q(n1635) );
  NOR21 U1341 ( .A(\u_inFIFO/n120 ), .B(\u_inFIFO/n162 ), .Q(\u_inFIFO/n161 )
         );
  INV3 U1342 ( .A(\u_inFIFO/n158 ), .Q(n1636) );
  NOR21 U1343 ( .A(\u_inFIFO/n142 ), .B(\u_inFIFO/n145 ), .Q(\u_inFIFO/n159 )
         );
  INV3 U1344 ( .A(\u_inFIFO/n156 ), .Q(n1637) );
  NOR21 U1345 ( .A(\u_inFIFO/n139 ), .B(\u_inFIFO/n145 ), .Q(\u_inFIFO/n157 )
         );
  INV3 U1346 ( .A(\u_inFIFO/n154 ), .Q(n1638) );
  NOR21 U1347 ( .A(\u_inFIFO/n136 ), .B(\u_inFIFO/n145 ), .Q(\u_inFIFO/n155 )
         );
  INV3 U1348 ( .A(\u_inFIFO/n152 ), .Q(n1639) );
  NOR21 U1349 ( .A(\u_inFIFO/n133 ), .B(\u_inFIFO/n145 ), .Q(\u_inFIFO/n153 )
         );
  INV3 U1350 ( .A(\u_inFIFO/n150 ), .Q(n1640) );
  NOR21 U1351 ( .A(\u_inFIFO/n130 ), .B(\u_inFIFO/n145 ), .Q(\u_inFIFO/n151 )
         );
  INV3 U1352 ( .A(\u_inFIFO/n148 ), .Q(n1641) );
  NOR21 U1353 ( .A(\u_inFIFO/n127 ), .B(\u_inFIFO/n145 ), .Q(\u_inFIFO/n149 )
         );
  INV3 U1354 ( .A(\u_inFIFO/n146 ), .Q(n1642) );
  NOR21 U1355 ( .A(\u_inFIFO/n124 ), .B(\u_inFIFO/n145 ), .Q(\u_inFIFO/n147 )
         );
  INV3 U1356 ( .A(\u_inFIFO/n143 ), .Q(n1643) );
  NOR21 U1357 ( .A(\u_inFIFO/n120 ), .B(\u_inFIFO/n145 ), .Q(\u_inFIFO/n144 )
         );
  INV3 U1358 ( .A(\u_inFIFO/n140 ), .Q(n1644) );
  NOR21 U1359 ( .A(\u_inFIFO/n121 ), .B(\u_inFIFO/n142 ), .Q(\u_inFIFO/n141 )
         );
  INV3 U1360 ( .A(\u_inFIFO/n137 ), .Q(n1645) );
  NOR21 U1361 ( .A(\u_inFIFO/n121 ), .B(\u_inFIFO/n139 ), .Q(\u_inFIFO/n138 )
         );
  INV3 U1362 ( .A(\u_inFIFO/n134 ), .Q(n1646) );
  NOR21 U1363 ( .A(\u_inFIFO/n121 ), .B(\u_inFIFO/n136 ), .Q(\u_inFIFO/n135 )
         );
  INV3 U1364 ( .A(\u_inFIFO/n131 ), .Q(n1647) );
  NOR21 U1365 ( .A(\u_inFIFO/n121 ), .B(\u_inFIFO/n133 ), .Q(\u_inFIFO/n132 )
         );
  INV3 U1366 ( .A(\u_inFIFO/n128 ), .Q(n1648) );
  NOR21 U1367 ( .A(\u_inFIFO/n121 ), .B(\u_inFIFO/n130 ), .Q(\u_inFIFO/n129 )
         );
  INV3 U1368 ( .A(\u_inFIFO/n125 ), .Q(n1649) );
  NOR21 U1369 ( .A(\u_inFIFO/n121 ), .B(\u_inFIFO/n127 ), .Q(\u_inFIFO/n126 )
         );
  INV3 U1370 ( .A(\u_inFIFO/n122 ), .Q(n1650) );
  NOR21 U1371 ( .A(\u_inFIFO/n121 ), .B(\u_inFIFO/n124 ), .Q(\u_inFIFO/n123 )
         );
  INV3 U1372 ( .A(\u_coder/n251 ), .Q(n1655) );
  NAND22 U1373 ( .A(n1749), .B(\u_coder/n212 ), .Q(\u_coder/n251 ) );
  INV3 U1374 ( .A(\u_inFIFO/n112 ), .Q(n1651) );
  NOR21 U1375 ( .A(\u_inFIFO/n120 ), .B(\u_inFIFO/n121 ), .Q(\u_inFIFO/n117 )
         );
  INV3 U1376 ( .A(\u_coder/n260 ), .Q(n1712) );
  NOR21 U1377 ( .A(\u_coder/n261 ), .B(\u_coder/n161 ), .Q(\u_coder/n260 ) );
  INV3 U1378 ( .A(\u_coder/n270 ), .Q(n1653) );
  NAND22 U1379 ( .A(\u_coder/n196 ), .B(\u_coder/n195 ), .Q(\u_coder/n270 ) );
  NOR21 U1380 ( .A(n229), .B(\u_decoder/I_prefilter [6]), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r164/CARRYB[7][3] ) );
  NOR21 U1381 ( .A(n230), .B(\u_decoder/Q_prefilter [6]), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r177/CARRYB[7][3] ) );
  NOR21 U1382 ( .A(n229), .B(\u_decoder/I_prefilter [6]), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r165/CARRYB[7][4] ) );
  NOR21 U1383 ( .A(n230), .B(\u_decoder/Q_prefilter [6]), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r178/CARRYB[7][4] ) );
  INV3 U1384 ( .A(\u_coder/n258 ), .Q(n1725) );
  NOR21 U1385 ( .A(\u_coder/n259 ), .B(\u_coder/n200 ), .Q(\u_coder/n258 ) );
  INV3 U1386 ( .A(\u_inFIFO/n204 ), .Q(n1478) );
  AOI221 U1387 ( .A(\u_inFIFO/n202 ), .B(n780), .C(\u_inFIFO/n203 ), .D(
        \u_inFIFO/N120 ), .Q(\u_inFIFO/n204 ) );
  INV3 U1388 ( .A(\u_outFIFO/n506 ), .Q(n1330) );
  AOI221 U1389 ( .A(\u_outFIFO/n504 ), .B(n775), .C(\u_outFIFO/n505 ), .D(
        \u_outFIFO/N198 ), .Q(\u_outFIFO/n506 ) );
  INV3 U1390 ( .A(\u_cordic/mycordic/n347 ), .Q(n1235) );
  AOI221 U1391 ( .A(n1579), .B(\u_cordic/mycordic/N257 ), .C(n787), .D(
        \u_cordic/mycordic/N265 ), .Q(\u_cordic/mycordic/n347 ) );
  INV3 U1392 ( .A(\u_cordic/mycordic/n346 ), .Q(n1236) );
  AOI221 U1393 ( .A(n1579), .B(\u_cordic/mycordic/N258 ), .C(n787), .D(
        \u_cordic/mycordic/N266 ), .Q(\u_cordic/mycordic/n346 ) );
  INV3 U1394 ( .A(\u_cordic/mycordic/n385 ), .Q(n1230) );
  AOI221 U1395 ( .A(n1579), .B(\u_cordic/mycordic/N289 ), .C(n787), .D(
        \u_cordic/mycordic/N257 ), .Q(\u_cordic/mycordic/n385 ) );
  INV3 U1396 ( .A(\u_cordic/mycordic/n384 ), .Q(n1231) );
  AOI221 U1397 ( .A(n1579), .B(\u_cordic/mycordic/N290 ), .C(n787), .D(
        \u_cordic/mycordic/N258 ), .Q(\u_cordic/mycordic/n384 ) );
  NOR21 U1398 ( .A(\u_coder/n315 ), .B(n1771), .Q(\u_coder/N508 ) );
  INV3 U1399 ( .A(\u_coder/N463 ), .Q(n1771) );
  NOR21 U1400 ( .A(n814), .B(n1772), .Q(\u_coder/N507 ) );
  INV3 U1401 ( .A(\u_coder/N462 ), .Q(n1772) );
  INV3 U1402 ( .A(\u_cordic/mycordic/n331 ), .Q(n1314) );
  AOI221 U1403 ( .A(\u_cordic/mycordic/N390 ), .B(n832), .C(
        \u_cordic/mycordic/N422 ), .D(n1582), .Q(\u_cordic/mycordic/n331 ) );
  INV3 U1404 ( .A(\u_cordic/mycordic/n371 ), .Q(n1307) );
  AOI221 U1405 ( .A(\u_cordic/mycordic/N383 ), .B(n832), .C(
        \u_cordic/mycordic/N415 ), .D(n1582), .Q(\u_cordic/mycordic/n371 ) );
  INV3 U1406 ( .A(\u_cordic/mycordic/n372 ), .Q(n1306) );
  AOI221 U1407 ( .A(\u_cordic/mycordic/N382 ), .B(n832), .C(
        \u_cordic/mycordic/N414 ), .D(n1582), .Q(\u_cordic/mycordic/n372 ) );
  INV3 U1408 ( .A(\u_cordic/mycordic/n553 ), .Q(n1283) );
  AOI221 U1409 ( .A(\u_cordic/mycordic/N391 ), .B(n831), .C(
        \u_cordic/mycordic/N423 ), .D(n1582), .Q(\u_cordic/mycordic/n553 ) );
  INV3 U1410 ( .A(\u_cordic/mycordic/n380 ), .Q(n1213) );
  AOI221 U1411 ( .A(\u_cordic/mycordic/N318 ), .B(n834), .C(
        \u_cordic/mycordic/N350 ), .D(n1578), .Q(\u_cordic/mycordic/n380 ) );
  INV3 U1412 ( .A(\u_cordic/mycordic/n379 ), .Q(n1214) );
  AOI221 U1413 ( .A(\u_cordic/mycordic/N319 ), .B(n834), .C(
        \u_cordic/mycordic/N351 ), .D(n1578), .Q(\u_cordic/mycordic/n379 ) );
  INV3 U1414 ( .A(\u_cordic/mycordic/n341 ), .Q(n1221) );
  AOI221 U1415 ( .A(\u_cordic/mycordic/N326 ), .B(n834), .C(
        \u_cordic/mycordic/N358 ), .D(n1578), .Q(\u_cordic/mycordic/n341 ) );
  INV3 U1416 ( .A(\u_cordic/mycordic/n340 ), .Q(n1222) );
  AOI221 U1417 ( .A(\u_cordic/mycordic/N327 ), .B(n834), .C(
        \u_cordic/mycordic/N359 ), .D(n1578), .Q(\u_cordic/mycordic/n340 ) );
  INV3 U1418 ( .A(\u_decoder/iq_demod/n51 ), .Q(n1933) );
  AOI221 U1419 ( .A(\u_decoder/iq_demod/add_Q_out [1]), .B(n790), .C(
        \u_decoder/Q_prefilter [1]), .D(n752), .Q(\u_decoder/iq_demod/n51 ) );
  INV3 U1420 ( .A(\u_decoder/iq_demod/n43 ), .Q(n1862) );
  AOI221 U1421 ( .A(\u_decoder/iq_demod/add_I_out [1]), .B(n790), .C(
        \u_decoder/I_prefilter [1]), .D(n753), .Q(\u_decoder/iq_demod/n43 ) );
  INV3 U1422 ( .A(\u_cordic/mycordic/n545 ), .Q(n1257) );
  AOI221 U1423 ( .A(\u_cordic/mycordic/N450 ), .B(n835), .C(
        \u_cordic/mycordic/N478 ), .D(n1581), .Q(\u_cordic/mycordic/n545 ) );
  INV3 U1424 ( .A(\u_cordic/mycordic/n544 ), .Q(n1258) );
  AOI221 U1425 ( .A(\u_cordic/mycordic/N451 ), .B(n835), .C(
        \u_cordic/mycordic/N479 ), .D(n1581), .Q(\u_cordic/mycordic/n544 ) );
  INV3 U1426 ( .A(\u_cordic/my_rotation/n80 ), .Q(n1524) );
  NAND22 U1427 ( .A(\u_cordic/my_rotation/next_delta [4]), .B(n974), .Q(
        \u_cordic/my_rotation/n80 ) );
  NAND22 U1428 ( .A(\u_outFIFO/n495 ), .B(\u_outFIFO/n288 ), .Q(
        \u_outFIFO/n438 ) );
  NAND22 U1429 ( .A(\u_outFIFO/n426 ), .B(\u_outFIFO/n288 ), .Q(
        \u_outFIFO/n369 ) );
  NAND22 U1430 ( .A(\u_outFIFO/n357 ), .B(\u_outFIFO/n288 ), .Q(
        \u_outFIFO/n300 ) );
  NAND22 U1431 ( .A(\u_outFIFO/n495 ), .B(\u_outFIFO/n291 ), .Q(
        \u_outFIFO/n441 ) );
  NAND22 U1432 ( .A(\u_outFIFO/n426 ), .B(\u_outFIFO/n291 ), .Q(
        \u_outFIFO/n372 ) );
  NAND22 U1433 ( .A(\u_outFIFO/n357 ), .B(\u_outFIFO/n291 ), .Q(
        \u_outFIFO/n303 ) );
  NAND22 U1434 ( .A(\u_outFIFO/n495 ), .B(\u_outFIFO/n294 ), .Q(
        \u_outFIFO/n444 ) );
  NAND22 U1435 ( .A(\u_outFIFO/n426 ), .B(\u_outFIFO/n294 ), .Q(
        \u_outFIFO/n375 ) );
  NAND22 U1436 ( .A(\u_outFIFO/n357 ), .B(\u_outFIFO/n294 ), .Q(
        \u_outFIFO/n306 ) );
  NAND22 U1437 ( .A(\u_outFIFO/n294 ), .B(\u_outFIFO/n285 ), .Q(
        \u_outFIFO/n227 ) );
  NAND22 U1438 ( .A(\u_outFIFO/n291 ), .B(\u_outFIFO/n285 ), .Q(
        \u_outFIFO/n224 ) );
  NAND22 U1439 ( .A(\u_outFIFO/n288 ), .B(\u_outFIFO/n285 ), .Q(
        \u_outFIFO/n221 ) );
  NOR21 U1440 ( .A(n982), .B(\u_outFIFO/n206 ), .Q(\u_outFIFO/n504 ) );
  NAND22 U1441 ( .A(\u_inFIFO/n109 ), .B(\u_inFIFO/n106 ), .Q(\u_inFIFO/n209 )
         );
  NOR21 U1442 ( .A(\u_cdr/n37 ), .B(n984), .Q(\u_cdr/n32 ) );
  NOR21 U1443 ( .A(n982), .B(\u_outFIFO/n504 ), .Q(\u_outFIFO/n505 ) );
  NAND22 U1444 ( .A(\u_decoder/iq_demod/cossin_dig/n37 ), .B(
        \u_decoder/iq_demod/cossin_dig/n26 ), .Q(
        \u_decoder/iq_demod/cossin_dig/n31 ) );
  NOR40 U1445 ( .A(n2229), .B(n2228), .C(n2227), .D(n2226), .Q(
        \u_cordic/my_rotation/n89 ) );
  INV3 U1446 ( .A(\u_cordic/mycordic/n386 ), .Q(n1229) );
  AOI221 U1447 ( .A(n1579), .B(\u_cordic/mycordic/N288 ), .C(n787), .D(
        \u_cordic/mycordic/N256 ), .Q(\u_cordic/mycordic/n386 ) );
  NAND22 U1448 ( .A(n976), .B(\u_decoder/iq_demod/cossin_dig/n26 ), .Q(
        \u_decoder/iq_demod/cossin_dig/n42 ) );
  NAND22 U1449 ( .A(n1698), .B(\u_inFIFO/n106 ), .Q(\u_inFIFO/n237 ) );
  NAND22 U1450 ( .A(\u_outFIFO/n206 ), .B(n969), .Q(\u_outFIFO/n525 ) );
  NOR21 U1451 ( .A(\u_coder/n315 ), .B(n1776), .Q(\u_coder/N504 ) );
  INV3 U1452 ( .A(\u_coder/N459 ), .Q(n1776) );
  NOR21 U1453 ( .A(n814), .B(n1775), .Q(\u_coder/N505 ) );
  INV3 U1454 ( .A(\u_coder/N460 ), .Q(n1775) );
  NOR21 U1455 ( .A(\u_coder/n315 ), .B(n1774), .Q(\u_coder/N506 ) );
  INV3 U1456 ( .A(\u_coder/N461 ), .Q(n1774) );
  BUF2 U1457 ( .A(\u_cordic/mycordic/n332 ), .Q(n831) );
  BUF2 U1458 ( .A(\u_cordic/mycordic/n336 ), .Q(n833) );
  INV3 U1459 ( .A(sig_MUX_outMUX8), .Q(n1663) );
  NOR21 U1460 ( .A(\u_coder/n208 ), .B(n776), .Q(\u_coder/n207 ) );
  NOR21 U1461 ( .A(\u_cordic/mycordic/present_Q_table[0][5] ), .B(n548), .Q(
        \u_cordic/mycordic/sub_add_151_b0/carry [6]) );
  INV3 U1462 ( .A(\u_cordic/mycordic/sub_add_151_b0/carry [5]), .Q(n548) );
  NOR21 U1463 ( .A(\u_cordic/mycordic/present_I_table[0][5] ), .B(n546), .Q(
        \u_cordic/mycordic/sub_add_150_b0/carry [6]) );
  INV3 U1464 ( .A(\u_cordic/mycordic/sub_add_150_b0/carry [5]), .Q(n546) );
  NOR21 U1465 ( .A(\u_cordic/mycordic/present_Q_table[0][4] ), .B(
        \u_cordic/mycordic/present_Q_table[0][3] ), .Q(
        \u_cordic/mycordic/sub_add_151_b0/carry [5]) );
  BUF2 U1466 ( .A(n166), .Q(n782) );
  INV3 U1467 ( .A(\u_coder/n314 ), .Q(n1757) );
  NAND22 U1468 ( .A(\u_inFIFO/n236 ), .B(\u_inFIFO/n237 ), .Q(\u_inFIFO/n234 )
         );
  INV3 U1469 ( .A(\u_coder/n220 ), .Q(n1707) );
  INV3 U1470 ( .A(\u_cordic/n18 ), .Q(n1777) );
  INV3 U1471 ( .A(\u_inFIFO/n241 ), .Q(n1698) );
  BUF2 U1472 ( .A(n166), .Q(n783) );
  INV3 U1473 ( .A(\u_coder/n219 ), .Q(n1727) );
  BUF2 U1474 ( .A(\u_outFIFO/n284 ), .Q(n806) );
  BUF2 U1475 ( .A(\u_outFIFO/n275 ), .Q(n803) );
  BUF2 U1476 ( .A(\u_outFIFO/n266 ), .Q(n801) );
  BUF2 U1477 ( .A(\u_outFIFO/n257 ), .Q(n799) );
  BUF2 U1478 ( .A(\u_outFIFO/n230 ), .Q(n793) );
  BUF2 U1479 ( .A(\u_outFIFO/n248 ), .Q(n797) );
  BUF2 U1480 ( .A(\u_outFIFO/n239 ), .Q(n795) );
  BUF2 U1481 ( .A(\u_outFIFO/n284 ), .Q(n807) );
  BUF2 U1482 ( .A(\u_outFIFO/n275 ), .Q(n804) );
  BUF2 U1483 ( .A(\u_outFIFO/n266 ), .Q(n802) );
  BUF2 U1484 ( .A(\u_outFIFO/n257 ), .Q(n800) );
  BUF2 U1485 ( .A(\u_outFIFO/n230 ), .Q(n794) );
  BUF2 U1486 ( .A(\u_outFIFO/n248 ), .Q(n798) );
  BUF2 U1487 ( .A(\u_outFIFO/n239 ), .Q(n796) );
  BUF2 U1488 ( .A(\u_outFIFO/n217 ), .Q(n791) );
  BUF2 U1489 ( .A(\u_outFIFO/n217 ), .Q(n792) );
  INV3 U1490 ( .A(\u_outFIFO/n537 ), .Q(n1789) );
  NOR21 U1491 ( .A(\u_cordic/mycordic/present_Q_table[0][6] ), .B(n549), .Q(
        \u_cordic/mycordic/sub_add_151_b0/carry [7]) );
  INV3 U1492 ( .A(\u_cordic/mycordic/sub_add_151_b0/carry [6]), .Q(n549) );
  INV3 U1493 ( .A(\u_outFIFO/n539 ), .Q(n1788) );
  BUF2 U1494 ( .A(\u_cordic/mycordic/n332 ), .Q(n832) );
  BUF2 U1495 ( .A(\u_cordic/mycordic/n336 ), .Q(n834) );
  INV3 U1496 ( .A(\u_inFIFO/n206 ), .Q(n1476) );
  AOI221 U1497 ( .A(\u_inFIFO/n202 ), .B(\u_inFIFO/N34 ), .C(\u_inFIFO/n203 ), 
        .D(\u_inFIFO/N118 ), .Q(\u_inFIFO/n206 ) );
  INV3 U1498 ( .A(\u_inFIFO/n205 ), .Q(n1477) );
  AOI221 U1499 ( .A(\u_inFIFO/n202 ), .B(n779), .C(\u_inFIFO/n203 ), .D(
        \u_inFIFO/N119 ), .Q(\u_inFIFO/n205 ) );
  NOR21 U1500 ( .A(\u_cordic/mycordic/present_I_table[0][4] ), .B(
        \u_cordic/mycordic/present_I_table[0][3] ), .Q(
        \u_cordic/mycordic/sub_add_150_b0/carry [5]) );
  NAND22 U1501 ( .A(n1506), .B(\u_decoder/iq_demod/cossin_dig/n37 ), .Q(
        \u_decoder/iq_demod/cossin_dig/n40 ) );
  INV3 U1502 ( .A(\u_decoder/iq_demod/cossin_dig/n42 ), .Q(n1506) );
  NOR21 U1503 ( .A(\u_cordic/mycordic/present_I_table[0][6] ), .B(n547), .Q(
        \u_cordic/mycordic/sub_add_150_b0/carry [7]) );
  INV3 U1504 ( .A(\u_cordic/mycordic/sub_add_150_b0/carry [6]), .Q(n547) );
  INV3 U1505 ( .A(\u_outFIFO/n509 ), .Q(n1327) );
  AOI221 U1506 ( .A(\u_outFIFO/n504 ), .B(n35), .C(\u_outFIFO/n505 ), .D(n215), 
        .Q(\u_outFIFO/n509 ) );
  INV3 U1507 ( .A(\u_outFIFO/n508 ), .Q(n1328) );
  AOI221 U1508 ( .A(\u_outFIFO/n504 ), .B(\u_outFIFO/N36 ), .C(
        \u_outFIFO/n505 ), .D(\u_outFIFO/N196 ), .Q(\u_outFIFO/n508 ) );
  INV3 U1509 ( .A(\u_outFIFO/n507 ), .Q(n1329) );
  AOI221 U1510 ( .A(\u_outFIFO/n504 ), .B(n774), .C(\u_outFIFO/n505 ), .D(
        \u_outFIFO/N197 ), .Q(\u_outFIFO/n507 ) );
  INV3 U1511 ( .A(\u_cordic/mycordic/n348 ), .Q(n1234) );
  AOI221 U1512 ( .A(n1579), .B(\u_cordic/mycordic/N256 ), .C(n787), .D(
        \u_cordic/mycordic/N264 ), .Q(\u_cordic/mycordic/n348 ) );
  INV3 U1513 ( .A(\u_cordic/mycordic/n333 ), .Q(n1313) );
  AOI221 U1514 ( .A(\u_cordic/mycordic/N389 ), .B(n832), .C(
        \u_cordic/mycordic/N421 ), .D(n1582), .Q(\u_cordic/mycordic/n333 ) );
  INV3 U1515 ( .A(\u_cordic/mycordic/n373 ), .Q(n1305) );
  AOI221 U1516 ( .A(\u_cordic/mycordic/N381 ), .B(n832), .C(
        \u_cordic/mycordic/N413 ), .D(n1582), .Q(\u_cordic/mycordic/n373 ) );
  INV3 U1517 ( .A(\u_cordic/mycordic/n381 ), .Q(n1212) );
  AOI221 U1518 ( .A(\u_cordic/mycordic/N317 ), .B(n834), .C(
        \u_cordic/mycordic/N349 ), .D(n1578), .Q(\u_cordic/mycordic/n381 ) );
  INV3 U1519 ( .A(\u_cordic/mycordic/n342 ), .Q(n1220) );
  AOI221 U1520 ( .A(\u_cordic/mycordic/N325 ), .B(n834), .C(
        \u_cordic/mycordic/N357 ), .D(n1578), .Q(\u_cordic/mycordic/n342 ) );
  INV3 U1521 ( .A(\u_decoder/iq_demod/n50 ), .Q(n1908) );
  AOI221 U1522 ( .A(\u_decoder/iq_demod/add_Q_out [0]), .B(n790), .C(n763), 
        .D(n753), .Q(\u_decoder/iq_demod/n50 ) );
  XOR21 U1523 ( .A(\u_decoder/iq_demod/dp_cluster_1/mult_I_sin_out [0]), .B(
        \u_decoder/iq_demod/dp_cluster_1/mult_Q_cos_out [0]), .Q(
        \u_decoder/iq_demod/add_Q_out [0]) );
  INV3 U1524 ( .A(\u_decoder/iq_demod/n41 ), .Q(n1837) );
  AOI221 U1525 ( .A(\u_decoder/iq_demod/add_I_out [0]), .B(n790), .C(n753), 
        .D(n773), .Q(\u_decoder/iq_demod/n41 ) );
  XNR21 U1526 ( .A(\u_decoder/iq_demod/dp_cluster_0/mult_I_cos_out [0]), .B(
        n1946), .Q(\u_decoder/iq_demod/add_I_out [0]) );
  INV3 U1527 ( .A(\u_cordic/mycordic/n546 ), .Q(n1256) );
  AOI221 U1528 ( .A(\u_cordic/mycordic/N449 ), .B(n835), .C(
        \u_cordic/mycordic/N477 ), .D(n1581), .Q(\u_cordic/mycordic/n546 ) );
  INV3 U1529 ( .A(\u_cordic/my_rotation/n82 ), .Q(n1526) );
  NAND22 U1530 ( .A(\u_cordic/my_rotation/next_delta [2]), .B(n974), .Q(
        \u_cordic/my_rotation/n82 ) );
  INV3 U1531 ( .A(\u_cordic/my_rotation/n81 ), .Q(n1525) );
  NAND22 U1532 ( .A(\u_cordic/my_rotation/next_delta [3]), .B(n974), .Q(
        \u_cordic/my_rotation/n81 ) );
  INV3 U1533 ( .A(\u_decoder/iq_demod/n70 ), .Q(n1583) );
  NAND22 U1534 ( .A(\u_decoder/iq_demod/n71 ), .B(n969), .Q(
        \u_decoder/iq_demod/n70 ) );
  INV3 U1535 ( .A(n790), .Q(n1961) );
  INV6 U1536 ( .A(\u_cordic/mycordic/n548 ), .Q(n1581) );
  NAND22 U1537 ( .A(n749), .B(n969), .Q(\u_cordic/mycordic/n548 ) );
  NOR21 U1538 ( .A(n985), .B(\u_inFIFO/n202 ), .Q(\u_inFIFO/n203 ) );
  INV3 U1539 ( .A(\u_cordic/mycordic/n349 ), .Q(n1233) );
  AOI221 U1540 ( .A(n1579), .B(\u_cordic/mycordic/N255 ), .C(n787), .D(
        \u_cordic/mycordic/N263 ), .Q(\u_cordic/mycordic/n349 ) );
  NOR21 U1541 ( .A(n983), .B(n749), .Q(\u_cordic/mycordic/n363 ) );
  NOR21 U1542 ( .A(\u_outFIFO/n546 ), .B(\u_outFIFO/n205 ), .Q(
        \u_outFIFO/n540 ) );
  INV3 U1543 ( .A(\u_inFIFO/n227 ), .Q(n1652) );
  INV3 U1544 ( .A(\u_cordic/mycordic/n391 ), .Q(n1575) );
  AOI211 U1545 ( .A(\u_decoder/fir_filter/n1153 ), .B(
        \u_decoder/fir_filter/n1154 ), .C(n980), .Q(\u_decoder/fir_filter/N11 ) );
  NAND22 U1546 ( .A(\u_decoder/fir_filter/n1151 ), .B(n314), .Q(
        \u_decoder/fir_filter/n1154 ) );
  BUF2 U1547 ( .A(\u_cordic/mycordic/n456 ), .Q(n788) );
  BUF2 U1548 ( .A(\u_cordic/mycordic/n456 ), .Q(n789) );
  BUF2 U1549 ( .A(\u_cordic/mycordic/n438 ), .Q(n785) );
  BUF2 U1550 ( .A(\u_cordic/mycordic/n438 ), .Q(n786) );
  INV3 U1551 ( .A(\u_coder/n218 ), .Q(n1706) );
  XNR21 U1552 ( .A(n771), .B(n773), .Q(n360) );
  XNR21 U1553 ( .A(n761), .B(n763), .Q(n361) );
  XNR21 U1554 ( .A(n769), .B(n772), .Q(n362) );
  XNR21 U1555 ( .A(n759), .B(n762), .Q(n363) );
  XNR21 U1556 ( .A(n772), .B(\u_decoder/I_prefilter [1]), .Q(n364) );
  XNR21 U1557 ( .A(n762), .B(\u_decoder/Q_prefilter [1]), .Q(n365) );
  XNR21 U1558 ( .A(n771), .B(n773), .Q(n366) );
  XNR21 U1559 ( .A(n761), .B(n763), .Q(n367) );
  INV3 U1560 ( .A(\u_inFIFO/n207 ), .Q(n1475) );
  AOI221 U1561 ( .A(\u_inFIFO/n202 ), .B(n34), .C(\u_inFIFO/n203 ), .D(n216), 
        .Q(\u_inFIFO/n207 ) );
  INV3 U1562 ( .A(\u_cdr/phd1/n15 ), .Q(n2252) );
  INV3 U1563 ( .A(\u_cordic/mycordic/n387 ), .Q(n1228) );
  AOI221 U1564 ( .A(n1579), .B(\u_cordic/mycordic/N287 ), .C(n787), .D(
        \u_cordic/mycordic/N255 ), .Q(\u_cordic/mycordic/n387 ) );
  INV3 U1565 ( .A(\u_cordic/mycordic/n536 ), .Q(n1227) );
  NOR21 U1566 ( .A(n787), .B(n1579), .Q(\u_cordic/mycordic/n536 ) );
  INV3 U1567 ( .A(n2649), .Q(n1500) );
  NAND22 U1568 ( .A(n977), .B(n1659), .Q(n2649) );
  INV3 U1569 ( .A(\u_cordic/my_rotation/n83 ), .Q(n1527) );
  NAND22 U1570 ( .A(\u_cordic/my_rotation/next_delta [1]), .B(n974), .Q(
        \u_cordic/my_rotation/n83 ) );
  NAND22 U1571 ( .A(n977), .B(\u_cdr/phd1/n16 ), .Q(\u_cdr/phd1/n18 ) );
  NOR21 U1572 ( .A(n987), .B(n1584), .Q(\u_decoder/iq_demod/n61 ) );
  NAND22 U1573 ( .A(n977), .B(sig_DEMUX_outDEMUX1[0]), .Q(
        \u_decoder/iq_demod/n69 ) );
  INV3 U1574 ( .A(n980), .Q(n978) );
  INV3 U1575 ( .A(n987), .Q(n977) );
  INV3 U1576 ( .A(n983), .Q(n976) );
  INV3 U1577 ( .A(n980), .Q(n974) );
  INV3 U1578 ( .A(n980), .Q(n975) );
  INV3 U1579 ( .A(n981), .Q(n970) );
  INV3 U1580 ( .A(n986), .Q(n971) );
  INV3 U1581 ( .A(n983), .Q(n972) );
  INV3 U1582 ( .A(n984), .Q(n973) );
  INV3 U1583 ( .A(n985), .Q(n969) );
  INV3 U1584 ( .A(n987), .Q(n979) );
  NOR21 U1585 ( .A(n1674), .B(n1696), .Q(sig_DEMUX_outDEMUX18[7]) );
  NOR21 U1586 ( .A(n1676), .B(n1696), .Q(sig_DEMUX_outDEMUX18[6]) );
  NOR21 U1587 ( .A(n1678), .B(n1696), .Q(sig_DEMUX_outDEMUX18[5]) );
  NOR21 U1588 ( .A(n1680), .B(n1696), .Q(sig_DEMUX_outDEMUX18[4]) );
  NOR21 U1589 ( .A(n1666), .B(n1696), .Q(sig_DEMUX_outDEMUX17[7]) );
  NOR21 U1590 ( .A(n1668), .B(n1696), .Q(sig_DEMUX_outDEMUX17[6]) );
  NOR21 U1591 ( .A(n1670), .B(n1696), .Q(sig_DEMUX_outDEMUX17[5]) );
  NOR21 U1592 ( .A(n1672), .B(n1696), .Q(sig_DEMUX_outDEMUX17[4]) );
  XNR21 U1593 ( .A(\u_coder/add_282/carry [19]), .B(\u_coder/j [19]), .Q(n368)
         );
  BUF2 U1594 ( .A(\u_coder/j [0]), .Q(n777) );
  BUF2 U1595 ( .A(\u_coder/i [0]), .Q(n778) );
  XNR21 U1596 ( .A(\u_coder/add_93/carry [19]), .B(\u_coder/c [19]), .Q(n369)
         );
  INV3 U1597 ( .A(\u_coder/n305 ), .Q(n1591) );
  AOI221 U1598 ( .A(n813), .B(\u_coder/i [19]), .C(n810), .D(\u_coder/N726 ), 
        .Q(\u_coder/n305 ) );
  XOR21 U1599 ( .A(\u_coder/add_206/carry [19]), .B(\u_coder/i [19]), .Q(
        \u_coder/N726 ) );
  INV3 U1600 ( .A(\u_coder/n284 ), .Q(n1610) );
  AOI221 U1601 ( .A(n812), .B(\u_coder/i [18]), .C(n811), .D(\u_coder/N725 ), 
        .Q(\u_coder/n284 ) );
  INV3 U1602 ( .A(\u_coder/N1031 ), .Q(n1728) );
  INV3 U1603 ( .A(\u_coder/N1030 ), .Q(n1729) );
  INV3 U1604 ( .A(n387), .Q(\u_cordic/my_rotation/sub_40/carry [1]) );
  NOR21 U1605 ( .A(n61), .B(\u_cordic/my_rotation/present_angle[0][0] ), .Q(
        n387) );
  BUF2 U1606 ( .A(\u_coder/j [3]), .Q(n776) );
  INV3 U1607 ( .A(\u_coder/n287 ), .Q(n1609) );
  AOI221 U1608 ( .A(n813), .B(\u_coder/i [17]), .C(n810), .D(\u_coder/N724 ), 
        .Q(\u_coder/n287 ) );
  INV3 U1609 ( .A(\u_coder/n288 ), .Q(n1608) );
  AOI221 U1610 ( .A(n812), .B(\u_coder/i [16]), .C(n811), .D(\u_coder/N723 ), 
        .Q(\u_coder/n288 ) );
  INV3 U1611 ( .A(\u_coder/N1029 ), .Q(n1730) );
  INV3 U1612 ( .A(\u_cordic/my_rotation/n69 ), .Q(n1513) );
  NAND22 U1613 ( .A(\u_cordic/my_rotation/next_delta [15]), .B(n975), .Q(
        \u_cordic/my_rotation/n69 ) );
  INV3 U1614 ( .A(\u_decoder/fir_filter/n1080 ), .Q(n1828) );
  AOI221 U1615 ( .A(\u_decoder/fir_filter/I_data_mult_4 [10]), .B(n844), .C(
        \u_decoder/fir_filter/I_data_mult_4_buff [10]), .D(n929), .Q(
        \u_decoder/fir_filter/n1080 ) );
  IMUX21 U1616 ( .A(n2502), .B(n2503), .S(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/A2[8] ), .Q(n2501) );
  INV3 U1617 ( .A(\u_decoder/fir_filter/n783 ), .Q(n1899) );
  AOI221 U1618 ( .A(\u_decoder/fir_filter/Q_data_mult_4 [10]), .B(n838), .C(
        \u_decoder/fir_filter/Q_data_mult_4_buff [10]), .D(n932), .Q(
        \u_decoder/fir_filter/n783 ) );
  IMUX21 U1619 ( .A(n2415), .B(n2416), .S(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/A2[8] ), .Q(n2414) );
  INV3 U1620 ( .A(n2540), .Q(n2105) );
  INV3 U1621 ( .A(n2521), .Q(n1985) );
  INV3 U1622 ( .A(n2542), .Q(n2103) );
  INV3 U1623 ( .A(n2523), .Q(n1983) );
  INV3 U1624 ( .A(n2544), .Q(n2101) );
  INV3 U1625 ( .A(n2525), .Q(n1981) );
  INV3 U1626 ( .A(n2538), .Q(n2107) );
  INV3 U1627 ( .A(n2519), .Q(n1987) );
  OAI2111 U1628 ( .A(\u_decoder/fir_filter/I_data_mult_0_buff [1]), .B(
        \u_decoder/fir_filter/I_data_add_1_buff [1]), .C(
        \u_decoder/fir_filter/I_data_mult_0_buff [0]), .D(
        \u_decoder/fir_filter/I_data_add_1_buff [0]), .Q(n2537) );
  OAI2111 U1629 ( .A(\u_decoder/fir_filter/Q_data_mult_0_buff [1]), .B(
        \u_decoder/fir_filter/Q_data_add_1_buff [1]), .C(
        \u_decoder/fir_filter/Q_data_mult_0_buff [0]), .D(
        \u_decoder/fir_filter/Q_data_add_1_buff [0]), .Q(n2518) );
  AOI211 U1630 ( .A(n2549), .B(\u_decoder/fir_filter/I_data_mult_0_buff [7]), 
        .C(n2096), .Q(n2551) );
  INV3 U1631 ( .A(n2548), .Q(n2096) );
  AOI211 U1632 ( .A(n2530), .B(\u_decoder/fir_filter/Q_data_mult_0_buff [7]), 
        .C(n1976), .Q(n2532) );
  INV3 U1633 ( .A(n2529), .Q(n1976) );
  AOI211 U1634 ( .A(n2553), .B(\u_decoder/fir_filter/I_data_mult_0_buff [9]), 
        .C(n2092), .Q(n2555) );
  INV3 U1635 ( .A(n2552), .Q(n2092) );
  AOI211 U1636 ( .A(n2534), .B(\u_decoder/fir_filter/Q_data_mult_0_buff [9]), 
        .C(n1972), .Q(n2536) );
  INV3 U1637 ( .A(n2533), .Q(n1972) );
  INV3 U1638 ( .A(\u_coder/N1028 ), .Q(n1731) );
  INV3 U1639 ( .A(n2551), .Q(n2095) );
  INV3 U1640 ( .A(n2532), .Q(n1975) );
  NOR21 U1641 ( .A(n87), .B(n9), .Q(\u_decoder/fir_filter/add_301/carry [1])
         );
  NOR21 U1642 ( .A(n88), .B(n10), .Q(\u_decoder/fir_filter/add_333/carry [1])
         );
  NOR21 U1643 ( .A(n89), .B(n11), .Q(\u_decoder/fir_filter/add_300/carry [1])
         );
  NOR21 U1644 ( .A(n90), .B(n12), .Q(\u_decoder/fir_filter/add_299/carry [1])
         );
  NOR21 U1645 ( .A(n91), .B(n21), .Q(\u_decoder/fir_filter/add_298/carry [1])
         );
  NOR21 U1646 ( .A(n92), .B(n13), .Q(\u_decoder/fir_filter/add_297/carry [1])
         );
  NOR21 U1647 ( .A(n93), .B(n14), .Q(\u_decoder/fir_filter/add_296/carry [1])
         );
  NOR21 U1648 ( .A(n94), .B(n15), .Q(\u_decoder/fir_filter/add_295/carry [1])
         );
  NOR21 U1649 ( .A(n95), .B(n16), .Q(\u_decoder/fir_filter/add_332/carry [1])
         );
  NOR21 U1650 ( .A(n96), .B(n17), .Q(\u_decoder/fir_filter/add_331/carry [1])
         );
  NOR21 U1651 ( .A(n97), .B(n22), .Q(\u_decoder/fir_filter/add_330/carry [1])
         );
  NOR21 U1652 ( .A(n98), .B(n18), .Q(\u_decoder/fir_filter/add_329/carry [1])
         );
  NOR21 U1653 ( .A(n99), .B(n19), .Q(\u_decoder/fir_filter/add_328/carry [1])
         );
  NOR21 U1654 ( .A(n100), .B(n20), .Q(\u_decoder/fir_filter/add_327/carry [1])
         );
  NAND22 U1655 ( .A(\u_decoder/fir_filter/I_data_mult_3_buff [10]), .B(n923), 
        .Q(\u_decoder/fir_filter/n1096 ) );
  NAND22 U1656 ( .A(\u_decoder/fir_filter/I_data_mult_5_buff [10]), .B(n921), 
        .Q(\u_decoder/fir_filter/n1064 ) );
  NAND22 U1657 ( .A(\u_decoder/fir_filter/Q_data_mult_3_buff [10]), .B(n916), 
        .Q(\u_decoder/fir_filter/n799 ) );
  NAND22 U1658 ( .A(\u_decoder/fir_filter/Q_data_mult_5_buff [10]), .B(n917), 
        .Q(\u_decoder/fir_filter/n767 ) );
  NAND22 U1659 ( .A(\u_decoder/fir_filter/I_data_mult_3_buff [13]), .B(n923), 
        .Q(\u_decoder/fir_filter/n1099 ) );
  NAND22 U1660 ( .A(\u_decoder/fir_filter/I_data_mult_5_buff [13]), .B(n922), 
        .Q(\u_decoder/fir_filter/n1067 ) );
  NAND22 U1661 ( .A(\u_decoder/fir_filter/Q_data_mult_3_buff [13]), .B(n919), 
        .Q(\u_decoder/fir_filter/n802 ) );
  NAND22 U1662 ( .A(\u_decoder/fir_filter/Q_data_mult_5_buff [13]), .B(n917), 
        .Q(\u_decoder/fir_filter/n770 ) );
  NAND22 U1663 ( .A(\u_decoder/fir_filter/I_data_mult_1_buff [12]), .B(n924), 
        .Q(\u_decoder/fir_filter/n1130 ) );
  NAND22 U1664 ( .A(\u_decoder/fir_filter/I_data_mult_7_buff [12]), .B(n919), 
        .Q(\u_decoder/fir_filter/n1032 ) );
  NAND22 U1665 ( .A(\u_decoder/fir_filter/Q_data_mult_1_buff [12]), .B(n915), 
        .Q(\u_decoder/fir_filter/n833 ) );
  NAND22 U1666 ( .A(\u_decoder/fir_filter/Q_data_mult_7_buff [12]), .B(n917), 
        .Q(\u_decoder/fir_filter/n735 ) );
  NAND22 U1667 ( .A(\u_decoder/fir_filter/I_data_mult_0_buff [11]), .B(n924), 
        .Q(\u_decoder/fir_filter/n1145 ) );
  NAND22 U1668 ( .A(\u_decoder/fir_filter/Q_data_mult_0_buff [11]), .B(n915), 
        .Q(\u_decoder/fir_filter/n848 ) );
  NAND22 U1669 ( .A(\u_decoder/fir_filter/I_data_mult_3_buff [12]), .B(n923), 
        .Q(\u_decoder/fir_filter/n1098 ) );
  NAND22 U1670 ( .A(\u_decoder/fir_filter/I_data_mult_5_buff [12]), .B(n922), 
        .Q(\u_decoder/fir_filter/n1066 ) );
  NAND22 U1671 ( .A(\u_decoder/fir_filter/Q_data_mult_3_buff [12]), .B(n918), 
        .Q(\u_decoder/fir_filter/n801 ) );
  NAND22 U1672 ( .A(\u_decoder/fir_filter/Q_data_mult_5_buff [12]), .B(n917), 
        .Q(\u_decoder/fir_filter/n769 ) );
  NAND22 U1673 ( .A(\u_decoder/fir_filter/I_data_mult_2_buff [12]), .B(n923), 
        .Q(\u_decoder/fir_filter/n1114 ) );
  NAND22 U1674 ( .A(\u_decoder/fir_filter/I_data_mult_3_buff [14]), .B(n923), 
        .Q(\u_decoder/fir_filter/n1100 ) );
  NAND22 U1675 ( .A(\u_decoder/fir_filter/I_data_mult_5_buff [14]), .B(n922), 
        .Q(\u_decoder/fir_filter/n1068 ) );
  NAND22 U1676 ( .A(\u_decoder/fir_filter/I_data_mult_6_buff [12]), .B(n920), 
        .Q(\u_decoder/fir_filter/n1049 ) );
  NAND22 U1677 ( .A(\u_decoder/fir_filter/Q_data_mult_2_buff [12]), .B(n932), 
        .Q(\u_decoder/fir_filter/n817 ) );
  NAND22 U1678 ( .A(\u_decoder/fir_filter/Q_data_mult_3_buff [14]), .B(n917), 
        .Q(\u_decoder/fir_filter/n803 ) );
  NAND22 U1679 ( .A(\u_decoder/fir_filter/Q_data_mult_5_buff [14]), .B(n917), 
        .Q(\u_decoder/fir_filter/n771 ) );
  NAND22 U1680 ( .A(\u_decoder/fir_filter/Q_data_mult_6_buff [12]), .B(n918), 
        .Q(\u_decoder/fir_filter/n752 ) );
  NAND22 U1681 ( .A(\u_decoder/fir_filter/n1019 ), .B(
        \u_decoder/fir_filter/n1148 ), .Q(\u_decoder/fir_filter/n1450 ) );
  NAND22 U1682 ( .A(\u_decoder/fir_filter/I_data_mult_0_buff [14]), .B(n913), 
        .Q(\u_decoder/fir_filter/n1148 ) );
  NAND22 U1683 ( .A(\u_decoder/fir_filter/n1019 ), .B(
        \u_decoder/fir_filter/n1147 ), .Q(\u_decoder/fir_filter/n1449 ) );
  NAND22 U1684 ( .A(\u_decoder/fir_filter/I_data_mult_0_buff [13]), .B(n919), 
        .Q(\u_decoder/fir_filter/n1147 ) );
  NAND22 U1685 ( .A(\u_decoder/fir_filter/n1019 ), .B(
        \u_decoder/fir_filter/n1146 ), .Q(\u_decoder/fir_filter/n1448 ) );
  NAND22 U1686 ( .A(\u_decoder/fir_filter/I_data_mult_0_buff [12]), .B(n914), 
        .Q(\u_decoder/fir_filter/n1146 ) );
  NAND22 U1687 ( .A(\u_decoder/fir_filter/n722 ), .B(
        \u_decoder/fir_filter/n851 ), .Q(\u_decoder/fir_filter/n1302 ) );
  NAND22 U1688 ( .A(\u_decoder/fir_filter/Q_data_mult_0_buff [14]), .B(n914), 
        .Q(\u_decoder/fir_filter/n851 ) );
  NAND22 U1689 ( .A(\u_decoder/fir_filter/n722 ), .B(
        \u_decoder/fir_filter/n850 ), .Q(\u_decoder/fir_filter/n1301 ) );
  NAND22 U1690 ( .A(\u_decoder/fir_filter/Q_data_mult_0_buff [13]), .B(n914), 
        .Q(\u_decoder/fir_filter/n850 ) );
  NAND22 U1691 ( .A(\u_decoder/fir_filter/n722 ), .B(
        \u_decoder/fir_filter/n849 ), .Q(\u_decoder/fir_filter/n1300 ) );
  NAND22 U1692 ( .A(\u_decoder/fir_filter/Q_data_mult_0_buff [12]), .B(n914), 
        .Q(\u_decoder/fir_filter/n849 ) );
  NAND22 U1693 ( .A(\u_decoder/fir_filter/n1033 ), .B(
        \u_decoder/fir_filter/n1132 ), .Q(\u_decoder/fir_filter/n1434 ) );
  NAND22 U1694 ( .A(\u_decoder/fir_filter/I_data_mult_1_buff [14]), .B(n924), 
        .Q(\u_decoder/fir_filter/n1132 ) );
  NAND22 U1695 ( .A(\u_decoder/fir_filter/n1033 ), .B(
        \u_decoder/fir_filter/n1131 ), .Q(\u_decoder/fir_filter/n1433 ) );
  NAND22 U1696 ( .A(\u_decoder/fir_filter/I_data_mult_1_buff [13]), .B(n924), 
        .Q(\u_decoder/fir_filter/n1131 ) );
  NAND22 U1697 ( .A(\u_decoder/fir_filter/n1033 ), .B(
        \u_decoder/fir_filter/n1035 ), .Q(\u_decoder/fir_filter/n1354 ) );
  NAND22 U1698 ( .A(\u_decoder/fir_filter/I_data_mult_7_buff [14]), .B(n919), 
        .Q(\u_decoder/fir_filter/n1035 ) );
  NAND22 U1699 ( .A(\u_decoder/fir_filter/n1033 ), .B(
        \u_decoder/fir_filter/n1034 ), .Q(\u_decoder/fir_filter/n1353 ) );
  NAND22 U1700 ( .A(\u_decoder/fir_filter/I_data_mult_7_buff [13]), .B(n919), 
        .Q(\u_decoder/fir_filter/n1034 ) );
  NAND22 U1701 ( .A(\u_decoder/fir_filter/n753 ), .B(
        \u_decoder/fir_filter/n755 ), .Q(\u_decoder/fir_filter/n1222 ) );
  NAND22 U1702 ( .A(\u_decoder/fir_filter/Q_data_mult_6_buff [14]), .B(n918), 
        .Q(\u_decoder/fir_filter/n755 ) );
  NAND22 U1703 ( .A(\u_decoder/fir_filter/n753 ), .B(
        \u_decoder/fir_filter/n754 ), .Q(\u_decoder/fir_filter/n1221 ) );
  NAND22 U1704 ( .A(\u_decoder/fir_filter/Q_data_mult_6_buff [13]), .B(n918), 
        .Q(\u_decoder/fir_filter/n754 ) );
  NAND22 U1705 ( .A(\u_decoder/fir_filter/n736 ), .B(
        \u_decoder/fir_filter/n738 ), .Q(\u_decoder/fir_filter/n1206 ) );
  NAND22 U1706 ( .A(\u_decoder/fir_filter/Q_data_mult_7_buff [14]), .B(n917), 
        .Q(\u_decoder/fir_filter/n738 ) );
  NAND22 U1707 ( .A(\u_decoder/fir_filter/n736 ), .B(
        \u_decoder/fir_filter/n737 ), .Q(\u_decoder/fir_filter/n1205 ) );
  NAND22 U1708 ( .A(\u_decoder/fir_filter/Q_data_mult_7_buff [13]), .B(n917), 
        .Q(\u_decoder/fir_filter/n737 ) );
  NAND22 U1709 ( .A(\u_decoder/fir_filter/n736 ), .B(
        \u_decoder/fir_filter/n835 ), .Q(\u_decoder/fir_filter/n1286 ) );
  NAND22 U1710 ( .A(\u_decoder/fir_filter/Q_data_mult_1_buff [14]), .B(n915), 
        .Q(\u_decoder/fir_filter/n835 ) );
  NAND22 U1711 ( .A(\u_decoder/fir_filter/n736 ), .B(
        \u_decoder/fir_filter/n834 ), .Q(\u_decoder/fir_filter/n1285 ) );
  NAND22 U1712 ( .A(\u_decoder/fir_filter/Q_data_mult_1_buff [13]), .B(n915), 
        .Q(\u_decoder/fir_filter/n834 ) );
  NAND22 U1713 ( .A(\u_decoder/fir_filter/n753 ), .B(
        \u_decoder/fir_filter/n819 ), .Q(\u_decoder/fir_filter/n1270 ) );
  NAND22 U1714 ( .A(\u_decoder/fir_filter/Q_data_mult_2_buff [14]), .B(n915), 
        .Q(\u_decoder/fir_filter/n819 ) );
  NAND22 U1715 ( .A(\u_decoder/fir_filter/n753 ), .B(
        \u_decoder/fir_filter/n818 ), .Q(\u_decoder/fir_filter/n1269 ) );
  NAND22 U1716 ( .A(\u_decoder/fir_filter/Q_data_mult_2_buff [13]), .B(n914), 
        .Q(\u_decoder/fir_filter/n818 ) );
  NAND22 U1717 ( .A(\u_decoder/fir_filter/n1050 ), .B(
        \u_decoder/fir_filter/n1116 ), .Q(\u_decoder/fir_filter/n1418 ) );
  NAND22 U1718 ( .A(\u_decoder/fir_filter/I_data_mult_2_buff [14]), .B(n921), 
        .Q(\u_decoder/fir_filter/n1116 ) );
  NAND22 U1719 ( .A(\u_decoder/fir_filter/n1050 ), .B(
        \u_decoder/fir_filter/n1115 ), .Q(\u_decoder/fir_filter/n1417 ) );
  NAND22 U1720 ( .A(\u_decoder/fir_filter/I_data_mult_2_buff [13]), .B(n923), 
        .Q(\u_decoder/fir_filter/n1115 ) );
  NAND22 U1721 ( .A(\u_decoder/fir_filter/n1050 ), .B(
        \u_decoder/fir_filter/n1052 ), .Q(\u_decoder/fir_filter/n1370 ) );
  NAND22 U1722 ( .A(\u_decoder/fir_filter/I_data_mult_6_buff [14]), .B(n921), 
        .Q(\u_decoder/fir_filter/n1052 ) );
  NAND22 U1723 ( .A(\u_decoder/fir_filter/n1050 ), .B(
        \u_decoder/fir_filter/n1051 ), .Q(\u_decoder/fir_filter/n1369 ) );
  NAND22 U1724 ( .A(\u_decoder/fir_filter/I_data_mult_6_buff [13]), .B(n920), 
        .Q(\u_decoder/fir_filter/n1051 ) );
  INV3 U1725 ( .A(\u_coder/n290 ), .Q(n1606) );
  AOI221 U1726 ( .A(n812), .B(\u_coder/i [14]), .C(n811), .D(\u_coder/N721 ), 
        .Q(\u_coder/n290 ) );
  INV3 U1727 ( .A(\u_coder/n289 ), .Q(n1607) );
  AOI221 U1728 ( .A(n813), .B(\u_coder/i [15]), .C(n810), .D(\u_coder/N722 ), 
        .Q(\u_coder/n289 ) );
  XNR21 U1729 ( .A(n961), .B(n2505), .Q(
        \u_decoder/fir_filter/I_data_mult_4 [14]) );
  XNR21 U1730 ( .A(n963), .B(n2418), .Q(
        \u_decoder/fir_filter/Q_data_mult_4 [14]) );
  INV3 U1731 ( .A(\u_decoder/fir_filter/n982 ), .Q(n2185) );
  AOI221 U1732 ( .A(\u_decoder/fir_filter/I_data_add_7 [14]), .B(n846), .C(
        \u_decoder/fir_filter/I_data_add_7_buff [14]), .D(n931), .Q(
        \u_decoder/fir_filter/n982 ) );
  INV3 U1733 ( .A(\u_decoder/fir_filter/n961 ), .Q(n2170) );
  AOI221 U1734 ( .A(\u_decoder/fir_filter/I_data_add_6 [14]), .B(n847), .C(
        \u_decoder/fir_filter/I_data_add_6_buff [14]), .D(n930), .Q(
        \u_decoder/fir_filter/n961 ) );
  INV3 U1735 ( .A(\u_decoder/fir_filter/n940 ), .Q(n2155) );
  AOI221 U1736 ( .A(\u_decoder/fir_filter/I_data_add_5 [14]), .B(n848), .C(
        \u_decoder/fir_filter/I_data_add_5_buff [14]), .D(n931), .Q(
        \u_decoder/fir_filter/n940 ) );
  INV3 U1737 ( .A(\u_decoder/fir_filter/n919 ), .Q(n2140) );
  AOI221 U1738 ( .A(\u_decoder/fir_filter/I_data_add_4 [14]), .B(n849), .C(
        \u_decoder/fir_filter/I_data_add_4_buff [14]), .D(n932), .Q(
        \u_decoder/fir_filter/n919 ) );
  INV3 U1739 ( .A(\u_decoder/fir_filter/n684 ), .Q(n2065) );
  AOI221 U1740 ( .A(\u_decoder/fir_filter/Q_data_add_7 [14]), .B(n841), .C(
        \u_decoder/fir_filter/Q_data_add_7_buff [14]), .D(n928), .Q(
        \u_decoder/fir_filter/n684 ) );
  INV3 U1741 ( .A(\u_decoder/fir_filter/n663 ), .Q(n2050) );
  AOI221 U1742 ( .A(\u_decoder/fir_filter/Q_data_add_6 [14]), .B(n840), .C(
        \u_decoder/fir_filter/Q_data_add_6_buff [14]), .D(n928), .Q(
        \u_decoder/fir_filter/n663 ) );
  INV3 U1743 ( .A(\u_decoder/fir_filter/n642 ), .Q(n2035) );
  AOI221 U1744 ( .A(\u_decoder/fir_filter/Q_data_add_5 [14]), .B(n840), .C(
        \u_decoder/fir_filter/Q_data_add_5_buff [14]), .D(n927), .Q(
        \u_decoder/fir_filter/n642 ) );
  INV3 U1745 ( .A(\u_decoder/fir_filter/n621 ), .Q(n2020) );
  AOI221 U1746 ( .A(\u_decoder/fir_filter/Q_data_add_4 [14]), .B(n841), .C(
        \u_decoder/fir_filter/Q_data_add_4_buff [14]), .D(n926), .Q(
        \u_decoder/fir_filter/n621 ) );
  INV3 U1747 ( .A(\u_decoder/fir_filter/n600 ), .Q(n2005) );
  AOI221 U1748 ( .A(\u_decoder/fir_filter/Q_data_add_3 [14]), .B(n842), .C(
        \u_decoder/fir_filter/Q_data_add_3_buff [14]), .D(n925), .Q(
        \u_decoder/fir_filter/n600 ) );
  INV3 U1749 ( .A(\u_decoder/fir_filter/n579 ), .Q(n1990) );
  AOI221 U1750 ( .A(\u_decoder/fir_filter/Q_data_add_2 [14]), .B(n843), .C(
        \u_decoder/fir_filter/Q_data_add_2_buff [14]), .D(n926), .Q(
        \u_decoder/fir_filter/n579 ) );
  INV3 U1751 ( .A(\u_decoder/fir_filter/n558 ), .Q(n1966) );
  AOI221 U1752 ( .A(\u_decoder/fir_filter/Q_data_add_1 [14]), .B(n844), .C(
        \u_decoder/fir_filter/Q_data_add_1_buff [14]), .D(n927), .Q(
        \u_decoder/fir_filter/n558 ) );
  INV3 U1753 ( .A(\u_decoder/fir_filter/n555 ), .Q(n1963) );
  AOI221 U1754 ( .A(\u_decoder/fir_filter/Q_data_add_0 [13]), .B(n844), .C(
        sig_decod_outQ[2]), .D(n927), .Q(\u_decoder/fir_filter/n555 ) );
  INV3 U1755 ( .A(\u_decoder/fir_filter/n553 ), .Q(n1962) );
  AOI221 U1756 ( .A(\u_decoder/fir_filter/Q_data_add_0 [14]), .B(n844), .C(
        sig_decod_outQ[3]), .D(n929), .Q(\u_decoder/fir_filter/n553 ) );
  INV3 U1757 ( .A(\u_decoder/fir_filter/n898 ), .Q(n2125) );
  AOI221 U1758 ( .A(\u_decoder/fir_filter/I_data_add_3 [14]), .B(n850), .C(
        \u_decoder/fir_filter/I_data_add_3_buff [14]), .D(n932), .Q(
        \u_decoder/fir_filter/n898 ) );
  INV3 U1759 ( .A(\u_decoder/fir_filter/n877 ), .Q(n2110) );
  AOI221 U1760 ( .A(\u_decoder/fir_filter/I_data_add_2 [14]), .B(n850), .C(
        \u_decoder/fir_filter/I_data_add_2_buff [14]), .D(n920), .Q(
        \u_decoder/fir_filter/n877 ) );
  INV3 U1761 ( .A(\u_decoder/fir_filter/n856 ), .Q(n2086) );
  AOI221 U1762 ( .A(\u_decoder/fir_filter/I_data_add_1 [14]), .B(n851), .C(
        \u_decoder/fir_filter/I_data_add_1_buff [14]), .D(n932), .Q(
        \u_decoder/fir_filter/n856 ) );
  INV3 U1763 ( .A(\u_decoder/fir_filter/n853 ), .Q(n2083) );
  AOI221 U1764 ( .A(\u_decoder/fir_filter/I_data_add_0 [13]), .B(n851), .C(
        sig_decod_outI[2]), .D(n927), .Q(\u_decoder/fir_filter/n853 ) );
  INV3 U1765 ( .A(\u_coder/N1027 ), .Q(n1732) );
  INV3 U1766 ( .A(\u_decoder/fir_filter/n852 ), .Q(n2082) );
  AOI221 U1767 ( .A(\u_decoder/fir_filter/I_data_add_0 [14]), .B(n839), .C(
        sig_decod_outI[3]), .D(n931), .Q(\u_decoder/fir_filter/n852 ) );
  NOR40 U1768 ( .A(n1129), .B(n1128), .C(n1127), .D(n1126), .Q(n1130) );
  NAND41 U1769 ( .A(n2616), .B(n2615), .C(n2614), .D(n2613), .Q(
        \u_cdr/phd1/cnt_phd/N76 ) );
  NAND41 U1770 ( .A(n2603), .B(n2602), .C(n2601), .D(n2600), .Q(
        \u_cdr/dec1/cnt_dec/N76 ) );
  NAND41 U1771 ( .A(n2599), .B(n2598), .C(n2597), .D(n2596), .Q(
        \u_cdr/div1/cnt_div/N76 ) );
  NAND31 U1772 ( .A(\u_cdr/cnt_d [1]), .B(\u_cdr/cnt_d [0]), .C(
        \u_cdr/phd1/cnt_phd/N76 ), .Q(n2629) );
  NAND31 U1773 ( .A(\u_cdr/cnt_d [1]), .B(\u_cdr/cnt_d [0]), .C(
        \u_cdr/dec1/cnt_dec/N76 ), .Q(n2642) );
  NAND31 U1774 ( .A(\u_cdr/cnt_d [1]), .B(\u_cdr/cnt_d [0]), .C(
        \u_cdr/div1/cnt_div/N76 ), .Q(\u_cdr/div1/cnt_div/n48 ) );
  NOR40 U1775 ( .A(n1087), .B(n1039), .C(n1038), .D(n1037), .Q(n2600) );
  NOR40 U1776 ( .A(n1087), .B(n1036), .C(n1035), .D(n1034), .Q(n2596) );
  NOR21 U1777 ( .A(\u_decoder/iq_demod/cos_out [1]), .B(
        \u_decoder/iq_demod/Q_if_buff[3] ), .Q(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/ab[3][1] ) );
  NOR40 U1778 ( .A(n1087), .B(n1076), .C(n1046), .D(n1061), .Q(n2613) );
  INV3 U1779 ( .A(\u_decoder/fir_filter/n1083 ), .Q(n1821) );
  AOI221 U1780 ( .A(\u_decoder/fir_filter/I_data_mult_4 [13]), .B(n848), .C(
        \u_decoder/fir_filter/I_data_mult_4_buff [13]), .D(n932), .Q(
        \u_decoder/fir_filter/n1083 ) );
  INV3 U1781 ( .A(\u_decoder/fir_filter/n786 ), .Q(n1892) );
  AOI221 U1782 ( .A(\u_decoder/fir_filter/Q_data_mult_4 [13]), .B(n837), .C(
        \u_decoder/fir_filter/Q_data_mult_4_buff [13]), .D(n920), .Q(
        \u_decoder/fir_filter/n786 ) );
  BUF6 U1783 ( .A(\u_decoder/I_prefilter [4]), .Q(n766) );
  BUF6 U1784 ( .A(\u_decoder/Q_prefilter [4]), .Q(n756) );
  NOR21 U1785 ( .A(\u_decoder/iq_demod/Q_if_signed [0]), .B(n5), .Q(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/ab[0][3] ) );
  NAND22 U1786 ( .A(\u_decoder/fir_filter/I_data_mult_1_buff [11]), .B(n924), 
        .Q(\u_decoder/fir_filter/n1129 ) );
  NAND22 U1787 ( .A(\u_decoder/fir_filter/I_data_mult_2_buff [11]), .B(n922), 
        .Q(\u_decoder/fir_filter/n1113 ) );
  NAND22 U1788 ( .A(\u_decoder/fir_filter/I_data_mult_6_buff [11]), .B(n920), 
        .Q(\u_decoder/fir_filter/n1048 ) );
  NAND22 U1789 ( .A(\u_decoder/fir_filter/I_data_mult_7_buff [11]), .B(n919), 
        .Q(\u_decoder/fir_filter/n1031 ) );
  NAND22 U1790 ( .A(\u_decoder/fir_filter/Q_data_mult_1_buff [11]), .B(n915), 
        .Q(\u_decoder/fir_filter/n832 ) );
  NAND22 U1791 ( .A(\u_decoder/fir_filter/Q_data_mult_2_buff [11]), .B(n927), 
        .Q(\u_decoder/fir_filter/n816 ) );
  NAND22 U1792 ( .A(\u_decoder/fir_filter/Q_data_mult_6_buff [11]), .B(n918), 
        .Q(\u_decoder/fir_filter/n751 ) );
  NAND22 U1793 ( .A(\u_decoder/fir_filter/Q_data_mult_7_buff [11]), .B(n917), 
        .Q(\u_decoder/fir_filter/n734 ) );
  NAND22 U1794 ( .A(\u_decoder/fir_filter/I_data_mult_0_buff [10]), .B(n924), 
        .Q(\u_decoder/fir_filter/n1144 ) );
  NAND22 U1795 ( .A(\u_decoder/fir_filter/Q_data_mult_0_buff [10]), .B(n914), 
        .Q(\u_decoder/fir_filter/n847 ) );
  NAND22 U1796 ( .A(\u_decoder/fir_filter/I_data_mult_3_buff [11]), .B(n923), 
        .Q(\u_decoder/fir_filter/n1097 ) );
  NAND22 U1797 ( .A(\u_decoder/fir_filter/I_data_mult_5_buff [11]), .B(n921), 
        .Q(\u_decoder/fir_filter/n1065 ) );
  NAND22 U1798 ( .A(\u_decoder/fir_filter/Q_data_mult_3_buff [11]), .B(n916), 
        .Q(\u_decoder/fir_filter/n800 ) );
  NAND22 U1799 ( .A(\u_decoder/fir_filter/Q_data_mult_5_buff [11]), .B(n917), 
        .Q(\u_decoder/fir_filter/n768 ) );
  NOR21 U1800 ( .A(\u_decoder/iq_demod/Q_if_signed [1]), .B(n5), .Q(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/ab[1][3] ) );
  NOR21 U1801 ( .A(n125), .B(n25), .Q(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/ab[2][2] ) );
  NOR21 U1802 ( .A(n708), .B(n709), .Q(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/CARRYB[1][2] ) );
  AOI221 U1803 ( .A(\u_cdr/dec1/cnt_r [0]), .B(n1140), .C(n250), .D(n1139), 
        .Q(\u_cdr/dec1/n33 ) );
  AOI221 U1804 ( .A(\u_cdr/dec1/cnt_r [5]), .B(n1140), .C(\u_cdr/dec1/N65 ), 
        .D(n1139), .Q(\u_cdr/dec1/n32 ) );
  XOR21 U1805 ( .A(\u_cdr/dec1/add_41/carry [5]), .B(\u_cdr/dec1/cnt_r [5]), 
        .Q(\u_cdr/dec1/N65 ) );
  AOI221 U1806 ( .A(\u_cdr/dec1/cnt_r [4]), .B(n1140), .C(\u_cdr/dec1/N64 ), 
        .D(n1139), .Q(\u_cdr/dec1/n26 ) );
  AOI221 U1807 ( .A(\u_cdr/dec1/cnt_r [3]), .B(n1140), .C(\u_cdr/dec1/N63 ), 
        .D(n1139), .Q(\u_cdr/dec1/n29 ) );
  AOI221 U1808 ( .A(\u_cdr/dec1/cnt_r [2]), .B(n1140), .C(\u_cdr/dec1/N62 ), 
        .D(n1139), .Q(\u_cdr/dec1/n30 ) );
  AOI221 U1809 ( .A(\u_cdr/dec1/cnt_r [1]), .B(n1140), .C(\u_cdr/dec1/N61 ), 
        .D(n1139), .Q(\u_cdr/dec1/n31 ) );
  INV3 U1810 ( .A(n2628), .Q(n1143) );
  AOI221 U1811 ( .A(n2622), .B(\u_cdr/phd1/cnt_phd/cnt [0]), .C(n2623), .D(
        n2620), .Q(n2628) );
  INV3 U1812 ( .A(n2627), .Q(n1144) );
  AOI221 U1813 ( .A(n2622), .B(\u_cdr/phd1/cnt_phd/cnt [5]), .C(n2623), .D(
        \u_cdr/phd1/cnt_phd/N84 ), .Q(n2627) );
  XOR21 U1814 ( .A(\u_cdr/phd1/cnt_phd/add_65/carry [5]), .B(
        \u_cdr/phd1/cnt_phd/cnt [5]), .Q(\u_cdr/phd1/cnt_phd/N84 ) );
  INV3 U1815 ( .A(n2621), .Q(n1148) );
  AOI221 U1816 ( .A(n2622), .B(\u_cdr/phd1/cnt_phd/cnt [4]), .C(n2623), .D(
        \u_cdr/phd1/cnt_phd/N83 ), .Q(n2621) );
  INV3 U1817 ( .A(n2624), .Q(n1147) );
  AOI221 U1818 ( .A(n2622), .B(\u_cdr/phd1/cnt_phd/cnt [3]), .C(n2623), .D(
        \u_cdr/phd1/cnt_phd/N82 ), .Q(n2624) );
  INV3 U1819 ( .A(n2625), .Q(n1146) );
  AOI221 U1820 ( .A(n2622), .B(\u_cdr/phd1/cnt_phd/cnt [2]), .C(n2623), .D(
        \u_cdr/phd1/cnt_phd/N81 ), .Q(n2625) );
  INV3 U1821 ( .A(n2626), .Q(n1145) );
  AOI221 U1822 ( .A(n2622), .B(\u_cdr/phd1/cnt_phd/cnt [1]), .C(n2623), .D(
        \u_cdr/phd1/cnt_phd/N80 ), .Q(n2626) );
  INV3 U1823 ( .A(n2641), .Q(n1149) );
  AOI221 U1824 ( .A(n2635), .B(\u_cdr/dec1/cnt_dec/cnt [0]), .C(n2636), .D(
        n196), .Q(n2641) );
  INV3 U1825 ( .A(n2640), .Q(n1150) );
  AOI221 U1826 ( .A(n2635), .B(\u_cdr/dec1/cnt_dec/cnt [5]), .C(n2636), .D(
        \u_cdr/dec1/cnt_dec/N84 ), .Q(n2640) );
  XOR21 U1827 ( .A(\u_cdr/dec1/cnt_dec/add_65/carry [5]), .B(
        \u_cdr/dec1/cnt_dec/cnt [5]), .Q(\u_cdr/dec1/cnt_dec/N84 ) );
  INV3 U1828 ( .A(n2634), .Q(n1154) );
  AOI221 U1829 ( .A(n2635), .B(\u_cdr/dec1/cnt_dec/cnt [4]), .C(n2636), .D(
        \u_cdr/dec1/cnt_dec/N83 ), .Q(n2634) );
  INV3 U1830 ( .A(n2637), .Q(n1153) );
  AOI221 U1831 ( .A(n2635), .B(\u_cdr/dec1/cnt_dec/cnt [3]), .C(n2636), .D(
        \u_cdr/dec1/cnt_dec/N82 ), .Q(n2637) );
  INV3 U1832 ( .A(n2638), .Q(n1152) );
  AOI221 U1833 ( .A(n2635), .B(\u_cdr/dec1/cnt_dec/cnt [2]), .C(n2636), .D(
        \u_cdr/dec1/cnt_dec/N81 ), .Q(n2638) );
  INV3 U1834 ( .A(n2639), .Q(n1151) );
  AOI221 U1835 ( .A(n2635), .B(\u_cdr/dec1/cnt_dec/cnt [1]), .C(n2636), .D(
        \u_cdr/dec1/cnt_dec/N80 ), .Q(n2639) );
  INV3 U1836 ( .A(\u_cdr/div1/cnt_div/n47 ), .Q(n1155) );
  AOI221 U1837 ( .A(\u_cdr/div1/cnt_div/n41 ), .B(\u_cdr/div1/cnt_div/cnt [0]), 
        .C(\u_cdr/div1/cnt_div/n42 ), .D(n197), .Q(\u_cdr/div1/cnt_div/n47 )
         );
  INV3 U1838 ( .A(\u_cdr/div1/cnt_div/n46 ), .Q(n1156) );
  AOI221 U1839 ( .A(\u_cdr/div1/cnt_div/n41 ), .B(\u_cdr/div1/cnt_div/cnt [5]), 
        .C(\u_cdr/div1/cnt_div/n42 ), .D(\u_cdr/div1/cnt_div/N84 ), .Q(
        \u_cdr/div1/cnt_div/n46 ) );
  XOR21 U1840 ( .A(\u_cdr/div1/cnt_div/add_65/carry [5]), .B(
        \u_cdr/div1/cnt_div/cnt [5]), .Q(\u_cdr/div1/cnt_div/N84 ) );
  INV3 U1841 ( .A(\u_cdr/div1/cnt_div/n40 ), .Q(n1160) );
  AOI221 U1842 ( .A(\u_cdr/div1/cnt_div/n41 ), .B(\u_cdr/div1/cnt_div/cnt [4]), 
        .C(\u_cdr/div1/cnt_div/n42 ), .D(\u_cdr/div1/cnt_div/N83 ), .Q(
        \u_cdr/div1/cnt_div/n40 ) );
  INV3 U1843 ( .A(\u_cdr/div1/cnt_div/n43 ), .Q(n1159) );
  AOI221 U1844 ( .A(\u_cdr/div1/cnt_div/n41 ), .B(\u_cdr/div1/cnt_div/cnt [3]), 
        .C(\u_cdr/div1/cnt_div/n42 ), .D(\u_cdr/div1/cnt_div/N82 ), .Q(
        \u_cdr/div1/cnt_div/n43 ) );
  INV3 U1845 ( .A(\u_cdr/div1/cnt_div/n44 ), .Q(n1158) );
  AOI221 U1846 ( .A(\u_cdr/div1/cnt_div/n41 ), .B(\u_cdr/div1/cnt_div/cnt [2]), 
        .C(\u_cdr/div1/cnt_div/n42 ), .D(\u_cdr/div1/cnt_div/N81 ), .Q(
        \u_cdr/div1/cnt_div/n44 ) );
  INV3 U1847 ( .A(\u_cdr/div1/cnt_div/n45 ), .Q(n1157) );
  AOI221 U1848 ( .A(\u_cdr/div1/cnt_div/n41 ), .B(\u_cdr/div1/cnt_div/cnt [1]), 
        .C(\u_cdr/div1/cnt_div/n42 ), .D(\u_cdr/div1/cnt_div/N80 ), .Q(
        \u_cdr/div1/cnt_div/n45 ) );
  INV3 U1849 ( .A(\u_coder/n291 ), .Q(n1605) );
  AOI221 U1850 ( .A(n813), .B(\u_coder/i [13]), .C(n810), .D(\u_coder/N720 ), 
        .Q(\u_coder/n291 ) );
  INV3 U1851 ( .A(\u_decoder/fir_filter/n785 ), .Q(n1890) );
  AOI221 U1852 ( .A(\u_decoder/fir_filter/Q_data_mult_4 [12]), .B(n837), .C(
        \u_decoder/fir_filter/Q_data_mult_4_buff [12]), .D(n924), .Q(
        \u_decoder/fir_filter/n785 ) );
  XOR21 U1853 ( .A(n2428), .B(n2429), .Q(
        \u_decoder/fir_filter/Q_data_mult_4 [12]) );
  NAND22 U1854 ( .A(n1891), .B(n2425), .Q(n2429) );
  INV3 U1855 ( .A(\u_decoder/fir_filter/n784 ), .Q(n1895) );
  AOI221 U1856 ( .A(\u_decoder/fir_filter/Q_data_mult_4 [11]), .B(n837), .C(
        \u_decoder/fir_filter/Q_data_mult_4_buff [11]), .D(n921), .Q(
        \u_decoder/fir_filter/n784 ) );
  XNR21 U1857 ( .A(n2409), .B(n2410), .Q(
        \u_decoder/fir_filter/Q_data_mult_4 [11]) );
  NAND22 U1858 ( .A(n1896), .B(n2411), .Q(n2410) );
  INV3 U1859 ( .A(\u_decoder/fir_filter/n1082 ), .Q(n1819) );
  AOI221 U1860 ( .A(\u_decoder/fir_filter/I_data_mult_4 [12]), .B(n844), .C(
        \u_decoder/fir_filter/I_data_mult_4_buff [12]), .D(n929), .Q(
        \u_decoder/fir_filter/n1082 ) );
  XOR21 U1861 ( .A(n2515), .B(n2516), .Q(
        \u_decoder/fir_filter/I_data_mult_4 [12]) );
  NAND22 U1862 ( .A(n1820), .B(n2512), .Q(n2516) );
  INV3 U1863 ( .A(\u_decoder/fir_filter/n1081 ), .Q(n1824) );
  AOI221 U1864 ( .A(\u_decoder/fir_filter/I_data_mult_4 [11]), .B(n844), .C(
        \u_decoder/fir_filter/I_data_mult_4_buff [11]), .D(n929), .Q(
        \u_decoder/fir_filter/n1081 ) );
  XNR21 U1865 ( .A(n2496), .B(n2497), .Q(
        \u_decoder/fir_filter/I_data_mult_4 [11]) );
  NAND22 U1866 ( .A(n1825), .B(n2498), .Q(n2497) );
  INV3 U1867 ( .A(\u_decoder/fir_filter/n984 ), .Q(n2187) );
  AOI221 U1868 ( .A(\u_decoder/fir_filter/I_data_add_7 [12]), .B(n846), .C(
        \u_decoder/fir_filter/I_data_add_7_buff [12]), .D(n931), .Q(
        \u_decoder/fir_filter/n984 ) );
  INV3 U1869 ( .A(\u_decoder/fir_filter/n983 ), .Q(n2186) );
  AOI221 U1870 ( .A(\u_decoder/fir_filter/I_data_add_7 [13]), .B(n846), .C(
        \u_decoder/fir_filter/I_data_add_7_buff [13]), .D(n931), .Q(
        \u_decoder/fir_filter/n983 ) );
  INV3 U1871 ( .A(\u_decoder/fir_filter/n963 ), .Q(n2172) );
  AOI221 U1872 ( .A(\u_decoder/fir_filter/I_data_add_6 [12]), .B(n847), .C(
        \u_decoder/fir_filter/I_data_add_6_buff [12]), .D(n931), .Q(
        \u_decoder/fir_filter/n963 ) );
  INV3 U1873 ( .A(\u_decoder/fir_filter/n962 ), .Q(n2171) );
  AOI221 U1874 ( .A(\u_decoder/fir_filter/I_data_add_6 [13]), .B(n847), .C(
        \u_decoder/fir_filter/I_data_add_6_buff [13]), .D(n931), .Q(
        \u_decoder/fir_filter/n962 ) );
  INV3 U1875 ( .A(\u_decoder/fir_filter/n942 ), .Q(n2157) );
  AOI221 U1876 ( .A(\u_decoder/fir_filter/I_data_add_5 [12]), .B(n848), .C(
        \u_decoder/fir_filter/I_data_add_5_buff [12]), .D(n928), .Q(
        \u_decoder/fir_filter/n942 ) );
  INV3 U1877 ( .A(\u_decoder/fir_filter/n941 ), .Q(n2156) );
  AOI221 U1878 ( .A(\u_decoder/fir_filter/I_data_add_5 [13]), .B(n848), .C(
        \u_decoder/fir_filter/I_data_add_5_buff [13]), .D(n929), .Q(
        \u_decoder/fir_filter/n941 ) );
  INV3 U1879 ( .A(\u_decoder/fir_filter/n921 ), .Q(n2142) );
  AOI221 U1880 ( .A(\u_decoder/fir_filter/I_data_add_4 [12]), .B(n849), .C(
        \u_decoder/fir_filter/I_data_add_4_buff [12]), .D(n932), .Q(
        \u_decoder/fir_filter/n921 ) );
  INV3 U1881 ( .A(\u_decoder/fir_filter/n920 ), .Q(n2141) );
  AOI221 U1882 ( .A(\u_decoder/fir_filter/I_data_add_4 [13]), .B(n849), .C(
        \u_decoder/fir_filter/I_data_add_4_buff [13]), .D(n932), .Q(
        \u_decoder/fir_filter/n920 ) );
  INV3 U1883 ( .A(\u_decoder/fir_filter/n900 ), .Q(n2127) );
  AOI221 U1884 ( .A(\u_decoder/fir_filter/I_data_add_3 [12]), .B(n849), .C(
        \u_decoder/fir_filter/I_data_add_3_buff [12]), .D(n919), .Q(
        \u_decoder/fir_filter/n900 ) );
  INV3 U1885 ( .A(\u_decoder/fir_filter/n899 ), .Q(n2126) );
  AOI221 U1886 ( .A(\u_decoder/fir_filter/I_data_add_3 [13]), .B(n849), .C(
        \u_decoder/fir_filter/I_data_add_3_buff [13]), .D(n918), .Q(
        \u_decoder/fir_filter/n899 ) );
  INV3 U1887 ( .A(\u_decoder/fir_filter/n686 ), .Q(n2067) );
  AOI221 U1888 ( .A(\u_decoder/fir_filter/Q_data_add_7 [12]), .B(n839), .C(
        \u_decoder/fir_filter/Q_data_add_7_buff [12]), .D(n928), .Q(
        \u_decoder/fir_filter/n686 ) );
  INV3 U1889 ( .A(\u_decoder/fir_filter/n685 ), .Q(n2066) );
  AOI221 U1890 ( .A(\u_decoder/fir_filter/Q_data_add_7 [13]), .B(n839), .C(
        \u_decoder/fir_filter/Q_data_add_7_buff [13]), .D(n928), .Q(
        \u_decoder/fir_filter/n685 ) );
  INV3 U1891 ( .A(\u_decoder/fir_filter/n665 ), .Q(n2052) );
  AOI221 U1892 ( .A(\u_decoder/fir_filter/Q_data_add_6 [12]), .B(n839), .C(
        \u_decoder/fir_filter/Q_data_add_6_buff [12]), .D(n928), .Q(
        \u_decoder/fir_filter/n665 ) );
  INV3 U1893 ( .A(\u_decoder/fir_filter/n664 ), .Q(n2051) );
  AOI221 U1894 ( .A(\u_decoder/fir_filter/Q_data_add_6 [13]), .B(n840), .C(
        \u_decoder/fir_filter/Q_data_add_6_buff [13]), .D(n928), .Q(
        \u_decoder/fir_filter/n664 ) );
  INV3 U1895 ( .A(\u_decoder/fir_filter/n644 ), .Q(n2037) );
  AOI221 U1896 ( .A(\u_decoder/fir_filter/Q_data_add_5 [12]), .B(n840), .C(
        \u_decoder/fir_filter/Q_data_add_5_buff [12]), .D(n927), .Q(
        \u_decoder/fir_filter/n644 ) );
  INV3 U1897 ( .A(\u_decoder/fir_filter/n643 ), .Q(n2036) );
  AOI221 U1898 ( .A(\u_decoder/fir_filter/Q_data_add_5 [13]), .B(n840), .C(
        \u_decoder/fir_filter/Q_data_add_5_buff [13]), .D(n927), .Q(
        \u_decoder/fir_filter/n643 ) );
  INV3 U1899 ( .A(\u_decoder/fir_filter/n623 ), .Q(n2022) );
  AOI221 U1900 ( .A(\u_decoder/fir_filter/Q_data_add_4 [12]), .B(n841), .C(
        \u_decoder/fir_filter/Q_data_add_4_buff [12]), .D(n926), .Q(
        \u_decoder/fir_filter/n623 ) );
  INV3 U1901 ( .A(\u_decoder/fir_filter/n622 ), .Q(n2021) );
  AOI221 U1902 ( .A(\u_decoder/fir_filter/Q_data_add_4 [13]), .B(n841), .C(
        \u_decoder/fir_filter/Q_data_add_4_buff [13]), .D(n926), .Q(
        \u_decoder/fir_filter/n622 ) );
  INV3 U1903 ( .A(\u_decoder/fir_filter/n602 ), .Q(n2007) );
  AOI221 U1904 ( .A(\u_decoder/fir_filter/Q_data_add_3 [12]), .B(n842), .C(
        \u_decoder/fir_filter/Q_data_add_3_buff [12]), .D(n927), .Q(
        \u_decoder/fir_filter/n602 ) );
  INV3 U1905 ( .A(\u_decoder/fir_filter/n601 ), .Q(n2006) );
  AOI221 U1906 ( .A(\u_decoder/fir_filter/Q_data_add_3 [13]), .B(n842), .C(
        \u_decoder/fir_filter/Q_data_add_3_buff [13]), .D(n925), .Q(
        \u_decoder/fir_filter/n601 ) );
  INV3 U1907 ( .A(\u_decoder/fir_filter/n581 ), .Q(n1992) );
  AOI221 U1908 ( .A(\u_decoder/fir_filter/Q_data_add_2 [12]), .B(n843), .C(
        \u_decoder/fir_filter/Q_data_add_2_buff [12]), .D(n925), .Q(
        \u_decoder/fir_filter/n581 ) );
  INV3 U1909 ( .A(\u_decoder/fir_filter/n580 ), .Q(n1991) );
  AOI221 U1910 ( .A(\u_decoder/fir_filter/Q_data_add_2 [13]), .B(n843), .C(
        \u_decoder/fir_filter/Q_data_add_2_buff [13]), .D(n926), .Q(
        \u_decoder/fir_filter/n580 ) );
  INV3 U1911 ( .A(\u_decoder/fir_filter/n560 ), .Q(n1968) );
  AOI221 U1912 ( .A(\u_decoder/fir_filter/Q_data_add_1 [12]), .B(n844), .C(
        \u_decoder/fir_filter/Q_data_add_1_buff [12]), .D(n927), .Q(
        \u_decoder/fir_filter/n560 ) );
  INV3 U1913 ( .A(\u_decoder/fir_filter/n559 ), .Q(n1967) );
  AOI221 U1914 ( .A(\u_decoder/fir_filter/Q_data_add_1 [13]), .B(n844), .C(
        \u_decoder/fir_filter/Q_data_add_1_buff [13]), .D(n927), .Q(
        \u_decoder/fir_filter/n559 ) );
  INV3 U1915 ( .A(\u_decoder/fir_filter/n556 ), .Q(n1964) );
  AOI221 U1916 ( .A(\u_decoder/fir_filter/Q_data_add_0 [12]), .B(n844), .C(
        sig_decod_outQ[1]), .D(n927), .Q(\u_decoder/fir_filter/n556 ) );
  INV3 U1917 ( .A(\u_decoder/fir_filter/n879 ), .Q(n2112) );
  AOI221 U1918 ( .A(\u_decoder/fir_filter/I_data_add_2 [12]), .B(n850), .C(
        \u_decoder/fir_filter/I_data_add_2_buff [12]), .D(n921), .Q(
        \u_decoder/fir_filter/n879 ) );
  INV3 U1919 ( .A(\u_decoder/fir_filter/n878 ), .Q(n2111) );
  AOI221 U1920 ( .A(\u_decoder/fir_filter/I_data_add_2 [13]), .B(n850), .C(
        \u_decoder/fir_filter/I_data_add_2_buff [13]), .D(n923), .Q(
        \u_decoder/fir_filter/n878 ) );
  INV3 U1921 ( .A(\u_decoder/fir_filter/n858 ), .Q(n2088) );
  AOI221 U1922 ( .A(\u_decoder/fir_filter/I_data_add_1 [12]), .B(n851), .C(
        \u_decoder/fir_filter/I_data_add_1_buff [12]), .D(n922), .Q(
        \u_decoder/fir_filter/n858 ) );
  INV3 U1923 ( .A(\u_decoder/fir_filter/n857 ), .Q(n2087) );
  AOI221 U1924 ( .A(\u_decoder/fir_filter/I_data_add_1 [13]), .B(n851), .C(
        \u_decoder/fir_filter/I_data_add_1_buff [13]), .D(n932), .Q(
        \u_decoder/fir_filter/n857 ) );
  INV3 U1925 ( .A(\u_decoder/fir_filter/n854 ), .Q(n2084) );
  AOI221 U1926 ( .A(\u_decoder/fir_filter/I_data_add_0 [12]), .B(n851), .C(
        sig_decod_outI[1]), .D(n919), .Q(\u_decoder/fir_filter/n854 ) );
  INV3 U1927 ( .A(\u_coder/N1026 ), .Q(n1733) );
  NAND41 U1928 ( .A(n2607), .B(n2606), .C(n2605), .D(n2604), .Q(n2612) );
  XNR21 U1929 ( .A(\u_cdr/phd1/cnt_phd/N12 ), .B(\u_cdr/phd1/cnt_phd/cnt [2]), 
        .Q(n2605) );
  XNR21 U1930 ( .A(\u_cdr/phd1/cnt_phd/N13 ), .B(\u_cdr/phd1/cnt_phd/cnt [3]), 
        .Q(n2606) );
  XNR21 U1931 ( .A(n2240), .B(\u_cdr/phd1/cnt_phd/cnt [5]), .Q(n2604) );
  NOR21 U1932 ( .A(\u_decoder/iq_demod/cos_out [1]), .B(
        \u_decoder/iq_demod/I_if_buff[3] ), .Q(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/ab[3][1] ) );
  NOR21 U1933 ( .A(\u_decoder/iq_demod/Q_if_signed [2]), .B(n5), .Q(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/ab[2][3] ) );
  NOR21 U1934 ( .A(\u_decoder/iq_demod/cos_out [2]), .B(
        \u_decoder/iq_demod/Q_if_buff[3] ), .Q(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/ab[3][2] ) );
  NOR21 U1935 ( .A(\u_decoder/iq_demod/I_if_signed [2]), .B(n5), .Q(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/ab[2][3] ) );
  NOR21 U1936 ( .A(\u_decoder/iq_demod/cos_out [2]), .B(
        \u_decoder/iq_demod/I_if_buff[3] ), .Q(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/ab[3][2] ) );
  NOR21 U1937 ( .A(\u_decoder/iq_demod/sin_out [1]), .B(
        \u_decoder/iq_demod/Q_if_buff[3] ), .Q(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/ab[3][1] ) );
  NOR21 U1938 ( .A(\u_decoder/iq_demod/sin_out [1]), .B(
        \u_decoder/iq_demod/I_if_buff[3] ), .Q(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/ab[3][1] ) );
  NOR21 U1939 ( .A(\u_decoder/iq_demod/Q_if_signed [2]), .B(n6), .Q(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/ab[2][3] ) );
  NOR21 U1940 ( .A(\u_decoder/iq_demod/sin_out [2]), .B(
        \u_decoder/iq_demod/Q_if_buff[3] ), .Q(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/ab[3][2] ) );
  NOR21 U1941 ( .A(\u_decoder/iq_demod/I_if_signed [2]), .B(n6), .Q(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/ab[2][3] ) );
  NOR21 U1942 ( .A(\u_decoder/iq_demod/sin_out [2]), .B(
        \u_decoder/iq_demod/I_if_buff[3] ), .Q(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/ab[3][2] ) );
  INV3 U1943 ( .A(\u_coder/N1025 ), .Q(n1734) );
  XNR21 U1944 ( .A(\u_cdr/phd1/cnt_phd/N14 ), .B(\u_cdr/phd1/cnt_phd/cnt [4]), 
        .Q(n2607) );
  NOR21 U1945 ( .A(\u_decoder/iq_demod/Q_if_signed [0]), .B(n6), .Q(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/ab[0][3] ) );
  NOR21 U1946 ( .A(\u_decoder/iq_demod/I_if_signed [0]), .B(n6), .Q(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/ab[0][3] ) );
  NOR21 U1947 ( .A(\u_decoder/iq_demod/I_if_signed [0]), .B(n5), .Q(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/ab[0][3] ) );
  NAND22 U1948 ( .A(\u_decoder/fir_filter/I_data_mult_1_buff [10]), .B(n924), 
        .Q(\u_decoder/fir_filter/n1128 ) );
  NAND22 U1949 ( .A(\u_decoder/fir_filter/I_data_mult_2_buff [10]), .B(n920), 
        .Q(\u_decoder/fir_filter/n1112 ) );
  NAND22 U1950 ( .A(\u_decoder/fir_filter/I_data_mult_2_buff [9]), .B(n921), 
        .Q(\u_decoder/fir_filter/n1111 ) );
  NAND22 U1951 ( .A(\u_decoder/fir_filter/I_data_mult_6_buff [10]), .B(n920), 
        .Q(\u_decoder/fir_filter/n1047 ) );
  NAND22 U1952 ( .A(\u_decoder/fir_filter/I_data_mult_6_buff [9]), .B(n920), 
        .Q(\u_decoder/fir_filter/n1046 ) );
  NAND22 U1953 ( .A(\u_decoder/fir_filter/I_data_mult_7_buff [10]), .B(n919), 
        .Q(\u_decoder/fir_filter/n1030 ) );
  NAND22 U1954 ( .A(\u_decoder/fir_filter/Q_data_mult_1_buff [10]), .B(n915), 
        .Q(\u_decoder/fir_filter/n831 ) );
  NAND22 U1955 ( .A(\u_decoder/fir_filter/Q_data_mult_2_buff [10]), .B(n932), 
        .Q(\u_decoder/fir_filter/n815 ) );
  NAND22 U1956 ( .A(\u_decoder/fir_filter/Q_data_mult_2_buff [9]), .B(n932), 
        .Q(\u_decoder/fir_filter/n814 ) );
  NAND22 U1957 ( .A(\u_decoder/fir_filter/Q_data_mult_6_buff [10]), .B(n917), 
        .Q(\u_decoder/fir_filter/n750 ) );
  NAND22 U1958 ( .A(\u_decoder/fir_filter/Q_data_mult_6_buff [9]), .B(n916), 
        .Q(\u_decoder/fir_filter/n749 ) );
  NAND22 U1959 ( .A(\u_decoder/fir_filter/Q_data_mult_7_buff [10]), .B(n917), 
        .Q(\u_decoder/fir_filter/n733 ) );
  NAND22 U1960 ( .A(\u_decoder/fir_filter/I_data_mult_0_buff [9]), .B(n924), 
        .Q(\u_decoder/fir_filter/n1143 ) );
  NAND22 U1961 ( .A(\u_decoder/fir_filter/Q_data_mult_0_buff [9]), .B(n914), 
        .Q(\u_decoder/fir_filter/n846 ) );
  NAND22 U1962 ( .A(\u_decoder/fir_filter/I_data_mult_0_buff [8]), .B(n919), 
        .Q(\u_decoder/fir_filter/n1142 ) );
  NAND22 U1963 ( .A(\u_decoder/fir_filter/Q_data_mult_0_buff [8]), .B(n915), 
        .Q(\u_decoder/fir_filter/n845 ) );
  NOR21 U1964 ( .A(\u_decoder/iq_demod/Q_if_signed [1]), .B(n6), .Q(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/ab[1][3] ) );
  NOR21 U1965 ( .A(n125), .B(n28), .Q(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/ab[2][2] ) );
  NOR21 U1966 ( .A(n684), .B(n685), .Q(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/CARRYB[1][2] ) );
  NOR21 U1967 ( .A(\u_decoder/iq_demod/I_if_signed [1]), .B(n6), .Q(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/ab[1][3] ) );
  NOR21 U1968 ( .A(n126), .B(n28), .Q(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/ab[2][2] ) );
  NOR21 U1969 ( .A(n720), .B(n721), .Q(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/CARRYB[1][2] ) );
  NOR21 U1970 ( .A(\u_decoder/iq_demod/I_if_signed [1]), .B(n5), .Q(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/ab[1][3] ) );
  NOR21 U1971 ( .A(n126), .B(n25), .Q(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/ab[2][2] ) );
  NOR21 U1972 ( .A(n696), .B(n697), .Q(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/CARRYB[1][2] ) );
  NOR21 U1973 ( .A(\u_decoder/iq_demod/sin_out [0]), .B(
        \u_decoder/iq_demod/Q_if_buff[3] ), .Q(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/ab[3][0] ) );
  NOR21 U1974 ( .A(\u_decoder/iq_demod/sin_out [0]), .B(
        \u_decoder/iq_demod/I_if_buff[3] ), .Q(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/ab[3][0] ) );
  NOR21 U1975 ( .A(\u_decoder/iq_demod/cos_out [0]), .B(
        \u_decoder/iq_demod/Q_if_buff[3] ), .Q(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/ab[3][0] ) );
  NOR21 U1976 ( .A(\u_decoder/iq_demod/cos_out [0]), .B(
        \u_decoder/iq_demod/I_if_buff[3] ), .Q(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/ab[3][0] ) );
  INV3 U1977 ( .A(\u_coder/n293 ), .Q(n1603) );
  AOI221 U1978 ( .A(n813), .B(\u_coder/i [11]), .C(n810), .D(\u_coder/N718 ), 
        .Q(\u_coder/n293 ) );
  INV3 U1979 ( .A(\u_coder/n292 ), .Q(n1604) );
  AOI221 U1980 ( .A(n812), .B(\u_coder/i [12]), .C(n811), .D(\u_coder/N719 ), 
        .Q(\u_coder/n292 ) );
  INV3 U1981 ( .A(\u_decoder/fir_filter/n985 ), .Q(n2188) );
  AOI221 U1982 ( .A(\u_decoder/fir_filter/I_data_add_7 [11]), .B(n846), .C(
        \u_decoder/fir_filter/I_data_add_7_buff [11]), .D(n931), .Q(
        \u_decoder/fir_filter/n985 ) );
  INV3 U1983 ( .A(\u_decoder/fir_filter/n964 ), .Q(n2173) );
  AOI221 U1984 ( .A(\u_decoder/fir_filter/I_data_add_6 [11]), .B(n847), .C(
        \u_decoder/fir_filter/I_data_add_6_buff [11]), .D(n931), .Q(
        \u_decoder/fir_filter/n964 ) );
  INV3 U1985 ( .A(\u_decoder/fir_filter/n943 ), .Q(n2158) );
  AOI221 U1986 ( .A(\u_decoder/fir_filter/I_data_add_5 [11]), .B(n848), .C(
        \u_decoder/fir_filter/I_data_add_5_buff [11]), .D(n930), .Q(
        \u_decoder/fir_filter/n943 ) );
  INV3 U1987 ( .A(\u_decoder/fir_filter/n922 ), .Q(n2143) );
  AOI221 U1988 ( .A(\u_decoder/fir_filter/I_data_add_4 [11]), .B(n848), .C(
        \u_decoder/fir_filter/I_data_add_4_buff [11]), .D(n932), .Q(
        \u_decoder/fir_filter/n922 ) );
  INV3 U1989 ( .A(\u_decoder/fir_filter/n901 ), .Q(n2128) );
  AOI221 U1990 ( .A(\u_decoder/fir_filter/I_data_add_3 [11]), .B(n849), .C(
        \u_decoder/fir_filter/I_data_add_3_buff [11]), .D(n917), .Q(
        \u_decoder/fir_filter/n901 ) );
  INV3 U1991 ( .A(\u_decoder/fir_filter/n687 ), .Q(n2068) );
  AOI221 U1992 ( .A(\u_decoder/fir_filter/Q_data_add_7 [11]), .B(n839), .C(
        \u_decoder/fir_filter/Q_data_add_7_buff [11]), .D(n929), .Q(
        \u_decoder/fir_filter/n687 ) );
  INV3 U1993 ( .A(\u_decoder/fir_filter/n666 ), .Q(n2053) );
  AOI221 U1994 ( .A(\u_decoder/fir_filter/Q_data_add_6 [11]), .B(n839), .C(
        \u_decoder/fir_filter/Q_data_add_6_buff [11]), .D(n928), .Q(
        \u_decoder/fir_filter/n666 ) );
  INV3 U1995 ( .A(\u_decoder/fir_filter/n645 ), .Q(n2038) );
  AOI221 U1996 ( .A(\u_decoder/fir_filter/Q_data_add_5 [11]), .B(n840), .C(
        \u_decoder/fir_filter/Q_data_add_5_buff [11]), .D(n927), .Q(
        \u_decoder/fir_filter/n645 ) );
  INV3 U1997 ( .A(\u_decoder/fir_filter/n624 ), .Q(n2023) );
  AOI221 U1998 ( .A(\u_decoder/fir_filter/Q_data_add_4 [11]), .B(n841), .C(
        \u_decoder/fir_filter/Q_data_add_4_buff [11]), .D(n926), .Q(
        \u_decoder/fir_filter/n624 ) );
  INV3 U1999 ( .A(\u_decoder/fir_filter/n603 ), .Q(n2008) );
  AOI221 U2000 ( .A(\u_decoder/fir_filter/Q_data_add_3 [11]), .B(n842), .C(
        \u_decoder/fir_filter/Q_data_add_3_buff [11]), .D(n925), .Q(
        \u_decoder/fir_filter/n603 ) );
  INV3 U2001 ( .A(\u_decoder/fir_filter/n582 ), .Q(n1993) );
  AOI221 U2002 ( .A(\u_decoder/fir_filter/Q_data_add_2 [11]), .B(n843), .C(
        \u_decoder/fir_filter/Q_data_add_2_buff [11]), .D(n925), .Q(
        \u_decoder/fir_filter/n582 ) );
  INV3 U2003 ( .A(\u_decoder/fir_filter/n561 ), .Q(n1969) );
  AOI221 U2004 ( .A(\u_decoder/fir_filter/Q_data_add_1 [11]), .B(n844), .C(
        \u_decoder/fir_filter/Q_data_add_1_buff [11]), .D(n927), .Q(
        \u_decoder/fir_filter/n561 ) );
  INV3 U2005 ( .A(\u_decoder/fir_filter/n557 ), .Q(n1965) );
  AOI221 U2006 ( .A(\u_decoder/fir_filter/Q_data_add_0 [11]), .B(n844), .C(
        sig_decod_outQ[0]), .D(n927), .Q(\u_decoder/fir_filter/n557 ) );
  INV3 U2007 ( .A(\u_decoder/fir_filter/n880 ), .Q(n2113) );
  AOI221 U2008 ( .A(\u_decoder/fir_filter/I_data_add_2 [11]), .B(n850), .C(
        \u_decoder/fir_filter/I_data_add_2_buff [11]), .D(n926), .Q(
        \u_decoder/fir_filter/n880 ) );
  INV3 U2009 ( .A(\u_decoder/fir_filter/n859 ), .Q(n2089) );
  AOI221 U2010 ( .A(\u_decoder/fir_filter/I_data_add_1 [11]), .B(n851), .C(
        \u_decoder/fir_filter/I_data_add_1_buff [11]), .D(n916), .Q(
        \u_decoder/fir_filter/n859 ) );
  INV3 U2011 ( .A(\u_decoder/fir_filter/n855 ), .Q(n2085) );
  AOI221 U2012 ( .A(\u_decoder/fir_filter/I_data_add_0 [11]), .B(n851), .C(
        sig_decod_outI[0]), .D(n923), .Q(\u_decoder/fir_filter/n855 ) );
  INV3 U2013 ( .A(\u_coder/N1024 ), .Q(n1735) );
  AOI221 U2014 ( .A(\sig_MUX_inMUX5[0] ), .B(n1687), .C(in_MUX_inSEL3), .D(
        sig_DEMUX_outDEMUX2[1]), .Q(n2688) );
  NOR31 U2015 ( .A(n2692), .B(in_DEMUX_inSEL2[2]), .C(in_DEMUX_inSEL2[1]), .Q(
        sig_DEMUX_outDEMUX2[1]) );
  AOI311 U2016 ( .A(n2265), .B(n2266), .C(n2260), .D(
        \u_inFIFO/outWriteCount[5] ), .Q(n2261) );
  OAI2111 U2017 ( .A(\u_inFIFO/outReadCount[3] ), .B(\u_inFIFO/n83 ), .C(n1703), .D(n2259), .Q(n2260) );
  NAND22 U2018 ( .A(\u_inFIFO/outWriteCount[2] ), .B(n106), .Q(n2259) );
  NOR40 U2019 ( .A(n1106), .B(n1105), .C(n1104), .D(n1103), .Q(
        \u_cdr/dec1/N73 ) );
  NAND22 U2020 ( .A(\u_coder/IorQ ), .B(n2688), .Q(\u_coder/n189 ) );
  NOR40 U2021 ( .A(n2232), .B(n2223), .C(n2231), .D(n2230), .Q(
        \u_cordic/my_rotation/n88 ) );
  INV3 U2022 ( .A(\u_cordic/my_rotation/n101 ), .Q(n2232) );
  AOI221 U2023 ( .A(\u_cordic/my_rotation/present_delta [1]), .B(n33), .C(
        \u_cordic/my_rotation/present_delta [1]), .D(n747), .Q(
        \u_cordic/my_rotation/n101 ) );
  NOR31 U2024 ( .A(n1135), .B(n985), .C(n289), .Q(n1094) );
  NOR21 U2025 ( .A(n303), .B(n75), .Q(\u_cordic/mycordic/r173/carry [4]) );
  NOR21 U2026 ( .A(n298), .B(n77), .Q(\u_cordic/mycordic/sub_196/carry[2] ) );
  NOR21 U2027 ( .A(n300), .B(n78), .Q(\u_cordic/mycordic/sub_229/carry[2] ) );
  NOR21 U2028 ( .A(n132), .B(n392), .Q(\u_cordic/mycordic/r173/carry [7]) );
  NOR21 U2029 ( .A(n395), .B(n4), .Q(\u_cordic/mycordic/add_191/carry[3] ) );
  NOR21 U2030 ( .A(n493), .B(n133), .Q(\u_cordic/mycordic/sub_196/carry[5] )
         );
  INV3 U2031 ( .A(\u_cordic/mycordic/sub_196/carry[4] ), .Q(n493) );
  NOR21 U2032 ( .A(n504), .B(n114), .Q(\u_cordic/mycordic/sub_207/carry [4])
         );
  INV3 U2033 ( .A(\u_cordic/mycordic/sub_207/carry [3]), .Q(n504) );
  NOR21 U2034 ( .A(n516), .B(n79), .Q(\u_cordic/mycordic/sub_218/carry[3] ) );
  INV3 U2035 ( .A(\u_cordic/mycordic/sub_218/carry[2] ), .Q(n516) );
  NAND22 U2036 ( .A(\u_inFIFO/outWriteCount[0] ), .B(n105), .Q(n2257) );
  NOR21 U2037 ( .A(n266), .B(n64), .Q(\u_cordic/my_rotation/add_43/carry [5])
         );
  NOR21 U2038 ( .A(n389), .B(n123), .Q(\u_cordic/my_rotation/add_43/carry [8])
         );
  INV3 U2039 ( .A(n395), .Q(\u_cordic/mycordic/add_191/carry[2] ) );
  NOR21 U2040 ( .A(\u_cordic/mycordic/present_ANGLE_table[1][0] ), .B(
        \u_cordic/mycordic/present_ANGLE_table[1][1] ), .Q(n395) );
  INV3 U2041 ( .A(n411), .Q(\u_cordic/mycordic/add_202/carry [3]) );
  NOR21 U2042 ( .A(\u_cordic/mycordic/present_ANGLE_table[2][1] ), .B(
        \u_cordic/mycordic/present_ANGLE_table[2][2] ), .Q(n411) );
  INV3 U2043 ( .A(n426), .Q(\u_cordic/mycordic/add_213/carry[2] ) );
  NOR21 U2044 ( .A(\u_cordic/mycordic/present_ANGLE_table[3][0] ), .B(
        \u_cordic/mycordic/present_ANGLE_table[3][1] ), .Q(n426) );
  INV3 U2045 ( .A(n459), .Q(\u_cordic/mycordic/sub_236/carry [3]) );
  NOR21 U2046 ( .A(\u_cordic/mycordic/present_ANGLE_table[5][1] ), .B(
        \u_cordic/mycordic/present_ANGLE_table[5][2] ), .Q(n459) );
  NOR21 U2047 ( .A(n297), .B(n80), .Q(\u_cordic/mycordic/sub_207/carry [3]) );
  NOR21 U2048 ( .A(n299), .B(n81), .Q(\u_cordic/mycordic/sub_218/carry[2] ) );
  NOR21 U2049 ( .A(n301), .B(n62), .Q(\u_cordic/mycordic/add_233/carry [3]) );
  NOR21 U2050 ( .A(n144), .B(n393), .Q(\u_cordic/mycordic/r173/carry [9]) );
  NOR21 U2051 ( .A(n404), .B(n115), .Q(\u_cordic/mycordic/sub_196/carry[4] )
         );
  NOR21 U2052 ( .A(n397), .B(n116), .Q(\u_cordic/mycordic/add_191/carry[6] )
         );
  NOR21 U2053 ( .A(n484), .B(n134), .Q(\u_cordic/mycordic/add_191/carry[7] )
         );
  INV3 U2054 ( .A(\u_cordic/mycordic/add_191/carry[6] ), .Q(n484) );
  NOR21 U2055 ( .A(n485), .B(n145), .Q(\u_cordic/mycordic/add_191/carry[8] )
         );
  INV3 U2056 ( .A(\u_cordic/mycordic/add_191/carry[7] ), .Q(n485) );
  NOR21 U2057 ( .A(n486), .B(n170), .Q(\u_cordic/mycordic/add_191/carry[9] )
         );
  INV3 U2058 ( .A(\u_cordic/mycordic/add_191/carry[8] ), .Q(n486) );
  NOR21 U2059 ( .A(n487), .B(n171), .Q(\u_cordic/mycordic/add_191/carry[10] )
         );
  INV3 U2060 ( .A(\u_cordic/mycordic/add_191/carry[9] ), .Q(n487) );
  NOR21 U2061 ( .A(n488), .B(n202), .Q(\u_cordic/mycordic/add_191/carry[11] )
         );
  INV3 U2062 ( .A(\u_cordic/mycordic/add_191/carry[10] ), .Q(n488) );
  NOR21 U2063 ( .A(n489), .B(n236), .Q(\u_cordic/mycordic/add_191/carry[12] )
         );
  INV3 U2064 ( .A(\u_cordic/mycordic/add_191/carry[11] ), .Q(n489) );
  NOR21 U2065 ( .A(n490), .B(n261), .Q(\u_cordic/mycordic/add_191/carry[13] )
         );
  INV3 U2066 ( .A(\u_cordic/mycordic/add_191/carry[12] ), .Q(n490) );
  NOR21 U2067 ( .A(n491), .B(n281), .Q(\u_cordic/mycordic/add_191/carry[14] )
         );
  INV3 U2068 ( .A(\u_cordic/mycordic/add_191/carry[13] ), .Q(n491) );
  NOR21 U2069 ( .A(n412), .B(n82), .Q(\u_cordic/mycordic/add_202/carry [5]) );
  NOR21 U2070 ( .A(n494), .B(n117), .Q(\u_cordic/mycordic/add_202/carry [6])
         );
  INV3 U2071 ( .A(\u_cordic/mycordic/add_202/carry [5]), .Q(n494) );
  NOR21 U2072 ( .A(n495), .B(n135), .Q(\u_cordic/mycordic/add_202/carry [7])
         );
  INV3 U2073 ( .A(\u_cordic/mycordic/add_202/carry [6]), .Q(n495) );
  NOR21 U2074 ( .A(n496), .B(n146), .Q(\u_cordic/mycordic/add_202/carry [8])
         );
  INV3 U2075 ( .A(\u_cordic/mycordic/add_202/carry [7]), .Q(n496) );
  NOR21 U2076 ( .A(n497), .B(n172), .Q(\u_cordic/mycordic/add_202/carry [9])
         );
  INV3 U2077 ( .A(\u_cordic/mycordic/add_202/carry [8]), .Q(n497) );
  NOR21 U2078 ( .A(n498), .B(n173), .Q(\u_cordic/mycordic/add_202/carry [10])
         );
  INV3 U2079 ( .A(\u_cordic/mycordic/add_202/carry [9]), .Q(n498) );
  NOR21 U2080 ( .A(n499), .B(n203), .Q(\u_cordic/mycordic/add_202/carry [11])
         );
  INV3 U2081 ( .A(\u_cordic/mycordic/add_202/carry [10]), .Q(n499) );
  NOR21 U2082 ( .A(n500), .B(n237), .Q(\u_cordic/mycordic/add_202/carry [12])
         );
  INV3 U2083 ( .A(\u_cordic/mycordic/add_202/carry [11]), .Q(n500) );
  NOR21 U2084 ( .A(n501), .B(n262), .Q(\u_cordic/mycordic/add_202/carry [13])
         );
  INV3 U2085 ( .A(\u_cordic/mycordic/add_202/carry [12]), .Q(n501) );
  NOR21 U2086 ( .A(n502), .B(n282), .Q(\u_cordic/mycordic/add_202/carry [14])
         );
  INV3 U2087 ( .A(\u_cordic/mycordic/add_202/carry [13]), .Q(n502) );
  NOR21 U2088 ( .A(n427), .B(n83), .Q(\u_cordic/mycordic/add_213/carry[4] ) );
  NOR21 U2089 ( .A(n505), .B(n84), .Q(\u_cordic/mycordic/add_213/carry[5] ) );
  INV3 U2090 ( .A(\u_cordic/mycordic/add_213/carry[4] ), .Q(n505) );
  NOR21 U2091 ( .A(n506), .B(n118), .Q(\u_cordic/mycordic/add_213/carry[6] )
         );
  INV3 U2092 ( .A(\u_cordic/mycordic/add_213/carry[5] ), .Q(n506) );
  NOR21 U2093 ( .A(n507), .B(n136), .Q(\u_cordic/mycordic/add_213/carry[7] )
         );
  INV3 U2094 ( .A(\u_cordic/mycordic/add_213/carry[6] ), .Q(n507) );
  NOR21 U2095 ( .A(n508), .B(n147), .Q(\u_cordic/mycordic/add_213/carry[8] )
         );
  INV3 U2096 ( .A(\u_cordic/mycordic/add_213/carry[7] ), .Q(n508) );
  NOR21 U2097 ( .A(n509), .B(n174), .Q(\u_cordic/mycordic/add_213/carry[9] )
         );
  INV3 U2098 ( .A(\u_cordic/mycordic/add_213/carry[8] ), .Q(n509) );
  NOR21 U2099 ( .A(n510), .B(n175), .Q(\u_cordic/mycordic/add_213/carry[10] )
         );
  INV3 U2100 ( .A(\u_cordic/mycordic/add_213/carry[9] ), .Q(n510) );
  NOR21 U2101 ( .A(n511), .B(n204), .Q(\u_cordic/mycordic/add_213/carry[11] )
         );
  INV3 U2102 ( .A(\u_cordic/mycordic/add_213/carry[10] ), .Q(n511) );
  NOR21 U2103 ( .A(n512), .B(n238), .Q(\u_cordic/mycordic/add_213/carry[12] )
         );
  INV3 U2104 ( .A(\u_cordic/mycordic/add_213/carry[11] ), .Q(n512) );
  NOR21 U2105 ( .A(n513), .B(n263), .Q(\u_cordic/mycordic/add_213/carry[13] )
         );
  INV3 U2106 ( .A(\u_cordic/mycordic/add_213/carry[12] ), .Q(n513) );
  NOR21 U2107 ( .A(n514), .B(n283), .Q(\u_cordic/mycordic/add_213/carry[14] )
         );
  INV3 U2108 ( .A(\u_cordic/mycordic/add_213/carry[13] ), .Q(n514) );
  NOR21 U2109 ( .A(n440), .B(n63), .Q(\u_cordic/mycordic/add_224/carry[3] ) );
  NOR21 U2110 ( .A(n517), .B(n85), .Q(\u_cordic/mycordic/add_224/carry[4] ) );
  INV3 U2111 ( .A(\u_cordic/mycordic/add_224/carry[3] ), .Q(n517) );
  NOR21 U2112 ( .A(n518), .B(n119), .Q(\u_cordic/mycordic/add_224/carry[5] )
         );
  INV3 U2113 ( .A(\u_cordic/mycordic/add_224/carry[4] ), .Q(n518) );
  NOR21 U2114 ( .A(n519), .B(n120), .Q(\u_cordic/mycordic/add_224/carry[6] )
         );
  INV3 U2115 ( .A(\u_cordic/mycordic/add_224/carry[5] ), .Q(n519) );
  NOR21 U2116 ( .A(n520), .B(n137), .Q(\u_cordic/mycordic/add_224/carry[7] )
         );
  INV3 U2117 ( .A(\u_cordic/mycordic/add_224/carry[6] ), .Q(n520) );
  NOR21 U2118 ( .A(n521), .B(n148), .Q(\u_cordic/mycordic/add_224/carry[8] )
         );
  INV3 U2119 ( .A(\u_cordic/mycordic/add_224/carry[7] ), .Q(n521) );
  NOR21 U2120 ( .A(n522), .B(n176), .Q(\u_cordic/mycordic/add_224/carry[9] )
         );
  INV3 U2121 ( .A(\u_cordic/mycordic/add_224/carry[8] ), .Q(n522) );
  NOR21 U2122 ( .A(n523), .B(n205), .Q(\u_cordic/mycordic/add_224/carry[10] )
         );
  INV3 U2123 ( .A(\u_cordic/mycordic/add_224/carry[9] ), .Q(n523) );
  NOR21 U2124 ( .A(n524), .B(n206), .Q(\u_cordic/mycordic/add_224/carry[11] )
         );
  INV3 U2125 ( .A(\u_cordic/mycordic/add_224/carry[10] ), .Q(n524) );
  NOR21 U2126 ( .A(n525), .B(n239), .Q(\u_cordic/mycordic/add_224/carry[12] )
         );
  INV3 U2127 ( .A(\u_cordic/mycordic/add_224/carry[11] ), .Q(n525) );
  NOR21 U2128 ( .A(n526), .B(n264), .Q(\u_cordic/mycordic/add_224/carry[13] )
         );
  INV3 U2129 ( .A(\u_cordic/mycordic/add_224/carry[12] ), .Q(n526) );
  NOR21 U2130 ( .A(n527), .B(n284), .Q(\u_cordic/mycordic/add_224/carry[14] )
         );
  INV3 U2131 ( .A(\u_cordic/mycordic/add_224/carry[13] ), .Q(n527) );
  NOR21 U2132 ( .A(n529), .B(n86), .Q(\u_cordic/mycordic/add_233/carry [4]) );
  INV3 U2133 ( .A(\u_cordic/mycordic/add_233/carry [3]), .Q(n529) );
  NOR21 U2134 ( .A(n530), .B(n121), .Q(\u_cordic/mycordic/add_233/carry [5])
         );
  INV3 U2135 ( .A(\u_cordic/mycordic/add_233/carry [4]), .Q(n530) );
  NOR21 U2136 ( .A(n531), .B(n122), .Q(\u_cordic/mycordic/add_233/carry [6])
         );
  INV3 U2137 ( .A(\u_cordic/mycordic/add_233/carry [5]), .Q(n531) );
  NOR21 U2138 ( .A(n532), .B(n138), .Q(\u_cordic/mycordic/add_233/carry [7])
         );
  INV3 U2139 ( .A(\u_cordic/mycordic/add_233/carry [6]), .Q(n532) );
  NOR21 U2140 ( .A(n533), .B(n149), .Q(\u_cordic/mycordic/add_233/carry [8])
         );
  INV3 U2141 ( .A(\u_cordic/mycordic/add_233/carry [7]), .Q(n533) );
  NOR21 U2142 ( .A(n536), .B(n207), .Q(\u_cordic/mycordic/add_233/carry [11])
         );
  INV3 U2143 ( .A(\u_cordic/mycordic/add_233/carry [10]), .Q(n536) );
  NOR21 U2144 ( .A(n537), .B(n240), .Q(\u_cordic/mycordic/add_233/carry [12])
         );
  INV3 U2145 ( .A(\u_cordic/mycordic/add_233/carry [11]), .Q(n537) );
  NOR21 U2146 ( .A(n169), .B(n478), .Q(\u_cordic/mycordic/r173/carry [10]) );
  INV3 U2147 ( .A(\u_cordic/mycordic/r173/carry [9]), .Q(n478) );
  NOR21 U2148 ( .A(n200), .B(n479), .Q(\u_cordic/mycordic/r173/carry [11]) );
  INV3 U2149 ( .A(\u_cordic/mycordic/r173/carry [10]), .Q(n479) );
  NOR21 U2150 ( .A(n234), .B(n480), .Q(\u_cordic/mycordic/r173/carry [12]) );
  INV3 U2151 ( .A(\u_cordic/mycordic/r173/carry [11]), .Q(n480) );
  NOR21 U2152 ( .A(n235), .B(n481), .Q(\u_cordic/mycordic/r173/carry [13]) );
  INV3 U2153 ( .A(\u_cordic/mycordic/r173/carry [12]), .Q(n481) );
  NOR21 U2154 ( .A(n260), .B(n482), .Q(\u_cordic/mycordic/r173/carry [14]) );
  INV3 U2155 ( .A(\u_cordic/mycordic/r173/carry [13]), .Q(n482) );
  NOR21 U2156 ( .A(\u_coder/stateI[0] ), .B(\u_coder/n189 ), .Q(\u_coder/n155 ) );
  NOR21 U2157 ( .A(n390), .B(n151), .Q(\u_cordic/my_rotation/add_43/carry [10]) );
  NOR21 U2158 ( .A(n473), .B(n152), .Q(\u_cordic/my_rotation/add_43/carry [11]) );
  INV3 U2159 ( .A(\u_cordic/my_rotation/add_43/carry [10]), .Q(n473) );
  NOR21 U2160 ( .A(n474), .B(n179), .Q(\u_cordic/my_rotation/add_43/carry [12]) );
  INV3 U2161 ( .A(\u_cordic/my_rotation/add_43/carry [11]), .Q(n474) );
  NOR21 U2162 ( .A(n475), .B(n213), .Q(\u_cordic/my_rotation/add_43/carry [13]) );
  INV3 U2163 ( .A(\u_cordic/my_rotation/add_43/carry [12]), .Q(n475) );
  NOR21 U2164 ( .A(n476), .B(n241), .Q(\u_cordic/my_rotation/add_43/carry [14]) );
  INV3 U2165 ( .A(\u_cordic/my_rotation/add_43/carry [13]), .Q(n476) );
  NAND22 U2166 ( .A(\u_decoder/fir_filter/I_data_mult_3_buff [9]), .B(n923), 
        .Q(\u_decoder/fir_filter/n1095 ) );
  NAND22 U2167 ( .A(\u_decoder/fir_filter/I_data_mult_5_buff [9]), .B(n921), 
        .Q(\u_decoder/fir_filter/n1063 ) );
  NAND22 U2168 ( .A(\u_decoder/fir_filter/Q_data_mult_3_buff [9]), .B(n919), 
        .Q(\u_decoder/fir_filter/n798 ) );
  NAND22 U2169 ( .A(\u_decoder/fir_filter/Q_data_mult_5_buff [9]), .B(n918), 
        .Q(\u_decoder/fir_filter/n766 ) );
  NAND22 U2170 ( .A(\u_decoder/fir_filter/I_data_mult_1_buff [9]), .B(n924), 
        .Q(\u_decoder/fir_filter/n1127 ) );
  NAND22 U2171 ( .A(\u_decoder/fir_filter/I_data_mult_7_buff [9]), .B(n919), 
        .Q(\u_decoder/fir_filter/n1029 ) );
  NAND22 U2172 ( .A(\u_decoder/fir_filter/Q_data_mult_1_buff [9]), .B(n915), 
        .Q(\u_decoder/fir_filter/n830 ) );
  NAND22 U2173 ( .A(\u_decoder/fir_filter/Q_data_mult_7_buff [9]), .B(n917), 
        .Q(\u_decoder/fir_filter/n732 ) );
  NAND22 U2174 ( .A(\u_decoder/fir_filter/I_data_mult_2_buff [8]), .B(n923), 
        .Q(\u_decoder/fir_filter/n1110 ) );
  NAND22 U2175 ( .A(\u_decoder/fir_filter/I_data_mult_6_buff [8]), .B(n920), 
        .Q(\u_decoder/fir_filter/n1045 ) );
  NAND22 U2176 ( .A(\u_decoder/fir_filter/Q_data_mult_2_buff [8]), .B(n913), 
        .Q(\u_decoder/fir_filter/n813 ) );
  NAND22 U2177 ( .A(\u_decoder/fir_filter/Q_data_mult_6_buff [8]), .B(n918), 
        .Q(\u_decoder/fir_filter/n748 ) );
  NAND22 U2178 ( .A(\u_decoder/fir_filter/I_data_mult_3_buff [8]), .B(n922), 
        .Q(\u_decoder/fir_filter/n1094 ) );
  NAND22 U2179 ( .A(\u_decoder/fir_filter/I_data_mult_5_buff [8]), .B(n921), 
        .Q(\u_decoder/fir_filter/n1062 ) );
  NAND22 U2180 ( .A(\u_decoder/fir_filter/Q_data_mult_3_buff [8]), .B(n918), 
        .Q(\u_decoder/fir_filter/n797 ) );
  NAND22 U2181 ( .A(\u_decoder/fir_filter/Q_data_mult_5_buff [8]), .B(n918), 
        .Q(\u_decoder/fir_filter/n765 ) );
  NAND22 U2182 ( .A(\u_decoder/fir_filter/I_data_mult_1_buff [8]), .B(n924), 
        .Q(\u_decoder/fir_filter/n1126 ) );
  NAND22 U2183 ( .A(\u_decoder/fir_filter/I_data_mult_7_buff [8]), .B(n919), 
        .Q(\u_decoder/fir_filter/n1028 ) );
  NAND22 U2184 ( .A(\u_decoder/fir_filter/Q_data_mult_1_buff [8]), .B(n915), 
        .Q(\u_decoder/fir_filter/n829 ) );
  NAND22 U2185 ( .A(\u_decoder/fir_filter/Q_data_mult_7_buff [8]), .B(n917), 
        .Q(\u_decoder/fir_filter/n731 ) );
  INV3 U2186 ( .A(\u_cordic/mycordic/n399 ), .Q(n1542) );
  NAND22 U2187 ( .A(\u_cordic/mycordic/next_ANGLE_table[6][15] ), .B(n973), 
        .Q(\u_cordic/mycordic/n399 ) );
  INV3 U2188 ( .A(n404), .Q(\u_cordic/mycordic/sub_196/carry[3] ) );
  NOR21 U2189 ( .A(\u_cordic/mycordic/sub_196/carry[2] ), .B(
        \u_cordic/mycordic/present_ANGLE_table[1][2] ), .Q(n404) );
  INV3 U2190 ( .A(n405), .Q(\u_cordic/mycordic/sub_196/carry[6] ) );
  NOR21 U2191 ( .A(\u_cordic/mycordic/sub_196/carry[5] ), .B(
        \u_cordic/mycordic/present_ANGLE_table[1][5] ), .Q(n405) );
  INV3 U2192 ( .A(n419), .Q(\u_cordic/mycordic/sub_207/carry [5]) );
  NOR21 U2193 ( .A(\u_cordic/mycordic/sub_207/carry [4]), .B(
        \u_cordic/mycordic/present_ANGLE_table[2][4] ), .Q(n419) );
  INV3 U2194 ( .A(n422), .Q(\u_cordic/mycordic/sub_207/carry [8]) );
  NOR21 U2195 ( .A(\u_cordic/mycordic/sub_207/carry [7]), .B(
        \u_cordic/mycordic/present_ANGLE_table[2][7] ), .Q(n422) );
  INV3 U2196 ( .A(n434), .Q(\u_cordic/mycordic/sub_218/carry[5] ) );
  NOR21 U2197 ( .A(\u_cordic/mycordic/sub_218/carry[4] ), .B(
        \u_cordic/mycordic/present_ANGLE_table[3][4] ), .Q(n434) );
  INV3 U2198 ( .A(n435), .Q(\u_cordic/mycordic/sub_218/carry[6] ) );
  NOR21 U2199 ( .A(\u_cordic/mycordic/sub_218/carry[5] ), .B(
        \u_cordic/mycordic/present_ANGLE_table[3][5] ), .Q(n435) );
  INV3 U2200 ( .A(n446), .Q(\u_cordic/mycordic/sub_229/carry[3] ) );
  NOR21 U2201 ( .A(\u_cordic/mycordic/sub_229/carry[2] ), .B(
        \u_cordic/mycordic/present_ANGLE_table[4][2] ), .Q(n446) );
  INV3 U2202 ( .A(n448), .Q(\u_cordic/mycordic/sub_229/carry[5] ) );
  NOR21 U2203 ( .A(\u_cordic/mycordic/sub_229/carry[4] ), .B(
        \u_cordic/mycordic/present_ANGLE_table[4][4] ), .Q(n448) );
  INV3 U2204 ( .A(n450), .Q(\u_cordic/mycordic/sub_229/carry[7] ) );
  NOR21 U2205 ( .A(\u_cordic/mycordic/sub_229/carry[6] ), .B(
        \u_cordic/mycordic/present_ANGLE_table[4][6] ), .Q(n450) );
  INV3 U2206 ( .A(n451), .Q(\u_cordic/mycordic/sub_229/carry[8] ) );
  NOR21 U2207 ( .A(\u_cordic/mycordic/sub_229/carry[7] ), .B(
        \u_cordic/mycordic/present_ANGLE_table[4][7] ), .Q(n451) );
  INV3 U2208 ( .A(n460), .Q(\u_cordic/mycordic/sub_236/carry [4]) );
  NOR21 U2209 ( .A(\u_cordic/mycordic/sub_236/carry [3]), .B(
        \u_cordic/mycordic/present_ANGLE_table[5][3] ), .Q(n460) );
  INV3 U2210 ( .A(n462), .Q(\u_cordic/mycordic/sub_236/carry [6]) );
  NOR21 U2211 ( .A(\u_cordic/mycordic/sub_236/carry [5]), .B(
        \u_cordic/mycordic/present_ANGLE_table[5][5] ), .Q(n462) );
  INV3 U2212 ( .A(n464), .Q(\u_cordic/mycordic/sub_236/carry [8]) );
  NOR21 U2213 ( .A(\u_cordic/mycordic/sub_236/carry [7]), .B(
        \u_cordic/mycordic/present_ANGLE_table[5][7] ), .Q(n464) );
  INV3 U2214 ( .A(n391), .Q(\u_cordic/mycordic/r173/carry [5]) );
  NOR21 U2215 ( .A(\u_cordic/mycordic/present_ANGLE_table[6][4] ), .B(
        \u_cordic/mycordic/r173/carry [4]), .Q(n391) );
  INV3 U2216 ( .A(\u_cordic/my_rotation/n99 ), .Q(n2231) );
  AOI221 U2217 ( .A(\u_cordic/my_rotation/present_delta [14]), .B(n33), .C(
        \u_cordic/my_rotation/N55 ), .D(n748), .Q(\u_cordic/my_rotation/n99 )
         );
  XOR21 U2218 ( .A(\u_cordic/my_rotation/present_delta [14]), .B(
        \u_cordic/my_rotation/add_43/carry [14]), .Q(
        \u_cordic/my_rotation/N55 ) );
  INV3 U2219 ( .A(n392), .Q(\u_cordic/mycordic/r173/carry [6]) );
  NOR21 U2220 ( .A(\u_cordic/mycordic/present_ANGLE_table[6][5] ), .B(
        \u_cordic/mycordic/r173/carry [5]), .Q(n392) );
  INV3 U2221 ( .A(n440), .Q(\u_cordic/mycordic/add_224/carry[2] ) );
  NOR21 U2222 ( .A(\u_cordic/mycordic/present_ANGLE_table[4][0] ), .B(
        \u_cordic/mycordic/present_ANGLE_table[4][1] ), .Q(n440) );
  INV3 U2223 ( .A(n393), .Q(\u_cordic/mycordic/r173/carry [8]) );
  NOR21 U2224 ( .A(\u_cordic/mycordic/present_ANGLE_table[6][7] ), .B(
        \u_cordic/mycordic/r173/carry [7]), .Q(n393) );
  INV3 U2225 ( .A(n390), .Q(\u_cordic/my_rotation/add_43/carry [9]) );
  NOR21 U2226 ( .A(\u_cordic/my_rotation/add_43/carry [8]), .B(
        \u_cordic/my_rotation/present_delta [8]), .Q(n390) );
  NOR21 U2227 ( .A(n492), .B(n285), .Q(\u_cordic/mycordic/add_191/carry[15] )
         );
  INV3 U2228 ( .A(\u_cordic/mycordic/add_191/carry[14] ), .Q(n492) );
  NOR21 U2229 ( .A(n503), .B(n286), .Q(\u_cordic/mycordic/add_202/carry [15])
         );
  INV3 U2230 ( .A(\u_cordic/mycordic/add_202/carry [14]), .Q(n503) );
  NOR21 U2231 ( .A(n515), .B(n287), .Q(\u_cordic/mycordic/add_213/carry[15] )
         );
  INV3 U2232 ( .A(\u_cordic/mycordic/add_213/carry[14] ), .Q(n515) );
  NOR21 U2233 ( .A(n528), .B(n306), .Q(\u_cordic/mycordic/add_224/carry[15] )
         );
  INV3 U2234 ( .A(\u_cordic/mycordic/add_224/carry[14] ), .Q(n528) );
  NOR21 U2235 ( .A(n540), .B(n307), .Q(\u_cordic/mycordic/add_233/carry [15])
         );
  INV3 U2236 ( .A(\u_cordic/mycordic/add_233/carry [14]), .Q(n540) );
  INV3 U2237 ( .A(n396), .Q(\u_cordic/mycordic/add_191/carry[4] ) );
  NOR21 U2238 ( .A(\u_cordic/mycordic/add_191/carry[3] ), .B(
        \u_cordic/mycordic/present_ANGLE_table[1][3] ), .Q(n396) );
  INV3 U2239 ( .A(n406), .Q(\u_cordic/mycordic/sub_196/carry[7] ) );
  NOR21 U2240 ( .A(\u_cordic/mycordic/sub_196/carry[6] ), .B(
        \u_cordic/mycordic/present_ANGLE_table[1][6] ), .Q(n406) );
  INV3 U2241 ( .A(n407), .Q(\u_cordic/mycordic/sub_196/carry[8] ) );
  NOR21 U2242 ( .A(\u_cordic/mycordic/sub_196/carry[7] ), .B(
        \u_cordic/mycordic/present_ANGLE_table[1][7] ), .Q(n407) );
  INV3 U2243 ( .A(n408), .Q(\u_cordic/mycordic/sub_196/carry[9] ) );
  NOR21 U2244 ( .A(\u_cordic/mycordic/sub_196/carry[8] ), .B(
        \u_cordic/mycordic/present_ANGLE_table[1][8] ), .Q(n408) );
  INV3 U2245 ( .A(n409), .Q(\u_cordic/mycordic/sub_196/carry[10] ) );
  NOR21 U2246 ( .A(\u_cordic/mycordic/sub_196/carry[9] ), .B(
        \u_cordic/mycordic/present_ANGLE_table[1][9] ), .Q(n409) );
  INV3 U2247 ( .A(n399), .Q(\u_cordic/mycordic/sub_196/carry[11] ) );
  NOR21 U2248 ( .A(\u_cordic/mycordic/sub_196/carry[10] ), .B(
        \u_cordic/mycordic/present_ANGLE_table[1][10] ), .Q(n399) );
  INV3 U2249 ( .A(n400), .Q(\u_cordic/mycordic/sub_196/carry[12] ) );
  NOR21 U2250 ( .A(\u_cordic/mycordic/sub_196/carry[11] ), .B(
        \u_cordic/mycordic/present_ANGLE_table[1][11] ), .Q(n400) );
  INV3 U2251 ( .A(n401), .Q(\u_cordic/mycordic/sub_196/carry[13] ) );
  NOR21 U2252 ( .A(\u_cordic/mycordic/sub_196/carry[12] ), .B(
        \u_cordic/mycordic/present_ANGLE_table[1][12] ), .Q(n401) );
  INV3 U2253 ( .A(n402), .Q(\u_cordic/mycordic/sub_196/carry[14] ) );
  NOR21 U2254 ( .A(\u_cordic/mycordic/sub_196/carry[13] ), .B(
        \u_cordic/mycordic/present_ANGLE_table[1][13] ), .Q(n402) );
  INV3 U2255 ( .A(n420), .Q(\u_cordic/mycordic/sub_207/carry [6]) );
  NOR21 U2256 ( .A(\u_cordic/mycordic/sub_207/carry [5]), .B(
        \u_cordic/mycordic/present_ANGLE_table[2][5] ), .Q(n420) );
  INV3 U2257 ( .A(n421), .Q(\u_cordic/mycordic/sub_207/carry [7]) );
  NOR21 U2258 ( .A(\u_cordic/mycordic/sub_207/carry [6]), .B(
        \u_cordic/mycordic/present_ANGLE_table[2][6] ), .Q(n421) );
  INV3 U2259 ( .A(n423), .Q(\u_cordic/mycordic/sub_207/carry [9]) );
  NOR21 U2260 ( .A(\u_cordic/mycordic/sub_207/carry [8]), .B(
        \u_cordic/mycordic/present_ANGLE_table[2][8] ), .Q(n423) );
  INV3 U2261 ( .A(n424), .Q(\u_cordic/mycordic/sub_207/carry [10]) );
  NOR21 U2262 ( .A(\u_cordic/mycordic/sub_207/carry [9]), .B(
        \u_cordic/mycordic/present_ANGLE_table[2][9] ), .Q(n424) );
  INV3 U2263 ( .A(n414), .Q(\u_cordic/mycordic/sub_207/carry [11]) );
  NOR21 U2264 ( .A(\u_cordic/mycordic/sub_207/carry [10]), .B(
        \u_cordic/mycordic/present_ANGLE_table[2][10] ), .Q(n414) );
  INV3 U2265 ( .A(n415), .Q(\u_cordic/mycordic/sub_207/carry [12]) );
  NOR21 U2266 ( .A(\u_cordic/mycordic/sub_207/carry [11]), .B(
        \u_cordic/mycordic/present_ANGLE_table[2][11] ), .Q(n415) );
  INV3 U2267 ( .A(n416), .Q(\u_cordic/mycordic/sub_207/carry [13]) );
  NOR21 U2268 ( .A(\u_cordic/mycordic/sub_207/carry [12]), .B(
        \u_cordic/mycordic/present_ANGLE_table[2][12] ), .Q(n416) );
  INV3 U2269 ( .A(n417), .Q(\u_cordic/mycordic/sub_207/carry [14]) );
  NOR21 U2270 ( .A(\u_cordic/mycordic/sub_207/carry [13]), .B(
        \u_cordic/mycordic/present_ANGLE_table[2][13] ), .Q(n417) );
  INV3 U2271 ( .A(n433), .Q(\u_cordic/mycordic/sub_218/carry[4] ) );
  NOR21 U2272 ( .A(\u_cordic/mycordic/sub_218/carry[3] ), .B(
        \u_cordic/mycordic/present_ANGLE_table[3][3] ), .Q(n433) );
  INV3 U2273 ( .A(n436), .Q(\u_cordic/mycordic/sub_218/carry[7] ) );
  NOR21 U2274 ( .A(\u_cordic/mycordic/sub_218/carry[6] ), .B(
        \u_cordic/mycordic/present_ANGLE_table[3][6] ), .Q(n436) );
  INV3 U2275 ( .A(n437), .Q(\u_cordic/mycordic/sub_218/carry[8] ) );
  NOR21 U2276 ( .A(\u_cordic/mycordic/sub_218/carry[7] ), .B(
        \u_cordic/mycordic/present_ANGLE_table[3][7] ), .Q(n437) );
  INV3 U2277 ( .A(n438), .Q(\u_cordic/mycordic/sub_218/carry[9] ) );
  NOR21 U2278 ( .A(\u_cordic/mycordic/sub_218/carry[8] ), .B(
        \u_cordic/mycordic/present_ANGLE_table[3][8] ), .Q(n438) );
  INV3 U2279 ( .A(n439), .Q(\u_cordic/mycordic/sub_218/carry[10] ) );
  NOR21 U2280 ( .A(\u_cordic/mycordic/sub_218/carry[9] ), .B(
        \u_cordic/mycordic/present_ANGLE_table[3][9] ), .Q(n439) );
  INV3 U2281 ( .A(n428), .Q(\u_cordic/mycordic/sub_218/carry[11] ) );
  NOR21 U2282 ( .A(\u_cordic/mycordic/sub_218/carry[10] ), .B(
        \u_cordic/mycordic/present_ANGLE_table[3][10] ), .Q(n428) );
  INV3 U2283 ( .A(n429), .Q(\u_cordic/mycordic/sub_218/carry[12] ) );
  NOR21 U2284 ( .A(\u_cordic/mycordic/sub_218/carry[11] ), .B(
        \u_cordic/mycordic/present_ANGLE_table[3][11] ), .Q(n429) );
  INV3 U2285 ( .A(n430), .Q(\u_cordic/mycordic/sub_218/carry[13] ) );
  NOR21 U2286 ( .A(\u_cordic/mycordic/sub_218/carry[12] ), .B(
        \u_cordic/mycordic/present_ANGLE_table[3][12] ), .Q(n430) );
  INV3 U2287 ( .A(n431), .Q(\u_cordic/mycordic/sub_218/carry[14] ) );
  NOR21 U2288 ( .A(\u_cordic/mycordic/sub_218/carry[13] ), .B(
        \u_cordic/mycordic/present_ANGLE_table[3][13] ), .Q(n431) );
  INV3 U2289 ( .A(n447), .Q(\u_cordic/mycordic/sub_229/carry[4] ) );
  NOR21 U2290 ( .A(\u_cordic/mycordic/sub_229/carry[3] ), .B(
        \u_cordic/mycordic/present_ANGLE_table[4][3] ), .Q(n447) );
  INV3 U2291 ( .A(n449), .Q(\u_cordic/mycordic/sub_229/carry[6] ) );
  NOR21 U2292 ( .A(\u_cordic/mycordic/sub_229/carry[5] ), .B(
        \u_cordic/mycordic/present_ANGLE_table[4][5] ), .Q(n449) );
  INV3 U2293 ( .A(n452), .Q(\u_cordic/mycordic/sub_229/carry[9] ) );
  NOR21 U2294 ( .A(\u_cordic/mycordic/sub_229/carry[8] ), .B(
        \u_cordic/mycordic/present_ANGLE_table[4][8] ), .Q(n452) );
  INV3 U2295 ( .A(n453), .Q(\u_cordic/mycordic/sub_229/carry[10] ) );
  NOR21 U2296 ( .A(\u_cordic/mycordic/sub_229/carry[9] ), .B(
        \u_cordic/mycordic/present_ANGLE_table[4][9] ), .Q(n453) );
  INV3 U2297 ( .A(n441), .Q(\u_cordic/mycordic/sub_229/carry[11] ) );
  NOR21 U2298 ( .A(\u_cordic/mycordic/sub_229/carry[10] ), .B(
        \u_cordic/mycordic/present_ANGLE_table[4][10] ), .Q(n441) );
  INV3 U2299 ( .A(n442), .Q(\u_cordic/mycordic/sub_229/carry[12] ) );
  NOR21 U2300 ( .A(\u_cordic/mycordic/sub_229/carry[11] ), .B(
        \u_cordic/mycordic/present_ANGLE_table[4][11] ), .Q(n442) );
  INV3 U2301 ( .A(n443), .Q(\u_cordic/mycordic/sub_229/carry[13] ) );
  NOR21 U2302 ( .A(\u_cordic/mycordic/sub_229/carry[12] ), .B(
        \u_cordic/mycordic/present_ANGLE_table[4][12] ), .Q(n443) );
  INV3 U2303 ( .A(n444), .Q(\u_cordic/mycordic/sub_229/carry[14] ) );
  NOR21 U2304 ( .A(\u_cordic/mycordic/sub_229/carry[13] ), .B(
        \u_cordic/mycordic/present_ANGLE_table[4][13] ), .Q(n444) );
  INV3 U2305 ( .A(n461), .Q(\u_cordic/mycordic/sub_236/carry [5]) );
  NOR21 U2306 ( .A(\u_cordic/mycordic/sub_236/carry [4]), .B(
        \u_cordic/mycordic/present_ANGLE_table[5][4] ), .Q(n461) );
  INV3 U2307 ( .A(n463), .Q(\u_cordic/mycordic/sub_236/carry [7]) );
  NOR21 U2308 ( .A(\u_cordic/mycordic/sub_236/carry [6]), .B(
        \u_cordic/mycordic/present_ANGLE_table[5][6] ), .Q(n463) );
  INV3 U2309 ( .A(n465), .Q(\u_cordic/mycordic/sub_236/carry [9]) );
  NOR21 U2310 ( .A(\u_cordic/mycordic/sub_236/carry [8]), .B(
        \u_cordic/mycordic/present_ANGLE_table[5][8] ), .Q(n465) );
  INV3 U2311 ( .A(n466), .Q(\u_cordic/mycordic/sub_236/carry [10]) );
  NOR21 U2312 ( .A(\u_cordic/mycordic/sub_236/carry [9]), .B(
        \u_cordic/mycordic/present_ANGLE_table[5][9] ), .Q(n466) );
  INV3 U2313 ( .A(n454), .Q(\u_cordic/mycordic/sub_236/carry [11]) );
  NOR21 U2314 ( .A(\u_cordic/mycordic/sub_236/carry [10]), .B(
        \u_cordic/mycordic/present_ANGLE_table[5][10] ), .Q(n454) );
  INV3 U2315 ( .A(n455), .Q(\u_cordic/mycordic/sub_236/carry [12]) );
  NOR21 U2316 ( .A(\u_cordic/mycordic/sub_236/carry [11]), .B(
        \u_cordic/mycordic/present_ANGLE_table[5][11] ), .Q(n455) );
  INV3 U2317 ( .A(n456), .Q(\u_cordic/mycordic/sub_236/carry [13]) );
  NOR21 U2318 ( .A(\u_cordic/mycordic/sub_236/carry [12]), .B(
        \u_cordic/mycordic/present_ANGLE_table[5][12] ), .Q(n456) );
  INV3 U2319 ( .A(n457), .Q(\u_cordic/mycordic/sub_236/carry [14]) );
  NOR21 U2320 ( .A(\u_cordic/mycordic/sub_236/carry [13]), .B(
        \u_cordic/mycordic/present_ANGLE_table[5][13] ), .Q(n457) );
  INV3 U2321 ( .A(n388), .Q(\u_cordic/my_rotation/add_43/carry [6]) );
  NOR21 U2322 ( .A(\u_cordic/my_rotation/add_43/carry [5]), .B(
        \u_cordic/my_rotation/present_delta [5]), .Q(n388) );
  INV3 U2323 ( .A(n397), .Q(\u_cordic/mycordic/add_191/carry[5] ) );
  NOR21 U2324 ( .A(\u_cordic/mycordic/add_191/carry[4] ), .B(
        \u_cordic/mycordic/present_ANGLE_table[1][4] ), .Q(n397) );
  INV3 U2325 ( .A(n412), .Q(\u_cordic/mycordic/add_202/carry [4]) );
  NOR21 U2326 ( .A(\u_cordic/mycordic/add_202/carry [3]), .B(
        \u_cordic/mycordic/present_ANGLE_table[2][3] ), .Q(n412) );
  INV3 U2327 ( .A(n427), .Q(\u_cordic/mycordic/add_213/carry[3] ) );
  NOR21 U2328 ( .A(\u_cordic/mycordic/add_213/carry[2] ), .B(
        \u_cordic/mycordic/present_ANGLE_table[3][2] ), .Q(n427) );
  INV3 U2329 ( .A(n389), .Q(\u_cordic/my_rotation/add_43/carry [7]) );
  NOR21 U2330 ( .A(\u_cordic/my_rotation/add_43/carry [6]), .B(
        \u_cordic/my_rotation/present_delta [6]), .Q(n389) );
  INV3 U2331 ( .A(\u_coder/n303 ), .Q(n1593) );
  AOI221 U2332 ( .A(\u_coder/i [1]), .B(n813), .C(n810), .D(\u_coder/N708 ), 
        .Q(\u_coder/n303 ) );
  INV3 U2333 ( .A(\u_coder/n302 ), .Q(n1594) );
  AOI221 U2334 ( .A(\u_coder/i [2]), .B(n813), .C(n811), .D(\u_coder/N709 ), 
        .Q(\u_coder/n302 ) );
  INV3 U2335 ( .A(n2258), .Q(n1703) );
  AOI2111 U2336 ( .A(n2257), .B(\u_inFIFO/outReadCount[1] ), .C(n1704), .D(
        n2267), .Q(n2258) );
  INV3 U2337 ( .A(n2256), .Q(n1704) );
  INV3 U2338 ( .A(\u_coder/n301 ), .Q(n1595) );
  AOI221 U2339 ( .A(\u_coder/i [3]), .B(n812), .C(n810), .D(\u_coder/N710 ), 
        .Q(\u_coder/n301 ) );
  INV3 U2340 ( .A(n403), .Q(\u_cordic/mycordic/sub_196/carry[15] ) );
  NOR21 U2341 ( .A(\u_cordic/mycordic/sub_196/carry[14] ), .B(
        \u_cordic/mycordic/present_ANGLE_table[1][14] ), .Q(n403) );
  INV3 U2342 ( .A(n418), .Q(\u_cordic/mycordic/sub_207/carry [15]) );
  NOR21 U2343 ( .A(\u_cordic/mycordic/sub_207/carry [14]), .B(
        \u_cordic/mycordic/present_ANGLE_table[2][14] ), .Q(n418) );
  INV3 U2344 ( .A(n432), .Q(\u_cordic/mycordic/sub_218/carry[15] ) );
  NOR21 U2345 ( .A(\u_cordic/mycordic/sub_218/carry[14] ), .B(
        \u_cordic/mycordic/present_ANGLE_table[3][14] ), .Q(n432) );
  INV3 U2346 ( .A(n445), .Q(\u_cordic/mycordic/sub_229/carry[15] ) );
  NOR21 U2347 ( .A(\u_cordic/mycordic/sub_229/carry[14] ), .B(
        \u_cordic/mycordic/present_ANGLE_table[4][14] ), .Q(n445) );
  INV3 U2348 ( .A(n458), .Q(\u_cordic/mycordic/sub_236/carry [15]) );
  NOR21 U2349 ( .A(\u_cordic/mycordic/sub_236/carry [14]), .B(
        \u_cordic/mycordic/present_ANGLE_table[5][14] ), .Q(n458) );
  NOR21 U2350 ( .A(n534), .B(n177), .Q(\u_cordic/mycordic/add_233/carry [9])
         );
  INV3 U2351 ( .A(\u_cordic/mycordic/add_233/carry [8]), .Q(n534) );
  NOR21 U2352 ( .A(n535), .B(n208), .Q(\u_cordic/mycordic/add_233/carry [10])
         );
  INV3 U2353 ( .A(\u_cordic/mycordic/add_233/carry [9]), .Q(n535) );
  NOR21 U2354 ( .A(n538), .B(n265), .Q(\u_cordic/mycordic/add_233/carry [13])
         );
  INV3 U2355 ( .A(\u_cordic/mycordic/add_233/carry [12]), .Q(n538) );
  NOR21 U2356 ( .A(n539), .B(n288), .Q(\u_cordic/mycordic/add_233/carry [14])
         );
  INV3 U2357 ( .A(\u_cordic/mycordic/add_233/carry [13]), .Q(n539) );
  INV3 U2358 ( .A(\u_coder/n294 ), .Q(n1602) );
  AOI221 U2359 ( .A(n812), .B(\u_coder/i [10]), .C(n811), .D(\u_coder/N717 ), 
        .Q(\u_coder/n294 ) );
  INV3 U2360 ( .A(\u_coder/n298 ), .Q(n1598) );
  AOI221 U2361 ( .A(n812), .B(\u_coder/i [6]), .C(n811), .D(\u_coder/N713 ), 
        .Q(\u_coder/n298 ) );
  INV3 U2362 ( .A(\u_coder/n299 ), .Q(n1597) );
  AOI221 U2363 ( .A(n813), .B(\u_coder/i [5]), .C(n810), .D(\u_coder/N712 ), 
        .Q(\u_coder/n299 ) );
  INV3 U2364 ( .A(\u_coder/n295 ), .Q(n1601) );
  AOI221 U2365 ( .A(n813), .B(\u_coder/i [9]), .C(n810), .D(\u_coder/N716 ), 
        .Q(\u_coder/n295 ) );
  INV3 U2366 ( .A(\u_coder/n296 ), .Q(n1600) );
  AOI221 U2367 ( .A(n812), .B(\u_coder/i [8]), .C(n811), .D(\u_coder/N715 ), 
        .Q(\u_coder/n296 ) );
  INV3 U2368 ( .A(\u_coder/n297 ), .Q(n1599) );
  AOI221 U2369 ( .A(n813), .B(\u_coder/i [7]), .C(n810), .D(\u_coder/N714 ), 
        .Q(\u_coder/n297 ) );
  INV3 U2370 ( .A(\u_coder/n300 ), .Q(n1596) );
  AOI221 U2371 ( .A(n812), .B(\u_coder/i [4]), .C(n811), .D(\u_coder/N711 ), 
        .Q(\u_coder/n300 ) );
  NOR21 U2372 ( .A(n279), .B(n483), .Q(\u_cordic/mycordic/r173/carry [15]) );
  INV3 U2373 ( .A(\u_decoder/fir_filter/n1079 ), .Q(n1830) );
  AOI221 U2374 ( .A(\u_decoder/fir_filter/I_data_mult_4 [9]), .B(n845), .C(
        \u_decoder/fir_filter/I_data_mult_4_buff [9]), .D(n929), .Q(
        \u_decoder/fir_filter/n1079 ) );
  INV3 U2375 ( .A(\u_decoder/fir_filter/n782 ), .Q(n1901) );
  AOI221 U2376 ( .A(\u_decoder/fir_filter/Q_data_mult_4 [9]), .B(n837), .C(
        \u_decoder/fir_filter/Q_data_mult_4_buff [9]), .D(n927), .Q(
        \u_decoder/fir_filter/n782 ) );
  INV3 U2377 ( .A(\u_cordic/mycordic/n488 ), .Q(n1303) );
  AOI221 U2378 ( .A(\u_cordic/mycordic/N411 ), .B(n832), .C(
        \u_cordic/mycordic/N443 ), .D(n1582), .Q(\u_cordic/mycordic/n488 ) );
  XOR21 U2379 ( .A(\u_cordic/mycordic/add_202/carry [15]), .B(
        \u_cordic/mycordic/present_ANGLE_table[2][15] ), .Q(
        \u_cordic/mycordic/N411 ) );
  XNR21 U2380 ( .A(\u_cordic/mycordic/sub_207/carry [15]), .B(
        \u_cordic/mycordic/present_ANGLE_table[2][15] ), .Q(
        \u_cordic/mycordic/N443 ) );
  INV3 U2381 ( .A(\u_cordic/mycordic/n505 ), .Q(n1209) );
  AOI221 U2382 ( .A(\u_cordic/mycordic/N346 ), .B(n833), .C(
        \u_cordic/mycordic/N378 ), .D(n1578), .Q(\u_cordic/mycordic/n505 ) );
  XOR21 U2383 ( .A(\u_cordic/mycordic/present_ANGLE_table[1][14] ), .B(
        \u_cordic/mycordic/add_191/carry[14] ), .Q(\u_cordic/mycordic/N346 )
         );
  XNR21 U2384 ( .A(\u_cordic/mycordic/present_ANGLE_table[1][14] ), .B(
        \u_cordic/mycordic/sub_196/carry[14] ), .Q(\u_cordic/mycordic/N378 )
         );
  INV3 U2385 ( .A(\u_cordic/mycordic/n504 ), .Q(n1210) );
  AOI221 U2386 ( .A(\u_cordic/mycordic/N347 ), .B(n834), .C(
        \u_cordic/mycordic/N379 ), .D(n1578), .Q(\u_cordic/mycordic/n504 ) );
  XOR21 U2387 ( .A(\u_cordic/mycordic/add_191/carry[15] ), .B(
        \u_cordic/mycordic/present_ANGLE_table[1][15] ), .Q(
        \u_cordic/mycordic/N347 ) );
  XNR21 U2388 ( .A(\u_cordic/mycordic/sub_196/carry[15] ), .B(
        \u_cordic/mycordic/present_ANGLE_table[1][15] ), .Q(
        \u_cordic/mycordic/N379 ) );
  INV3 U2389 ( .A(\u_decoder/fir_filter/n987 ), .Q(n2190) );
  AOI221 U2390 ( .A(\u_decoder/fir_filter/I_data_add_7 [9]), .B(n846), .C(
        \u_decoder/fir_filter/I_data_add_7_buff [9]), .D(n930), .Q(
        \u_decoder/fir_filter/n987 ) );
  INV3 U2391 ( .A(\u_decoder/fir_filter/n986 ), .Q(n2189) );
  AOI221 U2392 ( .A(\u_decoder/fir_filter/I_data_add_7 [10]), .B(n846), .C(
        \u_decoder/fir_filter/I_data_add_7_buff [10]), .D(n930), .Q(
        \u_decoder/fir_filter/n986 ) );
  INV3 U2393 ( .A(\u_decoder/fir_filter/n966 ), .Q(n2175) );
  AOI221 U2394 ( .A(\u_decoder/fir_filter/I_data_add_6 [9]), .B(n847), .C(
        \u_decoder/fir_filter/I_data_add_6_buff [9]), .D(n931), .Q(
        \u_decoder/fir_filter/n966 ) );
  INV3 U2395 ( .A(\u_decoder/fir_filter/n965 ), .Q(n2174) );
  AOI221 U2396 ( .A(\u_decoder/fir_filter/I_data_add_6 [10]), .B(n847), .C(
        \u_decoder/fir_filter/I_data_add_6_buff [10]), .D(n931), .Q(
        \u_decoder/fir_filter/n965 ) );
  INV3 U2397 ( .A(\u_decoder/fir_filter/n945 ), .Q(n2160) );
  AOI221 U2398 ( .A(\u_decoder/fir_filter/I_data_add_5 [9]), .B(n847), .C(
        \u_decoder/fir_filter/I_data_add_5_buff [9]), .D(n931), .Q(
        \u_decoder/fir_filter/n945 ) );
  INV3 U2399 ( .A(\u_decoder/fir_filter/n944 ), .Q(n2159) );
  AOI221 U2400 ( .A(\u_decoder/fir_filter/I_data_add_5 [10]), .B(n847), .C(
        \u_decoder/fir_filter/I_data_add_5_buff [10]), .D(n928), .Q(
        \u_decoder/fir_filter/n944 ) );
  INV3 U2401 ( .A(\u_decoder/fir_filter/n924 ), .Q(n2145) );
  AOI221 U2402 ( .A(\u_decoder/fir_filter/I_data_add_4 [9]), .B(n848), .C(
        \u_decoder/fir_filter/I_data_add_4_buff [9]), .D(n932), .Q(
        \u_decoder/fir_filter/n924 ) );
  INV3 U2403 ( .A(\u_decoder/fir_filter/n923 ), .Q(n2144) );
  AOI221 U2404 ( .A(\u_decoder/fir_filter/I_data_add_4 [10]), .B(n848), .C(
        \u_decoder/fir_filter/I_data_add_4_buff [10]), .D(n932), .Q(
        \u_decoder/fir_filter/n923 ) );
  INV3 U2405 ( .A(\u_decoder/fir_filter/n903 ), .Q(n2130) );
  AOI221 U2406 ( .A(\u_decoder/fir_filter/I_data_add_3 [9]), .B(n849), .C(
        \u_decoder/fir_filter/I_data_add_3_buff [9]), .D(n918), .Q(
        \u_decoder/fir_filter/n903 ) );
  INV3 U2407 ( .A(\u_decoder/fir_filter/n902 ), .Q(n2129) );
  AOI221 U2408 ( .A(\u_decoder/fir_filter/I_data_add_3 [10]), .B(n849), .C(
        \u_decoder/fir_filter/I_data_add_3_buff [10]), .D(n916), .Q(
        \u_decoder/fir_filter/n902 ) );
  INV3 U2409 ( .A(\u_decoder/fir_filter/n689 ), .Q(n2070) );
  AOI221 U2410 ( .A(\u_decoder/fir_filter/Q_data_add_7 [9]), .B(n839), .C(
        \u_decoder/fir_filter/Q_data_add_7_buff [9]), .D(n929), .Q(
        \u_decoder/fir_filter/n689 ) );
  INV3 U2411 ( .A(\u_decoder/fir_filter/n688 ), .Q(n2069) );
  AOI221 U2412 ( .A(\u_decoder/fir_filter/Q_data_add_7 [10]), .B(n838), .C(
        \u_decoder/fir_filter/Q_data_add_7_buff [10]), .D(n929), .Q(
        \u_decoder/fir_filter/n688 ) );
  INV3 U2413 ( .A(\u_decoder/fir_filter/n668 ), .Q(n2055) );
  AOI221 U2414 ( .A(\u_decoder/fir_filter/Q_data_add_6 [9]), .B(n839), .C(
        \u_decoder/fir_filter/Q_data_add_6_buff [9]), .D(n928), .Q(
        \u_decoder/fir_filter/n668 ) );
  INV3 U2415 ( .A(\u_decoder/fir_filter/n667 ), .Q(n2054) );
  AOI221 U2416 ( .A(\u_decoder/fir_filter/Q_data_add_6 [10]), .B(n839), .C(
        \u_decoder/fir_filter/Q_data_add_6_buff [10]), .D(n928), .Q(
        \u_decoder/fir_filter/n667 ) );
  INV3 U2417 ( .A(\u_decoder/fir_filter/n647 ), .Q(n2040) );
  AOI221 U2418 ( .A(\u_decoder/fir_filter/Q_data_add_5 [9]), .B(n840), .C(
        \u_decoder/fir_filter/Q_data_add_5_buff [9]), .D(n922), .Q(
        \u_decoder/fir_filter/n647 ) );
  INV3 U2419 ( .A(\u_decoder/fir_filter/n646 ), .Q(n2039) );
  AOI221 U2420 ( .A(\u_decoder/fir_filter/Q_data_add_5 [10]), .B(n840), .C(
        \u_decoder/fir_filter/Q_data_add_5_buff [10]), .D(n924), .Q(
        \u_decoder/fir_filter/n646 ) );
  INV3 U2421 ( .A(\u_decoder/fir_filter/n626 ), .Q(n2025) );
  AOI221 U2422 ( .A(\u_decoder/fir_filter/Q_data_add_4 [9]), .B(n841), .C(
        \u_decoder/fir_filter/Q_data_add_4_buff [9]), .D(n926), .Q(
        \u_decoder/fir_filter/n626 ) );
  INV3 U2423 ( .A(\u_decoder/fir_filter/n625 ), .Q(n2024) );
  AOI221 U2424 ( .A(\u_decoder/fir_filter/Q_data_add_4 [10]), .B(n841), .C(
        \u_decoder/fir_filter/Q_data_add_4_buff [10]), .D(n926), .Q(
        \u_decoder/fir_filter/n625 ) );
  INV3 U2425 ( .A(\u_decoder/fir_filter/n605 ), .Q(n2010) );
  AOI221 U2426 ( .A(\u_decoder/fir_filter/Q_data_add_3 [9]), .B(n842), .C(
        \u_decoder/fir_filter/Q_data_add_3_buff [9]), .D(n925), .Q(
        \u_decoder/fir_filter/n605 ) );
  INV3 U2427 ( .A(\u_decoder/fir_filter/n604 ), .Q(n2009) );
  AOI221 U2428 ( .A(\u_decoder/fir_filter/Q_data_add_3 [10]), .B(n842), .C(
        \u_decoder/fir_filter/Q_data_add_3_buff [10]), .D(n925), .Q(
        \u_decoder/fir_filter/n604 ) );
  INV3 U2429 ( .A(\u_decoder/fir_filter/n584 ), .Q(n1995) );
  AOI221 U2430 ( .A(\u_decoder/fir_filter/Q_data_add_2 [9]), .B(n843), .C(
        \u_decoder/fir_filter/Q_data_add_2_buff [9]), .D(n925), .Q(
        \u_decoder/fir_filter/n584 ) );
  INV3 U2431 ( .A(\u_decoder/fir_filter/n583 ), .Q(n1994) );
  AOI221 U2432 ( .A(\u_decoder/fir_filter/Q_data_add_2 [10]), .B(n843), .C(
        \u_decoder/fir_filter/Q_data_add_2_buff [10]), .D(n925), .Q(
        \u_decoder/fir_filter/n583 ) );
  INV3 U2433 ( .A(\u_decoder/fir_filter/n563 ), .Q(n1973) );
  AOI221 U2434 ( .A(\u_decoder/fir_filter/Q_data_add_1 [9]), .B(n844), .C(
        \u_decoder/fir_filter/Q_data_add_1_buff [9]), .D(n928), .Q(
        \u_decoder/fir_filter/n563 ) );
  INV3 U2435 ( .A(\u_decoder/fir_filter/n562 ), .Q(n1970) );
  AOI221 U2436 ( .A(\u_decoder/fir_filter/Q_data_add_1 [10]), .B(n844), .C(
        \u_decoder/fir_filter/Q_data_add_1_buff [10]), .D(n927), .Q(
        \u_decoder/fir_filter/n562 ) );
  INV3 U2437 ( .A(\u_decoder/fir_filter/n882 ), .Q(n2115) );
  AOI221 U2438 ( .A(\u_decoder/fir_filter/I_data_add_2 [9]), .B(n850), .C(
        \u_decoder/fir_filter/I_data_add_2_buff [9]), .D(n925), .Q(
        \u_decoder/fir_filter/n882 ) );
  INV3 U2439 ( .A(\u_decoder/fir_filter/n881 ), .Q(n2114) );
  AOI221 U2440 ( .A(\u_decoder/fir_filter/I_data_add_2 [10]), .B(n850), .C(
        \u_decoder/fir_filter/I_data_add_2_buff [10]), .D(n920), .Q(
        \u_decoder/fir_filter/n881 ) );
  INV3 U2441 ( .A(\u_decoder/fir_filter/n861 ), .Q(n2093) );
  AOI221 U2442 ( .A(\u_decoder/fir_filter/I_data_add_1 [9]), .B(n851), .C(
        \u_decoder/fir_filter/I_data_add_1_buff [9]), .D(n921), .Q(
        \u_decoder/fir_filter/n861 ) );
  INV3 U2443 ( .A(\u_decoder/fir_filter/n860 ), .Q(n2090) );
  AOI221 U2444 ( .A(\u_decoder/fir_filter/I_data_add_1 [10]), .B(n851), .C(
        \u_decoder/fir_filter/I_data_add_1_buff [10]), .D(n915), .Q(
        \u_decoder/fir_filter/n860 ) );
  INV3 U2445 ( .A(\u_cordic/mycordic/n473 ), .Q(n1277) );
  AOI221 U2446 ( .A(\u_cordic/mycordic/N470 ), .B(n836), .C(
        \u_cordic/mycordic/N498 ), .D(n1581), .Q(\u_cordic/mycordic/n473 ) );
  XOR21 U2447 ( .A(\u_cordic/mycordic/present_ANGLE_table[3][14] ), .B(
        \u_cordic/mycordic/add_213/carry[14] ), .Q(\u_cordic/mycordic/N470 )
         );
  XNR21 U2448 ( .A(\u_cordic/mycordic/present_ANGLE_table[3][14] ), .B(
        \u_cordic/mycordic/sub_218/carry[14] ), .Q(\u_cordic/mycordic/N498 )
         );
  INV3 U2449 ( .A(\u_cordic/mycordic/n472 ), .Q(n1278) );
  AOI221 U2450 ( .A(\u_cordic/mycordic/N471 ), .B(n836), .C(
        \u_cordic/mycordic/N499 ), .D(n1581), .Q(\u_cordic/mycordic/n472 ) );
  XOR21 U2451 ( .A(\u_cordic/mycordic/add_213/carry[15] ), .B(
        \u_cordic/mycordic/present_ANGLE_table[3][15] ), .Q(
        \u_cordic/mycordic/N471 ) );
  XNR21 U2452 ( .A(\u_cordic/mycordic/sub_218/carry[15] ), .B(
        \u_cordic/mycordic/present_ANGLE_table[3][15] ), .Q(
        \u_cordic/mycordic/N499 ) );
  INV3 U2453 ( .A(\u_cordic/mycordic/n458 ), .Q(n1252) );
  AOI221 U2454 ( .A(\u_cordic/mycordic/N514 ), .B(n789), .C(
        \u_cordic/mycordic/N531 ), .D(n1580), .Q(\u_cordic/mycordic/n458 ) );
  XOR21 U2455 ( .A(\u_cordic/mycordic/present_ANGLE_table[4][13] ), .B(
        \u_cordic/mycordic/add_224/carry[13] ), .Q(\u_cordic/mycordic/N514 )
         );
  XNR21 U2456 ( .A(\u_cordic/mycordic/present_ANGLE_table[4][13] ), .B(
        \u_cordic/mycordic/sub_229/carry[13] ), .Q(\u_cordic/mycordic/N531 )
         );
  INV3 U2457 ( .A(\u_cordic/mycordic/n457 ), .Q(n1253) );
  AOI221 U2458 ( .A(\u_cordic/mycordic/N515 ), .B(n789), .C(
        \u_cordic/mycordic/N532 ), .D(n1580), .Q(\u_cordic/mycordic/n457 ) );
  XOR21 U2459 ( .A(\u_cordic/mycordic/present_ANGLE_table[4][14] ), .B(
        \u_cordic/mycordic/add_224/carry[14] ), .Q(\u_cordic/mycordic/N515 )
         );
  XNR21 U2460 ( .A(\u_cordic/mycordic/present_ANGLE_table[4][14] ), .B(
        \u_cordic/mycordic/sub_229/carry[14] ), .Q(\u_cordic/mycordic/N532 )
         );
  INV3 U2461 ( .A(\u_cordic/mycordic/n439 ), .Q(n1193) );
  AOI221 U2462 ( .A(\u_cordic/mycordic/N548 ), .B(n786), .C(
        \u_cordic/mycordic/N564 ), .D(n1577), .Q(\u_cordic/mycordic/n439 ) );
  XOR21 U2463 ( .A(\u_cordic/mycordic/present_ANGLE_table[5][14] ), .B(
        \u_cordic/mycordic/add_233/carry [14]), .Q(\u_cordic/mycordic/N548 )
         );
  XNR21 U2464 ( .A(\u_cordic/mycordic/present_ANGLE_table[5][14] ), .B(
        \u_cordic/mycordic/sub_236/carry [14]), .Q(\u_cordic/mycordic/N564 )
         );
  INV3 U2465 ( .A(\u_cordic/mycordic/n455 ), .Q(n1254) );
  AOI221 U2466 ( .A(\u_cordic/mycordic/N516 ), .B(n789), .C(
        \u_cordic/mycordic/N533 ), .D(n1580), .Q(\u_cordic/mycordic/n455 ) );
  XOR21 U2467 ( .A(\u_cordic/mycordic/add_224/carry[15] ), .B(
        \u_cordic/mycordic/present_ANGLE_table[4][15] ), .Q(
        \u_cordic/mycordic/N516 ) );
  XNR21 U2468 ( .A(\u_cordic/mycordic/sub_229/carry[15] ), .B(
        \u_cordic/mycordic/present_ANGLE_table[4][15] ), .Q(
        \u_cordic/mycordic/N533 ) );
  INV3 U2469 ( .A(\u_cordic/mycordic/n437 ), .Q(n1194) );
  AOI221 U2470 ( .A(\u_cordic/mycordic/N549 ), .B(n786), .C(
        \u_cordic/mycordic/N565 ), .D(n1577), .Q(\u_cordic/mycordic/n437 ) );
  XOR21 U2471 ( .A(\u_cordic/mycordic/add_233/carry [15]), .B(
        \u_cordic/mycordic/present_ANGLE_table[5][15] ), .Q(
        \u_cordic/mycordic/N549 ) );
  XNR21 U2472 ( .A(\u_cordic/mycordic/sub_236/carry [15]), .B(
        \u_cordic/mycordic/present_ANGLE_table[5][15] ), .Q(
        \u_cordic/mycordic/N565 ) );
  INV3 U2473 ( .A(\u_coder/N1023 ), .Q(n1736) );
  INV3 U2474 ( .A(n2643), .Q(n1494) );
  NAND22 U2475 ( .A(\u_cdr/dec1/cnt_dec/N43 ), .B(n976), .Q(n2643) );
  NOR40 U2476 ( .A(n1088), .B(\u_cdr/dec1/cnt_dec/cnt [5]), .C(n1087), .D(
        n1086), .Q(\u_cdr/dec1/cnt_dec/N43 ) );
  NOR21 U2477 ( .A(\u_cordic/mycordic/present_I_table[4][1] ), .B(n2216), .Q(
        n2579) );
  INV3 U2478 ( .A(n2580), .Q(n2216) );
  INV3 U2479 ( .A(n2569), .Q(n2211) );
  NAND22 U2480 ( .A(n156), .B(n2570), .Q(n2569) );
  AOI221 U2481 ( .A(n2568), .B(\u_cordic/mycordic/present_Q_table[5][1] ), .C(
        n32), .D(n2213), .Q(n2570) );
  NOR21 U2482 ( .A(\u_coder/stateQ[0] ), .B(\u_coder/n234 ), .Q(\u_coder/n205 ) );
  AOI211 U2483 ( .A(\u_cordic/mycordic/present_I_table[4][1] ), .B(
        \u_cordic/mycordic/present_Q_table[4][4] ), .C(n2220), .Q(n2587) );
  INV3 U2484 ( .A(n2585), .Q(n2220) );
  OAI2111 U2485 ( .A(\u_cordic/mycordic/present_I_table[4][1] ), .B(
        \u_cordic/mycordic/present_Q_table[4][4] ), .C(
        \u_cordic/mycordic/present_I_table[4][0] ), .D(
        \u_cordic/mycordic/present_Q_table[4][3] ), .Q(n2585) );
  NAND22 U2486 ( .A(n2688), .B(\u_coder/n139 ), .Q(\u_coder/n234 ) );
  INV3 U2487 ( .A(n2587), .Q(n2219) );
  INV3 U2488 ( .A(n2562), .Q(n2208) );
  AOI211 U2489 ( .A(n2560), .B(\u_cordic/mycordic/present_Q_table[5][3] ), .C(
        n2209), .Q(n2562) );
  INV3 U2490 ( .A(n2557), .Q(n2212) );
  XNR21 U2491 ( .A(\u_outFIFO/r98/carry [5]), .B(\u_outFIFO/outWriteCount[5] ), 
        .Q(\u_outFIFO/N136 ) );
  XNR21 U2492 ( .A(\u_inFIFO/r96/carry [5]), .B(\u_inFIFO/outWriteCount[5] ), 
        .Q(\u_inFIFO/N128 ) );
  OAI2111 U2493 ( .A(\u_cordic/mycordic/present_Q_table[5][1] ), .B(
        \u_cordic/mycordic/present_I_table[5][5] ), .C(
        \u_cordic/mycordic/present_Q_table[5][0] ), .D(
        \u_cordic/mycordic/present_I_table[5][4] ), .Q(n2556) );
  NOR40 U2494 ( .A(n2236), .B(n2235), .C(n2234), .D(n2233), .Q(
        \u_cordic/my_rotation/n87 ) );
  INV3 U2495 ( .A(\u_cordic/my_rotation/n102 ), .Q(n2233) );
  AOI221 U2496 ( .A(\u_cordic/my_rotation/N41 ), .B(n33), .C(
        \u_cordic/my_rotation/N41 ), .D(n747), .Q(\u_cordic/my_rotation/n102 )
         );
  INV3 U2497 ( .A(n2566), .Q(n2204) );
  AOI211 U2498 ( .A(n2564), .B(\u_cordic/mycordic/present_Q_table[5][5] ), .C(
        n2205), .Q(n2566) );
  OAI2111 U2499 ( .A(\u_coder/n226 ), .B(n1661), .C(\u_coder/n227 ), .D(
        \u_coder/n228 ), .Q(\u_coder/n337 ) );
  AOI221 U2500 ( .A(\u_coder/n220 ), .B(\u_coder/n239 ), .C(\u_coder/n218 ), 
        .D(\u_coder/n239 ), .Q(\u_coder/n226 ) );
  NAND31 U2501 ( .A(\u_coder/my_clk_10M ), .B(\u_coder/n236 ), .C(
        \u_coder/stateQ[0] ), .Q(\u_coder/n227 ) );
  NAND22 U2502 ( .A(sig_coder_outSinQ[0]), .B(n1472), .Q(\u_coder/n228 ) );
  OAI2111 U2503 ( .A(\u_coder/n182 ), .B(n1660), .C(\u_coder/n183 ), .D(
        \u_coder/n184 ), .Q(\u_coder/n334 ) );
  AOI221 U2504 ( .A(\u_coder/n154 ), .B(\u_coder/n194 ), .C(\u_coder/n168 ), 
        .D(\u_coder/n194 ), .Q(\u_coder/n182 ) );
  NAND31 U2505 ( .A(\u_coder/stateI[0] ), .B(\u_coder/n192 ), .C(
        \u_coder/my_clk_10M ), .Q(\u_coder/n183 ) );
  NAND22 U2506 ( .A(sig_coder_outSinI[0]), .B(n1589), .Q(\u_coder/n184 ) );
  INV3 U2507 ( .A(n2571), .Q(n2210) );
  INV3 U2508 ( .A(\u_coder/N1021 ), .Q(n1738) );
  INV3 U2509 ( .A(\u_coder/N1020 ), .Q(n1739) );
  INV3 U2510 ( .A(\u_coder/N1019 ), .Q(n1740) );
  INV3 U2511 ( .A(\u_coder/N1018 ), .Q(n1741) );
  INV3 U2512 ( .A(\u_coder/N1017 ), .Q(n1742) );
  INV3 U2513 ( .A(\u_coder/N1016 ), .Q(n1743) );
  INV3 U2514 ( .A(\u_coder/N1015 ), .Q(n1744) );
  INV3 U2515 ( .A(\u_coder/N1014 ), .Q(n1745) );
  NOR21 U2516 ( .A(n385), .B(n303), .Q(\u_cordic/mycordic/add_262/carry [5])
         );
  NOR21 U2517 ( .A(n106), .B(\u_inFIFO/outWriteCount[2] ), .Q(n2267) );
  NOR21 U2518 ( .A(n377), .B(n468), .Q(\u_cordic/mycordic/add_262/carry [8])
         );
  NAND22 U2519 ( .A(\u_coder/n271 ), .B(\u_coder/n272 ), .Q(\u_coder/n348 ) );
  NAND22 U2520 ( .A(sig_coder_outSinIMasked[0]), .B(\u_coder/n265 ), .Q(
        \u_coder/n271 ) );
  NOR21 U2521 ( .A(\u_cordic/mycordic/present_I_table[4][3] ), .B(n2214), .Q(
        n2583) );
  INV3 U2522 ( .A(n2584), .Q(n2214) );
  AOI211 U2523 ( .A(\u_coder/n266 ), .B(\u_coder/n141 ), .C(n1653), .Q(
        \u_coder/n263 ) );
  NAND22 U2524 ( .A(sig_coder_outSinIMasked[3]), .B(\u_coder/n265 ), .Q(
        \u_coder/n264 ) );
  AOI211 U2525 ( .A(\u_coder/n247 ), .B(\u_coder/n144 ), .C(n1655), .Q(
        \u_coder/n244 ) );
  NAND22 U2526 ( .A(sig_coder_outSinQMasked[3]), .B(\u_coder/n246 ), .Q(
        \u_coder/n245 ) );
  NOR21 U2527 ( .A(n169), .B(n469), .Q(\u_cordic/mycordic/add_262/carry [10])
         );
  NOR21 U2528 ( .A(n200), .B(n541), .Q(\u_cordic/mycordic/add_262/carry [11])
         );
  INV3 U2529 ( .A(\u_cordic/mycordic/add_262/carry [10]), .Q(n541) );
  NOR21 U2530 ( .A(n234), .B(n542), .Q(\u_cordic/mycordic/add_262/carry [12])
         );
  INV3 U2531 ( .A(\u_cordic/mycordic/add_262/carry [11]), .Q(n542) );
  NOR21 U2532 ( .A(n235), .B(n543), .Q(\u_cordic/mycordic/add_262/carry [13])
         );
  INV3 U2533 ( .A(\u_cordic/mycordic/add_262/carry [12]), .Q(n543) );
  NOR21 U2534 ( .A(n260), .B(n544), .Q(\u_cordic/mycordic/add_262/carry [14])
         );
  INV3 U2535 ( .A(\u_cordic/mycordic/add_262/carry [13]), .Q(n544) );
  XOR21 U2536 ( .A(\u_cordic/mycordic/present_ANGLE_table[6][15] ), .B(
        \u_cordic/mycordic/add_262/carry [15]), .Q(\u_cordic/mycordic/N630 )
         );
  NOR21 U2537 ( .A(n279), .B(n545), .Q(\u_cordic/mycordic/add_262/carry [15])
         );
  XOR21 U2538 ( .A(\u_cordic/mycordic/add_262/carry [13]), .B(
        \u_cordic/mycordic/present_ANGLE_table[6][13] ), .Q(
        \u_cordic/mycordic/N628 ) );
  XOR21 U2539 ( .A(\u_cordic/mycordic/add_262/carry [14]), .B(
        \u_cordic/mycordic/present_ANGLE_table[6][14] ), .Q(
        \u_cordic/mycordic/N629 ) );
  NOR21 U2540 ( .A(n158), .B(n209), .Q(\u_cordic/mycordic/add_200/carry [1])
         );
  NOR21 U2541 ( .A(n157), .B(n210), .Q(\u_cordic/mycordic/add_206/carry [1])
         );
  NOR21 U2542 ( .A(n159), .B(n178), .Q(\u_cordic/mycordic/add_189/carry [1])
         );
  NOR21 U2543 ( .A(n160), .B(n211), .Q(\u_cordic/mycordic/add_195/carry [1])
         );
  NOR21 U2544 ( .A(n155), .B(n212), .Q(\u_cordic/mycordic/add_217/carry [1])
         );
  INV3 U2545 ( .A(n2590), .Q(n2217) );
  AOI211 U2546 ( .A(n2589), .B(\u_cordic/mycordic/present_I_table[4][3] ), .C(
        n2218), .Q(n2590) );
  INV3 U2547 ( .A(n2588), .Q(n2218) );
  INV3 U2548 ( .A(n413), .Q(\u_cordic/mycordic/sub_205/carry [1]) );
  NOR21 U2549 ( .A(n158), .B(\u_cordic/mycordic/present_I_table[3][0] ), .Q(
        n413) );
  INV3 U2550 ( .A(n410), .Q(\u_cordic/mycordic/sub_201/carry [1]) );
  NOR21 U2551 ( .A(n157), .B(\u_cordic/mycordic/present_Q_table[3][0] ), .Q(
        n410) );
  INV3 U2552 ( .A(n398), .Q(\u_cordic/mycordic/sub_194/carry [1]) );
  NOR21 U2553 ( .A(n159), .B(\u_cordic/mycordic/present_I_table[2][0] ), .Q(
        n398) );
  INV3 U2554 ( .A(n394), .Q(\u_cordic/mycordic/sub_190/carry [1]) );
  NOR21 U2555 ( .A(n160), .B(\u_cordic/mycordic/present_Q_table[2][0] ), .Q(
        n394) );
  INV3 U2556 ( .A(n425), .Q(\u_cordic/mycordic/sub_212/carry [1]) );
  NOR21 U2557 ( .A(n155), .B(\u_cordic/mycordic/present_Q_table[4][0] ), .Q(
        n425) );
  INV3 U2558 ( .A(n472), .Q(\u_inFIFO/r96/carry [1]) );
  NOR21 U2559 ( .A(n105), .B(\u_inFIFO/outWriteCount[0] ), .Q(n472) );
  INV3 U2560 ( .A(n471), .Q(\u_outFIFO/r98/carry [1]) );
  NOR21 U2561 ( .A(n154), .B(\u_outFIFO/outWriteCount[0] ), .Q(n471) );
  NAND22 U2562 ( .A(\u_cordic/mycordic/present_I_table[5][4] ), .B(n150), .Q(
        n2568) );
  NAND22 U2563 ( .A(\u_decoder/fir_filter/I_data_mult_2_buff [7]), .B(n922), 
        .Q(\u_decoder/fir_filter/n1109 ) );
  NAND22 U2564 ( .A(\u_decoder/fir_filter/I_data_mult_3_buff [7]), .B(n922), 
        .Q(\u_decoder/fir_filter/n1093 ) );
  NAND22 U2565 ( .A(\u_decoder/fir_filter/I_data_mult_5_buff [7]), .B(n921), 
        .Q(\u_decoder/fir_filter/n1061 ) );
  NAND22 U2566 ( .A(\u_decoder/fir_filter/I_data_mult_6_buff [7]), .B(n920), 
        .Q(\u_decoder/fir_filter/n1044 ) );
  NAND22 U2567 ( .A(\u_decoder/fir_filter/Q_data_mult_2_buff [7]), .B(n913), 
        .Q(\u_decoder/fir_filter/n812 ) );
  NAND22 U2568 ( .A(\u_decoder/fir_filter/Q_data_mult_3_buff [7]), .B(n917), 
        .Q(\u_decoder/fir_filter/n796 ) );
  NAND22 U2569 ( .A(\u_decoder/fir_filter/Q_data_mult_5_buff [7]), .B(n918), 
        .Q(\u_decoder/fir_filter/n764 ) );
  NAND22 U2570 ( .A(\u_decoder/fir_filter/Q_data_mult_6_buff [7]), .B(n918), 
        .Q(\u_decoder/fir_filter/n747 ) );
  NAND22 U2571 ( .A(\u_decoder/fir_filter/I_data_mult_0_buff [7]), .B(n916), 
        .Q(\u_decoder/fir_filter/n1141 ) );
  NAND22 U2572 ( .A(\u_decoder/fir_filter/Q_data_mult_0_buff [7]), .B(n926), 
        .Q(\u_decoder/fir_filter/n844 ) );
  NOR21 U2573 ( .A(n167), .B(\u_cordic/mycordic/present_I_table[4][0] ), .Q(
        n2580) );
  AOI221 U2574 ( .A(n2582), .B(\u_cordic/mycordic/present_I_table[4][2] ), .C(
        n231), .D(n2215), .Q(n2584) );
  INV3 U2575 ( .A(n2581), .Q(n2215) );
  NOR21 U2576 ( .A(\u_cordic/mycordic/present_I_table[4][2] ), .B(n2582), .Q(
        n2581) );
  INV3 U2577 ( .A(n2567), .Q(n2213) );
  NOR21 U2578 ( .A(\u_cordic/mycordic/present_Q_table[5][1] ), .B(n2568), .Q(
        n2567) );
  INV3 U2579 ( .A(n467), .Q(\u_cordic/mycordic/add_262/carry [6]) );
  NOR21 U2580 ( .A(\u_cordic/mycordic/present_ANGLE_table[6][5] ), .B(
        \u_cordic/mycordic/add_262/carry [5]), .Q(n467) );
  INV3 U2581 ( .A(\u_cordic/my_rotation/n98 ), .Q(n2230) );
  AOI221 U2582 ( .A(\u_cordic/my_rotation/present_delta [13]), .B(n33), .C(
        \u_cordic/my_rotation/N54 ), .D(n748), .Q(\u_cordic/my_rotation/n98 )
         );
  XOR21 U2583 ( .A(\u_cordic/my_rotation/present_delta [13]), .B(
        \u_cordic/my_rotation/add_43/carry [13]), .Q(
        \u_cordic/my_rotation/N54 ) );
  INV3 U2584 ( .A(\u_cordic/my_rotation/n105 ), .Q(n2236) );
  AOI221 U2585 ( .A(\u_cordic/my_rotation/present_delta [12]), .B(n33), .C(
        \u_cordic/my_rotation/N53 ), .D(n747), .Q(\u_cordic/my_rotation/n105 )
         );
  XOR21 U2586 ( .A(\u_cordic/my_rotation/present_delta [12]), .B(
        \u_cordic/my_rotation/add_43/carry [12]), .Q(
        \u_cordic/my_rotation/N53 ) );
  INV3 U2587 ( .A(n468), .Q(\u_cordic/mycordic/add_262/carry [7]) );
  NOR21 U2588 ( .A(\u_cordic/mycordic/present_ANGLE_table[6][6] ), .B(
        \u_cordic/mycordic/add_262/carry [6]), .Q(n468) );
  INV3 U2589 ( .A(n469), .Q(\u_cordic/mycordic/add_262/carry [9]) );
  NOR21 U2590 ( .A(\u_cordic/mycordic/present_ANGLE_table[6][8] ), .B(
        \u_cordic/mycordic/add_262/carry [8]), .Q(n469) );
  NAND22 U2591 ( .A(\u_coder/n248 ), .B(\u_coder/n249 ), .Q(\u_coder/n340 ) );
  NAND22 U2592 ( .A(sig_coder_outSinQMasked[2]), .B(\u_coder/n246 ), .Q(
        \u_coder/n249 ) );
  NAND22 U2593 ( .A(\u_coder/n248 ), .B(\u_coder/n250 ), .Q(\u_coder/n341 ) );
  NAND22 U2594 ( .A(sig_coder_outSinQMasked[1]), .B(\u_coder/n246 ), .Q(
        \u_coder/n250 ) );
  NAND22 U2595 ( .A(\u_coder/n267 ), .B(\u_coder/n268 ), .Q(\u_coder/n346 ) );
  NAND22 U2596 ( .A(sig_coder_outSinIMasked[2]), .B(\u_coder/n265 ), .Q(
        \u_coder/n268 ) );
  NAND22 U2597 ( .A(\u_coder/n267 ), .B(\u_coder/n269 ), .Q(\u_coder/n347 ) );
  NAND22 U2598 ( .A(sig_coder_outSinIMasked[1]), .B(\u_coder/n265 ), .Q(
        \u_coder/n269 ) );
  NAND22 U2599 ( .A(\u_coder/n252 ), .B(\u_coder/n253 ), .Q(\u_coder/n342 ) );
  NAND22 U2600 ( .A(sig_coder_outSinQMasked[0]), .B(\u_coder/n246 ), .Q(
        \u_coder/n252 ) );
  INV3 U2601 ( .A(n2559), .Q(n2209) );
  INV3 U2602 ( .A(n2563), .Q(n2205) );
  INV3 U2603 ( .A(n2609), .Q(n2241) );
  AOI221 U2604 ( .A(n276), .B(n2608), .C(n2608), .D(n1142), .Q(n2609) );
  NAND22 U2605 ( .A(\u_coder/n202 ), .B(\u_coder/n203 ), .Q(\u_coder/n335 ) );
  AOI221 U2606 ( .A(n1756), .B(\u_coder/n204 ), .C(\u_coder/n205 ), .D(
        \u_coder/n206 ), .Q(\u_coder/n202 ) );
  NAND22 U2607 ( .A(sig_coder_outSinQ[2]), .B(n1472), .Q(\u_coder/n203 ) );
  NAND22 U2608 ( .A(\u_coder/n213 ), .B(\u_coder/n214 ), .Q(\u_coder/n336 ) );
  AOI221 U2609 ( .A(n1756), .B(\u_coder/n215 ), .C(\u_coder/n205 ), .D(
        \u_coder/n216 ), .Q(\u_coder/n213 ) );
  NAND22 U2610 ( .A(sig_coder_outSinQ[1]), .B(n1472), .Q(\u_coder/n214 ) );
  INV3 U2611 ( .A(n2575), .Q(n2206) );
  INV3 U2612 ( .A(n2573), .Q(n2207) );
  AOI211 U2613 ( .A(n217), .B(n2574), .C(
        \u_cordic/mycordic/present_I_table[5][7] ), .Q(n2573) );
  AOI211 U2614 ( .A(n2572), .B(\u_cordic/mycordic/present_Q_table[5][3] ), .C(
        n2210), .Q(n2574) );
  INV3 U2615 ( .A(n2577), .Q(n2203) );
  AOI211 U2616 ( .A(n269), .B(n2578), .C(
        \u_cordic/mycordic/present_I_table[5][7] ), .Q(n2577) );
  AOI211 U2617 ( .A(n2576), .B(\u_cordic/mycordic/present_Q_table[5][5] ), .C(
        n2206), .Q(n2578) );
  XNR21 U2618 ( .A(\u_cordic/mycordic/r173/carry [12]), .B(
        \u_cordic/mycordic/present_ANGLE_table[6][12] ), .Q(n370) );
  XNR21 U2619 ( .A(\u_cordic/mycordic/r173/carry [13]), .B(
        \u_cordic/mycordic/present_ANGLE_table[6][13] ), .Q(n371) );
  XNR21 U2620 ( .A(\u_cordic/mycordic/r173/carry [14]), .B(
        \u_cordic/mycordic/present_ANGLE_table[6][14] ), .Q(n372) );
  INV3 U2621 ( .A(\u_cordic/mycordic/n367 ), .Q(n1311) );
  AOI221 U2622 ( .A(\u_cordic/mycordic/N387 ), .B(n832), .C(
        \u_cordic/mycordic/N419 ), .D(n1582), .Q(\u_cordic/mycordic/n367 ) );
  INV3 U2623 ( .A(\u_cordic/mycordic/n549 ), .Q(n1287) );
  AOI221 U2624 ( .A(\u_cordic/mycordic/N395 ), .B(n831), .C(
        \u_cordic/mycordic/N427 ), .D(n1582), .Q(\u_cordic/mycordic/n549 ) );
  INV3 U2625 ( .A(\u_cordic/mycordic/n491 ), .Q(n1300) );
  AOI221 U2626 ( .A(\u_cordic/mycordic/N408 ), .B(n832), .C(
        \u_cordic/mycordic/N440 ), .D(n1582), .Q(\u_cordic/mycordic/n491 ) );
  XOR21 U2627 ( .A(\u_cordic/mycordic/present_ANGLE_table[2][12] ), .B(
        \u_cordic/mycordic/add_202/carry [12]), .Q(\u_cordic/mycordic/N408 )
         );
  XNR21 U2628 ( .A(\u_cordic/mycordic/present_ANGLE_table[2][12] ), .B(
        \u_cordic/mycordic/sub_207/carry [12]), .Q(\u_cordic/mycordic/N440 )
         );
  INV3 U2629 ( .A(\u_cordic/mycordic/n490 ), .Q(n1301) );
  AOI221 U2630 ( .A(\u_cordic/mycordic/N409 ), .B(n832), .C(
        \u_cordic/mycordic/N441 ), .D(n1582), .Q(\u_cordic/mycordic/n490 ) );
  XOR21 U2631 ( .A(\u_cordic/mycordic/present_ANGLE_table[2][13] ), .B(
        \u_cordic/mycordic/add_202/carry [13]), .Q(\u_cordic/mycordic/N409 )
         );
  XNR21 U2632 ( .A(\u_cordic/mycordic/present_ANGLE_table[2][13] ), .B(
        \u_cordic/mycordic/sub_207/carry [13]), .Q(\u_cordic/mycordic/N441 )
         );
  INV3 U2633 ( .A(\u_cordic/mycordic/n489 ), .Q(n1302) );
  AOI221 U2634 ( .A(\u_cordic/mycordic/N410 ), .B(n831), .C(
        \u_cordic/mycordic/N442 ), .D(n1582), .Q(\u_cordic/mycordic/n489 ) );
  XOR21 U2635 ( .A(\u_cordic/mycordic/present_ANGLE_table[2][14] ), .B(
        \u_cordic/mycordic/add_202/carry [14]), .Q(\u_cordic/mycordic/N410 )
         );
  XNR21 U2636 ( .A(\u_cordic/mycordic/present_ANGLE_table[2][14] ), .B(
        \u_cordic/mycordic/sub_207/carry [14]), .Q(\u_cordic/mycordic/N442 )
         );
  INV3 U2637 ( .A(\u_cordic/mycordic/n375 ), .Q(n1218) );
  AOI221 U2638 ( .A(\u_cordic/mycordic/N323 ), .B(n833), .C(
        \u_cordic/mycordic/N355 ), .D(n1578), .Q(\u_cordic/mycordic/n375 ) );
  INV3 U2639 ( .A(\u_cordic/mycordic/n335 ), .Q(n1226) );
  AOI221 U2640 ( .A(\u_cordic/mycordic/N331 ), .B(n834), .C(
        \u_cordic/mycordic/N363 ), .D(n1578), .Q(\u_cordic/mycordic/n335 ) );
  INV3 U2641 ( .A(\u_cordic/mycordic/n507 ), .Q(n1207) );
  AOI221 U2642 ( .A(\u_cordic/mycordic/N344 ), .B(n833), .C(
        \u_cordic/mycordic/N376 ), .D(n1578), .Q(\u_cordic/mycordic/n507 ) );
  XOR21 U2643 ( .A(\u_cordic/mycordic/present_ANGLE_table[1][12] ), .B(
        \u_cordic/mycordic/add_191/carry[12] ), .Q(\u_cordic/mycordic/N344 )
         );
  XNR21 U2644 ( .A(\u_cordic/mycordic/present_ANGLE_table[1][12] ), .B(
        \u_cordic/mycordic/sub_196/carry[12] ), .Q(\u_cordic/mycordic/N376 )
         );
  INV3 U2645 ( .A(\u_cordic/mycordic/n506 ), .Q(n1208) );
  AOI221 U2646 ( .A(\u_cordic/mycordic/N345 ), .B(n834), .C(
        \u_cordic/mycordic/N377 ), .D(n1578), .Q(\u_cordic/mycordic/n506 ) );
  XOR21 U2647 ( .A(\u_cordic/mycordic/present_ANGLE_table[1][13] ), .B(
        \u_cordic/mycordic/add_191/carry[13] ), .Q(\u_cordic/mycordic/N345 )
         );
  XNR21 U2648 ( .A(\u_cordic/mycordic/present_ANGLE_table[1][13] ), .B(
        \u_cordic/mycordic/sub_196/carry[13] ), .Q(\u_cordic/mycordic/N377 )
         );
  INV3 U2649 ( .A(\u_decoder/fir_filter/n781 ), .Q(n1902) );
  AOI221 U2650 ( .A(\u_decoder/fir_filter/Q_data_mult_4 [8]), .B(n837), .C(
        \u_decoder/fir_filter/Q_data_mult_4_buff [8]), .D(n915), .Q(
        \u_decoder/fir_filter/n781 ) );
  AOI211 U2651 ( .A(n353), .B(n339), .C(n2417), .Q(
        \u_decoder/fir_filter/Q_data_mult_4 [8]) );
  INV3 U2652 ( .A(\u_decoder/fir_filter/n1078 ), .Q(n1831) );
  AOI221 U2653 ( .A(\u_decoder/fir_filter/I_data_mult_4 [8]), .B(n845), .C(
        \u_decoder/fir_filter/I_data_mult_4_buff [8]), .D(n929), .Q(
        \u_decoder/fir_filter/n1078 ) );
  AOI211 U2654 ( .A(n352), .B(n338), .C(n2504), .Q(
        \u_decoder/fir_filter/I_data_mult_4 [8]) );
  INV3 U2655 ( .A(\u_decoder/fir_filter/n988 ), .Q(n2191) );
  AOI221 U2656 ( .A(\u_decoder/fir_filter/I_data_add_7 [8]), .B(n846), .C(
        \u_decoder/fir_filter/I_data_add_7_buff [8]), .D(n930), .Q(
        \u_decoder/fir_filter/n988 ) );
  INV3 U2657 ( .A(\u_decoder/fir_filter/n967 ), .Q(n2176) );
  AOI221 U2658 ( .A(\u_decoder/fir_filter/I_data_add_6 [8]), .B(n846), .C(
        \u_decoder/fir_filter/I_data_add_6_buff [8]), .D(n931), .Q(
        \u_decoder/fir_filter/n967 ) );
  INV3 U2659 ( .A(\u_decoder/fir_filter/n946 ), .Q(n2161) );
  AOI221 U2660 ( .A(\u_decoder/fir_filter/I_data_add_5 [8]), .B(n847), .C(
        \u_decoder/fir_filter/I_data_add_5_buff [8]), .D(n929), .Q(
        \u_decoder/fir_filter/n946 ) );
  INV3 U2661 ( .A(\u_decoder/fir_filter/n925 ), .Q(n2146) );
  AOI221 U2662 ( .A(\u_decoder/fir_filter/I_data_add_4 [8]), .B(n848), .C(
        \u_decoder/fir_filter/I_data_add_4_buff [8]), .D(n932), .Q(
        \u_decoder/fir_filter/n925 ) );
  INV3 U2663 ( .A(\u_decoder/fir_filter/n904 ), .Q(n2131) );
  AOI221 U2664 ( .A(\u_decoder/fir_filter/I_data_add_3 [8]), .B(n849), .C(
        \u_decoder/fir_filter/I_data_add_3_buff [8]), .D(n915), .Q(
        \u_decoder/fir_filter/n904 ) );
  INV3 U2665 ( .A(\u_decoder/fir_filter/n690 ), .Q(n2071) );
  AOI221 U2666 ( .A(\u_decoder/fir_filter/Q_data_add_7 [8]), .B(n838), .C(
        \u_decoder/fir_filter/Q_data_add_7_buff [8]), .D(n929), .Q(
        \u_decoder/fir_filter/n690 ) );
  INV3 U2667 ( .A(\u_decoder/fir_filter/n669 ), .Q(n2056) );
  AOI221 U2668 ( .A(\u_decoder/fir_filter/Q_data_add_6 [8]), .B(n839), .C(
        \u_decoder/fir_filter/Q_data_add_6_buff [8]), .D(n928), .Q(
        \u_decoder/fir_filter/n669 ) );
  INV3 U2669 ( .A(\u_decoder/fir_filter/n648 ), .Q(n2041) );
  AOI221 U2670 ( .A(\u_decoder/fir_filter/Q_data_add_5 [8]), .B(n840), .C(
        \u_decoder/fir_filter/Q_data_add_5_buff [8]), .D(n929), .Q(
        \u_decoder/fir_filter/n648 ) );
  INV3 U2671 ( .A(\u_decoder/fir_filter/n627 ), .Q(n2026) );
  AOI221 U2672 ( .A(\u_decoder/fir_filter/Q_data_add_4 [8]), .B(n841), .C(
        \u_decoder/fir_filter/Q_data_add_4_buff [8]), .D(n926), .Q(
        \u_decoder/fir_filter/n627 ) );
  INV3 U2673 ( .A(\u_decoder/fir_filter/n606 ), .Q(n2011) );
  AOI221 U2674 ( .A(\u_decoder/fir_filter/Q_data_add_3 [8]), .B(n842), .C(
        \u_decoder/fir_filter/Q_data_add_3_buff [8]), .D(n925), .Q(
        \u_decoder/fir_filter/n606 ) );
  INV3 U2675 ( .A(\u_decoder/fir_filter/n585 ), .Q(n1996) );
  AOI221 U2676 ( .A(\u_decoder/fir_filter/Q_data_add_2 [8]), .B(n843), .C(
        \u_decoder/fir_filter/Q_data_add_2_buff [8]), .D(n925), .Q(
        \u_decoder/fir_filter/n585 ) );
  INV3 U2677 ( .A(\u_decoder/fir_filter/n564 ), .Q(n1974) );
  AOI221 U2678 ( .A(\u_decoder/fir_filter/Q_data_add_1 [8]), .B(n844), .C(
        \u_decoder/fir_filter/Q_data_add_1_buff [8]), .D(n931), .Q(
        \u_decoder/fir_filter/n564 ) );
  INV3 U2679 ( .A(\u_decoder/fir_filter/n883 ), .Q(n2116) );
  AOI221 U2680 ( .A(\u_decoder/fir_filter/I_data_add_2 [8]), .B(n850), .C(
        \u_decoder/fir_filter/I_data_add_2_buff [8]), .D(n923), .Q(
        \u_decoder/fir_filter/n883 ) );
  INV3 U2681 ( .A(\u_decoder/fir_filter/n862 ), .Q(n2094) );
  AOI221 U2682 ( .A(\u_decoder/fir_filter/I_data_add_1 [8]), .B(n851), .C(
        \u_decoder/fir_filter/I_data_add_1_buff [8]), .D(n927), .Q(
        \u_decoder/fir_filter/n862 ) );
  INV3 U2683 ( .A(\u_cordic/mycordic/n362 ), .Q(n1282) );
  AOI221 U2684 ( .A(\u_cordic/mycordic/N447 ), .B(n836), .C(
        \u_cordic/mycordic/N475 ), .D(n1581), .Q(\u_cordic/mycordic/n362 ) );
  INV3 U2685 ( .A(\u_cordic/mycordic/n540 ), .Q(n1262) );
  AOI221 U2686 ( .A(\u_cordic/mycordic/N455 ), .B(n835), .C(
        \u_cordic/mycordic/N483 ), .D(n1581), .Q(\u_cordic/mycordic/n540 ) );
  INV3 U2687 ( .A(\u_cordic/mycordic/n476 ), .Q(n1274) );
  AOI221 U2688 ( .A(\u_cordic/mycordic/N467 ), .B(n836), .C(
        \u_cordic/mycordic/N495 ), .D(n1581), .Q(\u_cordic/mycordic/n476 ) );
  XOR21 U2689 ( .A(\u_cordic/mycordic/present_ANGLE_table[3][11] ), .B(
        \u_cordic/mycordic/add_213/carry[11] ), .Q(\u_cordic/mycordic/N467 )
         );
  XNR21 U2690 ( .A(\u_cordic/mycordic/present_ANGLE_table[3][11] ), .B(
        \u_cordic/mycordic/sub_218/carry[11] ), .Q(\u_cordic/mycordic/N495 )
         );
  INV3 U2691 ( .A(\u_cordic/mycordic/n475 ), .Q(n1275) );
  AOI221 U2692 ( .A(\u_cordic/mycordic/N468 ), .B(n836), .C(
        \u_cordic/mycordic/N496 ), .D(n1581), .Q(\u_cordic/mycordic/n475 ) );
  XOR21 U2693 ( .A(\u_cordic/mycordic/present_ANGLE_table[3][12] ), .B(
        \u_cordic/mycordic/add_213/carry[12] ), .Q(\u_cordic/mycordic/N468 )
         );
  XNR21 U2694 ( .A(\u_cordic/mycordic/present_ANGLE_table[3][12] ), .B(
        \u_cordic/mycordic/sub_218/carry[12] ), .Q(\u_cordic/mycordic/N496 )
         );
  INV3 U2695 ( .A(\u_cordic/mycordic/n474 ), .Q(n1276) );
  AOI221 U2696 ( .A(\u_cordic/mycordic/N469 ), .B(n836), .C(
        \u_cordic/mycordic/N497 ), .D(n1581), .Q(\u_cordic/mycordic/n474 ) );
  XOR21 U2697 ( .A(\u_cordic/mycordic/present_ANGLE_table[3][13] ), .B(
        \u_cordic/mycordic/add_213/carry[13] ), .Q(\u_cordic/mycordic/N469 )
         );
  XNR21 U2698 ( .A(\u_cordic/mycordic/present_ANGLE_table[3][13] ), .B(
        \u_cordic/mycordic/sub_218/carry[13] ), .Q(\u_cordic/mycordic/N497 )
         );
  INV3 U2699 ( .A(\u_cordic/mycordic/n460 ), .Q(n1250) );
  AOI221 U2700 ( .A(\u_cordic/mycordic/N512 ), .B(n789), .C(
        \u_cordic/mycordic/N529 ), .D(n1580), .Q(\u_cordic/mycordic/n460 ) );
  XOR21 U2701 ( .A(\u_cordic/mycordic/present_ANGLE_table[4][11] ), .B(
        \u_cordic/mycordic/add_224/carry[11] ), .Q(\u_cordic/mycordic/N512 )
         );
  XNR21 U2702 ( .A(\u_cordic/mycordic/present_ANGLE_table[4][11] ), .B(
        \u_cordic/mycordic/sub_229/carry[11] ), .Q(\u_cordic/mycordic/N529 )
         );
  INV3 U2703 ( .A(\u_cordic/mycordic/n459 ), .Q(n1251) );
  AOI221 U2704 ( .A(\u_cordic/mycordic/N513 ), .B(n789), .C(
        \u_cordic/mycordic/N530 ), .D(n1580), .Q(\u_cordic/mycordic/n459 ) );
  XOR21 U2705 ( .A(\u_cordic/mycordic/present_ANGLE_table[4][12] ), .B(
        \u_cordic/mycordic/add_224/carry[12] ), .Q(\u_cordic/mycordic/N513 )
         );
  XNR21 U2706 ( .A(\u_cordic/mycordic/present_ANGLE_table[4][12] ), .B(
        \u_cordic/mycordic/sub_229/carry[12] ), .Q(\u_cordic/mycordic/N530 )
         );
  INV3 U2707 ( .A(\u_cordic/mycordic/n441 ), .Q(n1191) );
  AOI221 U2708 ( .A(\u_cordic/mycordic/N546 ), .B(n786), .C(
        \u_cordic/mycordic/N562 ), .D(n1577), .Q(\u_cordic/mycordic/n441 ) );
  XOR21 U2709 ( .A(\u_cordic/mycordic/present_ANGLE_table[5][12] ), .B(
        \u_cordic/mycordic/add_233/carry [12]), .Q(\u_cordic/mycordic/N546 )
         );
  XNR21 U2710 ( .A(\u_cordic/mycordic/present_ANGLE_table[5][12] ), .B(
        \u_cordic/mycordic/sub_236/carry [12]), .Q(\u_cordic/mycordic/N562 )
         );
  INV3 U2711 ( .A(\u_cordic/mycordic/n440 ), .Q(n1192) );
  AOI221 U2712 ( .A(\u_cordic/mycordic/N547 ), .B(n786), .C(
        \u_cordic/mycordic/N563 ), .D(n1577), .Q(\u_cordic/mycordic/n440 ) );
  XOR21 U2713 ( .A(\u_cordic/mycordic/present_ANGLE_table[5][13] ), .B(
        \u_cordic/mycordic/add_233/carry [13]), .Q(\u_cordic/mycordic/N547 )
         );
  XNR21 U2714 ( .A(\u_cordic/mycordic/present_ANGLE_table[5][13] ), .B(
        \u_cordic/mycordic/sub_236/carry [13]), .Q(\u_cordic/mycordic/N563 )
         );
  INV3 U2715 ( .A(\u_coder/n255 ), .Q(n1474) );
  AOI221 U2716 ( .A(\u_coder/sin_was_positiveQ ), .B(\u_coder/n256 ), .C(
        \u_coder/isPositiveQ ), .D(\u_coder/n205 ), .Q(\u_coder/n255 ) );
  INV3 U2717 ( .A(\u_cordic/mycordic/n538 ), .Q(n1238) );
  AOI221 U2718 ( .A(\u_cordic/mycordic/N500 ), .B(n788), .C(
        \u_cordic/mycordic/N517 ), .D(n1580), .Q(\u_cordic/mycordic/n538 ) );
  INV3 U2719 ( .A(\u_coder/N1022 ), .Q(n1737) );
  INV3 U2720 ( .A(\u_coder/n198 ), .Q(n1471) );
  AOI211 U2721 ( .A(n1472), .B(sig_coder_outSinQ[3]), .C(\u_coder/n199 ), .Q(
        \u_coder/n198 ) );
  INV3 U2722 ( .A(\u_coder/n157 ), .Q(n1587) );
  AOI211 U2723 ( .A(sig_coder_outSinI[2]), .B(n1589), .C(\u_coder/n158 ), .Q(
        \u_coder/n157 ) );
  AOI221 U2724 ( .A(\u_coder/n168 ), .B(n1720), .C(\u_coder/n154 ), .D(
        \u_coder/n163 ), .Q(\u_coder/n159 ) );
  INV3 U2725 ( .A(\u_coder/n169 ), .Q(n1588) );
  AOI211 U2726 ( .A(sig_coder_outSinI[1]), .B(n1589), .C(\u_coder/n170 ), .Q(
        \u_coder/n169 ) );
  AOI221 U2727 ( .A(\u_coder/n168 ), .B(\u_coder/n177 ), .C(\u_coder/n154 ), 
        .D(\u_coder/n173 ), .Q(\u_coder/n171 ) );
  INV3 U2728 ( .A(\u_cdr/div1/cnt_div/n50 ), .Q(n1503) );
  NAND22 U2729 ( .A(\u_cdr/div1/cnt_div/N67 ), .B(n975), .Q(
        \u_cdr/div1/cnt_div/n50 ) );
  NOR40 U2730 ( .A(n1120), .B(n1119), .C(n1118), .D(n1117), .Q(
        \u_cdr/div1/cnt_div/N67 ) );
  INV3 U2731 ( .A(\u_cordic/mycordic/n402 ), .Q(n1545) );
  NAND22 U2732 ( .A(\u_cordic/mycordic/next_ANGLE_table[6][12] ), .B(n972), 
        .Q(\u_cordic/mycordic/n402 ) );
  INV3 U2733 ( .A(\u_cordic/mycordic/n401 ), .Q(n1544) );
  NAND22 U2734 ( .A(\u_cordic/mycordic/next_ANGLE_table[6][13] ), .B(n972), 
        .Q(\u_cordic/mycordic/n401 ) );
  INV3 U2735 ( .A(\u_cordic/mycordic/n400 ), .Q(n1543) );
  NAND22 U2736 ( .A(\u_cordic/mycordic/next_ANGLE_table[6][14] ), .B(n973), 
        .Q(\u_cordic/mycordic/n400 ) );
  AOI311 U2737 ( .A(\u_cdr/div1/w_en_freq_synch ), .B(\u_cdr/w_sT ), .C(
        \u_cdr/div1/n31 ), .D(n987), .Q(n990) );
  NAND41 U2738 ( .A(\u_coder/n325 ), .B(\u_coder/n326 ), .C(\u_coder/n327 ), 
        .D(\u_coder/n328 ), .Q(\u_coder/n262 ) );
  NOR40 U2739 ( .A(\u_coder/j [9]), .B(\u_coder/j [8]), .C(\u_coder/j [7]), 
        .D(\u_coder/j [6]), .Q(\u_coder/n328 ) );
  NOR40 U2740 ( .A(\u_coder/j [5]), .B(\u_coder/j [4]), .C(\u_coder/j [19]), 
        .D(\u_coder/j [18]), .Q(\u_coder/n327 ) );
  NOR40 U2741 ( .A(\u_coder/j [17]), .B(\u_coder/j [16]), .C(\u_coder/j [15]), 
        .D(\u_coder/j [14]), .Q(\u_coder/n326 ) );
  NOR31 U2742 ( .A(\u_coder/i [2]), .B(\u_coder/i [4]), .C(\u_coder/i [3]), 
        .Q(n2295) );
  NAND31 U2743 ( .A(\u_cdr/div1/n7 ), .B(\u_cdr/w_nb_P [4]), .C(n988), .Q(n989) );
  OAI311 U2744 ( .A(n989), .B(\u_cdr/div1/n8 ), .C(\u_cdr/w_nb_P [2]), .D(
        \u_cdr/w_sE ), .Q(n1008) );
  NOR40 U2745 ( .A(\u_coder/j [13]), .B(\u_coder/j [12]), .C(\u_coder/j [11]), 
        .D(\u_coder/j [10]), .Q(\u_coder/n325 ) );
  OAI311 U2746 ( .A(n989), .B(\u_cdr/div1/n9 ), .C(\u_cdr/w_nb_P [3]), .D(
        \u_cdr/phd1/n9 ), .Q(n1003) );
  NOR31 U2747 ( .A(\u_coder/i [7]), .B(\u_coder/i [9]), .C(\u_coder/i [8]), 
        .Q(n2293) );
  OAI2111 U2748 ( .A(n1002), .B(n1016), .C(n1020), .D(n1001), .Q(
        \u_cdr/div1/n34 ) );
  IMUX21 U2749 ( .A(n1000), .B(n999), .S(\u_cdr/w_nb_P [4]), .Q(n1001) );
  OAI2111 U2750 ( .A(n995), .B(n1016), .C(n1020), .D(n994), .Q(
        \u_cdr/div1/n35 ) );
  IMUX21 U2751 ( .A(n993), .B(n992), .S(\u_cdr/w_nb_P [3]), .Q(n994) );
  NOR21 U2752 ( .A(\u_decoder/fir_filter/state [1]), .B(
        \u_decoder/fir_filter/state [0]), .Q(\u_decoder/fir_filter/n1149 ) );
  NOR21 U2753 ( .A(n1718), .B(\u_coder/n141 ), .Q(\u_coder/n176 ) );
  NOR21 U2754 ( .A(n1718), .B(\u_coder/isPositiveI ), .Q(\u_coder/n162 ) );
  NAND22 U2755 ( .A(\u_coder/N1149 ), .B(\u_coder/n76 ), .Q(\u_coder/n313 ) );
  NAND22 U2756 ( .A(\u_coder/N1143 ), .B(\u_coder/n72 ), .Q(\u_coder/n306 ) );
  NAND22 U2757 ( .A(\u_decoder/fir_filter/state [1]), .B(
        \u_decoder/fir_filter/n410 ), .Q(\u_decoder/fir_filter/n1153 ) );
  NOR21 U2758 ( .A(n105), .B(\u_inFIFO/outWriteCount[0] ), .Q(n2263) );
  NAND22 U2759 ( .A(\u_inFIFO/outReadCount[4] ), .B(\u_inFIFO/n82 ), .Q(n2265)
         );
  XOR21 U2760 ( .A(\u_cordic/mycordic/add_262/carry [11]), .B(
        \u_cordic/mycordic/present_ANGLE_table[6][11] ), .Q(
        \u_cordic/mycordic/N626 ) );
  XOR21 U2761 ( .A(\u_cordic/mycordic/add_262/carry [12]), .B(
        \u_cordic/mycordic/present_ANGLE_table[6][12] ), .Q(
        \u_cordic/mycordic/N627 ) );
  AOI221 U2762 ( .A(\u_coder/n154 ), .B(\u_coder/n155 ), .C(n1724), .D(n1654), 
        .Q(\u_coder/n153 ) );
  INV3 U2763 ( .A(\u_coder/n156 ), .Q(n1654) );
  NAND22 U2764 ( .A(\u_inFIFO/outReadCount[3] ), .B(\u_inFIFO/n83 ), .Q(n2266)
         );
  NAND22 U2765 ( .A(\u_decoder/fir_filter/I_data_mult_1_buff [7]), .B(n924), 
        .Q(\u_decoder/fir_filter/n1125 ) );
  NAND22 U2766 ( .A(\u_decoder/fir_filter/I_data_mult_7_buff [7]), .B(n924), 
        .Q(\u_decoder/fir_filter/n1027 ) );
  NAND22 U2767 ( .A(\u_decoder/fir_filter/Q_data_mult_1_buff [7]), .B(n915), 
        .Q(\u_decoder/fir_filter/n828 ) );
  NAND22 U2768 ( .A(\u_decoder/fir_filter/Q_data_mult_7_buff [7]), .B(n917), 
        .Q(\u_decoder/fir_filter/n730 ) );
  NAND22 U2769 ( .A(\u_decoder/fir_filter/I_data_mult_0_buff [6]), .B(n921), 
        .Q(\u_decoder/fir_filter/n1140 ) );
  NAND22 U2770 ( .A(\u_decoder/fir_filter/Q_data_mult_0_buff [6]), .B(n914), 
        .Q(\u_decoder/fir_filter/n843 ) );
  NAND22 U2771 ( .A(\u_decoder/fir_filter/I_data_mult_3_buff [6]), .B(n922), 
        .Q(\u_decoder/fir_filter/n1092 ) );
  NAND22 U2772 ( .A(\u_decoder/fir_filter/I_data_mult_5_buff [6]), .B(n921), 
        .Q(\u_decoder/fir_filter/n1060 ) );
  NAND22 U2773 ( .A(\u_decoder/fir_filter/Q_data_mult_3_buff [6]), .B(n916), 
        .Q(\u_decoder/fir_filter/n795 ) );
  NAND22 U2774 ( .A(\u_decoder/fir_filter/Q_data_mult_5_buff [6]), .B(n918), 
        .Q(\u_decoder/fir_filter/n763 ) );
  INV3 U2775 ( .A(\u_coder/N668 ), .Q(n1718) );
  NAND41 U2776 ( .A(n2300), .B(n2299), .C(n2298), .D(n2297), .Q(\u_coder/N668 ) );
  NOR21 U2777 ( .A(\u_coder/i [10]), .B(n778), .Q(n2300) );
  NOR31 U2778 ( .A(\u_coder/i [11]), .B(\u_coder/i [13]), .C(\u_coder/i [12]), 
        .Q(n2299) );
  AOI211 U2779 ( .A(\u_inFIFO/n231 ), .B(\u_inFIFO/n232 ), .C(n984), .Q(
        \u_inFIFO/N44 ) );
  NAND22 U2780 ( .A(n1700), .B(\u_inFIFO/n233 ), .Q(\u_inFIFO/n232 ) );
  AOI221 U2781 ( .A(\u_inFIFO/currentState [0]), .B(\u_inFIFO/n109 ), .C(
        \u_inFIFO/N249 ), .D(\u_inFIFO/n234 ), .Q(\u_inFIFO/n231 ) );
  AOI211 U2782 ( .A(\u_outFIFO/n535 ), .B(\u_outFIFO/n536 ), .C(n981), .Q(
        \u_outFIFO/N44 ) );
  AOI221 U2783 ( .A(n1787), .B(\u_outFIFO/currentState [1]), .C(n1792), .D(
        \u_outFIFO/n537 ), .Q(\u_outFIFO/n536 ) );
  AOI221 U2784 ( .A(\u_outFIFO/N473 ), .B(\u_outFIFO/n539 ), .C(
        \u_outFIFO/N474 ), .D(\u_outFIFO/n540 ), .Q(\u_outFIFO/n535 ) );
  INV3 U2785 ( .A(\u_outFIFO/n538 ), .Q(n1787) );
  INV3 U2786 ( .A(\u_cordic/my_rotation/n103 ), .Q(n2234) );
  AOI221 U2787 ( .A(\u_cordic/my_rotation/present_delta [10]), .B(n33), .C(
        \u_cordic/my_rotation/N51 ), .D(n747), .Q(\u_cordic/my_rotation/n103 )
         );
  XOR21 U2788 ( .A(\u_cordic/my_rotation/present_delta [10]), .B(
        \u_cordic/my_rotation/add_43/carry [10]), .Q(
        \u_cordic/my_rotation/N51 ) );
  INV3 U2789 ( .A(\u_cordic/my_rotation/n104 ), .Q(n2235) );
  AOI221 U2790 ( .A(\u_cordic/my_rotation/present_delta [11]), .B(n33), .C(
        \u_cordic/my_rotation/N52 ), .D(n747), .Q(\u_cordic/my_rotation/n104 )
         );
  XOR21 U2791 ( .A(\u_cordic/my_rotation/present_delta [11]), .B(
        \u_cordic/my_rotation/add_43/carry [11]), .Q(
        \u_cordic/my_rotation/N52 ) );
  INV3 U2792 ( .A(\u_cordic/my_rotation/n92 ), .Q(n2224) );
  AOI221 U2793 ( .A(\u_cordic/my_rotation/present_delta [9]), .B(n33), .C(
        \u_cordic/my_rotation/N50 ), .D(n748), .Q(\u_cordic/my_rotation/n92 )
         );
  XOR21 U2794 ( .A(\u_cordic/my_rotation/present_delta [9]), .B(
        \u_cordic/my_rotation/add_43/carry [9]), .Q(\u_cordic/my_rotation/N50 ) );
  OAI311 U2795 ( .A(n1018), .B(n1017), .C(\u_cdr/w_sE ), .D(\u_cdr/div1/N34 ), 
        .Q(n1019) );
  NOR40 U2796 ( .A(n2296), .B(n1721), .C(\u_coder/i [1]), .D(\u_coder/i [19]), 
        .Q(n2297) );
  NAND22 U2797 ( .A(n2294), .B(n2293), .Q(n2296) );
  INV3 U2798 ( .A(n2295), .Q(n1721) );
  NOR21 U2799 ( .A(\u_coder/i [6]), .B(\u_coder/i [5]), .Q(n2294) );
  INV3 U2800 ( .A(\u_decoder/fir_filter/n774 ), .Q(n1932) );
  AOI221 U2801 ( .A(\u_decoder/Q_prefilter [1]), .B(n838), .C(
        \u_decoder/fir_filter/Q_data_mult_4_buff [1]), .D(n920), .Q(
        \u_decoder/fir_filter/n774 ) );
  XNR21 U2802 ( .A(\u_cordic/mycordic/r173/carry [10]), .B(
        \u_cordic/mycordic/present_ANGLE_table[6][10] ), .Q(n373) );
  XNR21 U2803 ( .A(\u_cordic/mycordic/r173/carry [11]), .B(
        \u_cordic/mycordic/present_ANGLE_table[6][11] ), .Q(n374) );
  INV3 U2804 ( .A(\u_decoder/fir_filter/n773 ), .Q(n1889) );
  AOI221 U2805 ( .A(n763), .B(n838), .C(
        \u_decoder/fir_filter/Q_data_mult_4_buff [0]), .D(n921), .Q(
        \u_decoder/fir_filter/n773 ) );
  INV3 U2806 ( .A(\u_cordic/mycordic/n493 ), .Q(n1298) );
  AOI221 U2807 ( .A(\u_cordic/mycordic/N406 ), .B(n832), .C(
        \u_cordic/mycordic/N438 ), .D(n1582), .Q(\u_cordic/mycordic/n493 ) );
  XOR21 U2808 ( .A(\u_cordic/mycordic/present_ANGLE_table[2][10] ), .B(
        \u_cordic/mycordic/add_202/carry [10]), .Q(\u_cordic/mycordic/N406 )
         );
  XNR21 U2809 ( .A(\u_cordic/mycordic/present_ANGLE_table[2][10] ), .B(
        \u_cordic/mycordic/sub_207/carry [10]), .Q(\u_cordic/mycordic/N438 )
         );
  INV3 U2810 ( .A(\u_cordic/mycordic/n492 ), .Q(n1299) );
  AOI221 U2811 ( .A(\u_cordic/mycordic/N407 ), .B(n831), .C(
        \u_cordic/mycordic/N439 ), .D(n1582), .Q(\u_cordic/mycordic/n492 ) );
  XOR21 U2812 ( .A(\u_cordic/mycordic/present_ANGLE_table[2][11] ), .B(
        \u_cordic/mycordic/add_202/carry [11]), .Q(\u_cordic/mycordic/N407 )
         );
  XNR21 U2813 ( .A(\u_cordic/mycordic/present_ANGLE_table[2][11] ), .B(
        \u_cordic/mycordic/sub_207/carry [11]), .Q(\u_cordic/mycordic/N439 )
         );
  INV3 U2814 ( .A(\u_cordic/mycordic/n510 ), .Q(n1204) );
  AOI221 U2815 ( .A(\u_cordic/mycordic/N341 ), .B(n833), .C(
        \u_cordic/mycordic/N373 ), .D(n1578), .Q(\u_cordic/mycordic/n510 ) );
  XNR21 U2816 ( .A(\u_cordic/mycordic/present_ANGLE_table[1][9] ), .B(
        \u_cordic/mycordic/sub_196/carry[9] ), .Q(\u_cordic/mycordic/N373 ) );
  XOR21 U2817 ( .A(\u_cordic/mycordic/present_ANGLE_table[1][9] ), .B(
        \u_cordic/mycordic/add_191/carry[9] ), .Q(\u_cordic/mycordic/N341 ) );
  INV3 U2818 ( .A(\u_cordic/mycordic/n509 ), .Q(n1205) );
  AOI221 U2819 ( .A(\u_cordic/mycordic/N342 ), .B(n833), .C(
        \u_cordic/mycordic/N374 ), .D(n1578), .Q(\u_cordic/mycordic/n509 ) );
  XOR21 U2820 ( .A(\u_cordic/mycordic/present_ANGLE_table[1][10] ), .B(
        \u_cordic/mycordic/add_191/carry[10] ), .Q(\u_cordic/mycordic/N342 )
         );
  XNR21 U2821 ( .A(\u_cordic/mycordic/present_ANGLE_table[1][10] ), .B(
        \u_cordic/mycordic/sub_196/carry[10] ), .Q(\u_cordic/mycordic/N374 )
         );
  INV3 U2822 ( .A(\u_cordic/mycordic/n508 ), .Q(n1206) );
  AOI221 U2823 ( .A(\u_cordic/mycordic/N343 ), .B(n833), .C(
        \u_cordic/mycordic/N375 ), .D(n1578), .Q(\u_cordic/mycordic/n508 ) );
  XOR21 U2824 ( .A(\u_cordic/mycordic/present_ANGLE_table[1][11] ), .B(
        \u_cordic/mycordic/add_191/carry[11] ), .Q(\u_cordic/mycordic/N343 )
         );
  XNR21 U2825 ( .A(\u_cordic/mycordic/present_ANGLE_table[1][11] ), .B(
        \u_cordic/mycordic/sub_196/carry[11] ), .Q(\u_cordic/mycordic/N375 )
         );
  INV3 U2826 ( .A(\u_decoder/fir_filter/n780 ), .Q(n1903) );
  AOI221 U2827 ( .A(\u_decoder/fir_filter/Q_data_mult_4 [7]), .B(n837), .C(
        \u_decoder/fir_filter/Q_data_mult_4_buff [7]), .D(n914), .Q(
        \u_decoder/fir_filter/n780 ) );
  XOR21 U2828 ( .A(n962), .B(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/SUMB[7][0] ), .Q(
        \u_decoder/fir_filter/Q_data_mult_4 [7]) );
  INV3 U2829 ( .A(\u_decoder/fir_filter/n779 ), .Q(n1904) );
  AOI221 U2830 ( .A(\u_decoder/fir_filter/Q_data_mult_4 [6]), .B(n837), .C(
        \u_decoder/fir_filter/Q_data_mult_4_buff [6]), .D(n930), .Q(
        \u_decoder/fir_filter/n779 ) );
  INV3 U2831 ( .A(\u_decoder/fir_filter/n775 ), .Q(n1934) );
  AOI221 U2832 ( .A(n760), .B(n838), .C(
        \u_decoder/fir_filter/Q_data_mult_4_buff [2]), .D(n920), .Q(
        \u_decoder/fir_filter/n775 ) );
  INV3 U2833 ( .A(\u_decoder/fir_filter/n1077 ), .Q(n1832) );
  AOI221 U2834 ( .A(\u_decoder/fir_filter/I_data_mult_4 [7]), .B(n845), .C(
        \u_decoder/fir_filter/I_data_mult_4_buff [7]), .D(n929), .Q(
        \u_decoder/fir_filter/n1077 ) );
  XOR21 U2835 ( .A(n960), .B(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/SUMB[7][0] ), .Q(
        \u_decoder/fir_filter/I_data_mult_4 [7]) );
  INV3 U2836 ( .A(\u_decoder/fir_filter/n990 ), .Q(n2193) );
  AOI221 U2837 ( .A(\u_decoder/fir_filter/I_data_add_7 [6]), .B(n845), .C(
        \u_decoder/fir_filter/I_data_add_7_buff [6]), .D(n930), .Q(
        \u_decoder/fir_filter/n990 ) );
  INV3 U2838 ( .A(\u_decoder/fir_filter/n989 ), .Q(n2192) );
  AOI221 U2839 ( .A(\u_decoder/fir_filter/I_data_add_7 [7]), .B(n846), .C(
        \u_decoder/fir_filter/I_data_add_7_buff [7]), .D(n930), .Q(
        \u_decoder/fir_filter/n989 ) );
  INV3 U2840 ( .A(\u_decoder/fir_filter/n969 ), .Q(n2178) );
  AOI221 U2841 ( .A(\u_decoder/fir_filter/I_data_add_6 [6]), .B(n846), .C(
        \u_decoder/fir_filter/I_data_add_6_buff [6]), .D(n931), .Q(
        \u_decoder/fir_filter/n969 ) );
  INV3 U2842 ( .A(\u_decoder/fir_filter/n968 ), .Q(n2177) );
  AOI221 U2843 ( .A(\u_decoder/fir_filter/I_data_add_6 [7]), .B(n846), .C(
        \u_decoder/fir_filter/I_data_add_6_buff [7]), .D(n931), .Q(
        \u_decoder/fir_filter/n968 ) );
  INV3 U2844 ( .A(\u_decoder/fir_filter/n948 ), .Q(n2163) );
  AOI221 U2845 ( .A(\u_decoder/fir_filter/I_data_add_5 [6]), .B(n847), .C(
        \u_decoder/fir_filter/I_data_add_5_buff [6]), .D(n930), .Q(
        \u_decoder/fir_filter/n948 ) );
  INV3 U2846 ( .A(\u_decoder/fir_filter/n947 ), .Q(n2162) );
  AOI221 U2847 ( .A(\u_decoder/fir_filter/I_data_add_5 [7]), .B(n847), .C(
        \u_decoder/fir_filter/I_data_add_5_buff [7]), .D(n931), .Q(
        \u_decoder/fir_filter/n947 ) );
  INV3 U2848 ( .A(\u_decoder/fir_filter/n927 ), .Q(n2148) );
  AOI221 U2849 ( .A(\u_decoder/fir_filter/I_data_add_4 [6]), .B(n848), .C(
        \u_decoder/fir_filter/I_data_add_4_buff [6]), .D(n932), .Q(
        \u_decoder/fir_filter/n927 ) );
  INV3 U2850 ( .A(\u_decoder/fir_filter/n926 ), .Q(n2147) );
  AOI221 U2851 ( .A(\u_decoder/fir_filter/I_data_add_4 [7]), .B(n848), .C(
        \u_decoder/fir_filter/I_data_add_4_buff [7]), .D(n932), .Q(
        \u_decoder/fir_filter/n926 ) );
  INV3 U2852 ( .A(\u_decoder/fir_filter/n906 ), .Q(n2133) );
  AOI221 U2853 ( .A(\u_decoder/fir_filter/I_data_add_3 [6]), .B(n849), .C(
        \u_decoder/fir_filter/I_data_add_3_buff [6]), .D(n914), .Q(
        \u_decoder/fir_filter/n906 ) );
  INV3 U2854 ( .A(\u_decoder/fir_filter/n905 ), .Q(n2132) );
  AOI221 U2855 ( .A(\u_decoder/fir_filter/I_data_add_3 [7]), .B(n849), .C(
        \u_decoder/fir_filter/I_data_add_3_buff [7]), .D(n914), .Q(
        \u_decoder/fir_filter/n905 ) );
  INV3 U2856 ( .A(\u_decoder/fir_filter/n778 ), .Q(n1905) );
  AOI221 U2857 ( .A(\u_decoder/fir_filter/Q_data_mult_4 [5]), .B(n838), .C(
        \u_decoder/fir_filter/Q_data_mult_4_buff [5]), .D(n922), .Q(
        \u_decoder/fir_filter/n778 ) );
  INV3 U2858 ( .A(\u_decoder/fir_filter/n777 ), .Q(n1906) );
  AOI221 U2859 ( .A(\u_decoder/fir_filter/Q_data_mult_4 [4]), .B(n838), .C(
        \u_decoder/fir_filter/Q_data_mult_4_buff [4]), .D(n923), .Q(
        \u_decoder/fir_filter/n777 ) );
  INV3 U2860 ( .A(\u_decoder/fir_filter/n776 ), .Q(n1907) );
  AOI221 U2861 ( .A(\u_decoder/fir_filter/Q_data_mult_4 [3]), .B(n838), .C(
        \u_decoder/fir_filter/Q_data_mult_4_buff [3]), .D(n921), .Q(
        \u_decoder/fir_filter/n776 ) );
  XOR21 U2862 ( .A(n758), .B(n763), .Q(\u_decoder/fir_filter/Q_data_mult_4 [3]) );
  INV3 U2863 ( .A(\u_decoder/fir_filter/n698 ), .Q(n2079) );
  AOI221 U2864 ( .A(\u_decoder/fir_filter/Q_data_add_7 [0]), .B(n838), .C(
        \u_decoder/fir_filter/Q_data_add_7_buff [0]), .D(n925), .Q(
        \u_decoder/fir_filter/n698 ) );
  XOR21 U2865 ( .A(\u_decoder/fir_filter/Q_data_mult_7_buff [0]), .B(
        \u_decoder/fir_filter/Q_data_mult_8_buff [0]), .Q(
        \u_decoder/fir_filter/Q_data_add_7 [0]) );
  INV3 U2866 ( .A(\u_decoder/fir_filter/n697 ), .Q(n2078) );
  AOI221 U2867 ( .A(\u_decoder/fir_filter/Q_data_add_7 [1]), .B(n838), .C(
        \u_decoder/fir_filter/Q_data_add_7_buff [1]), .D(n929), .Q(
        \u_decoder/fir_filter/n697 ) );
  INV3 U2868 ( .A(\u_decoder/fir_filter/n696 ), .Q(n2077) );
  AOI221 U2869 ( .A(\u_decoder/fir_filter/Q_data_add_7 [2]), .B(n838), .C(
        \u_decoder/fir_filter/Q_data_add_7_buff [2]), .D(n929), .Q(
        \u_decoder/fir_filter/n696 ) );
  INV3 U2870 ( .A(\u_decoder/fir_filter/n695 ), .Q(n2076) );
  AOI221 U2871 ( .A(\u_decoder/fir_filter/Q_data_add_7 [3]), .B(n838), .C(
        \u_decoder/fir_filter/Q_data_add_7_buff [3]), .D(n929), .Q(
        \u_decoder/fir_filter/n695 ) );
  INV3 U2872 ( .A(\u_decoder/fir_filter/n694 ), .Q(n2075) );
  AOI221 U2873 ( .A(\u_decoder/fir_filter/Q_data_add_7 [4]), .B(n838), .C(
        \u_decoder/fir_filter/Q_data_add_7_buff [4]), .D(n929), .Q(
        \u_decoder/fir_filter/n694 ) );
  INV3 U2874 ( .A(\u_decoder/fir_filter/n693 ), .Q(n2074) );
  AOI221 U2875 ( .A(\u_decoder/fir_filter/Q_data_add_7 [5]), .B(n838), .C(
        \u_decoder/fir_filter/Q_data_add_7_buff [5]), .D(n929), .Q(
        \u_decoder/fir_filter/n693 ) );
  INV3 U2876 ( .A(\u_decoder/fir_filter/n692 ), .Q(n2073) );
  AOI221 U2877 ( .A(\u_decoder/fir_filter/Q_data_add_7 [6]), .B(n838), .C(
        \u_decoder/fir_filter/Q_data_add_7_buff [6]), .D(n929), .Q(
        \u_decoder/fir_filter/n692 ) );
  INV3 U2878 ( .A(\u_decoder/fir_filter/n691 ), .Q(n2072) );
  AOI221 U2879 ( .A(\u_decoder/fir_filter/Q_data_add_7 [7]), .B(n838), .C(
        \u_decoder/fir_filter/Q_data_add_7_buff [7]), .D(n929), .Q(
        \u_decoder/fir_filter/n691 ) );
  INV3 U2880 ( .A(\u_decoder/fir_filter/n677 ), .Q(n2064) );
  AOI221 U2881 ( .A(\u_decoder/fir_filter/Q_data_add_6 [0]), .B(n839), .C(
        \u_decoder/fir_filter/Q_data_add_6_buff [0]), .D(n928), .Q(
        \u_decoder/fir_filter/n677 ) );
  XOR21 U2882 ( .A(\u_decoder/fir_filter/Q_data_mult_6_buff [0]), .B(
        \u_decoder/fir_filter/Q_data_add_7_buff [0]), .Q(
        \u_decoder/fir_filter/Q_data_add_6 [0]) );
  INV3 U2883 ( .A(\u_decoder/fir_filter/n676 ), .Q(n2063) );
  AOI221 U2884 ( .A(\u_decoder/fir_filter/Q_data_add_6 [1]), .B(n839), .C(
        \u_decoder/fir_filter/Q_data_add_6_buff [1]), .D(n928), .Q(
        \u_decoder/fir_filter/n676 ) );
  INV3 U2885 ( .A(\u_decoder/fir_filter/n675 ), .Q(n2062) );
  AOI221 U2886 ( .A(\u_decoder/fir_filter/Q_data_add_6 [2]), .B(n839), .C(
        \u_decoder/fir_filter/Q_data_add_6_buff [2]), .D(n928), .Q(
        \u_decoder/fir_filter/n675 ) );
  INV3 U2887 ( .A(\u_decoder/fir_filter/n674 ), .Q(n2061) );
  AOI221 U2888 ( .A(\u_decoder/fir_filter/Q_data_add_6 [3]), .B(n839), .C(
        \u_decoder/fir_filter/Q_data_add_6_buff [3]), .D(n928), .Q(
        \u_decoder/fir_filter/n674 ) );
  INV3 U2889 ( .A(\u_decoder/fir_filter/n673 ), .Q(n2060) );
  AOI221 U2890 ( .A(\u_decoder/fir_filter/Q_data_add_6 [4]), .B(n839), .C(
        \u_decoder/fir_filter/Q_data_add_6_buff [4]), .D(n928), .Q(
        \u_decoder/fir_filter/n673 ) );
  INV3 U2891 ( .A(\u_decoder/fir_filter/n672 ), .Q(n2059) );
  AOI221 U2892 ( .A(\u_decoder/fir_filter/Q_data_add_6 [5]), .B(n839), .C(
        \u_decoder/fir_filter/Q_data_add_6_buff [5]), .D(n928), .Q(
        \u_decoder/fir_filter/n672 ) );
  INV3 U2893 ( .A(\u_decoder/fir_filter/n671 ), .Q(n2058) );
  AOI221 U2894 ( .A(\u_decoder/fir_filter/Q_data_add_6 [6]), .B(n839), .C(
        \u_decoder/fir_filter/Q_data_add_6_buff [6]), .D(n928), .Q(
        \u_decoder/fir_filter/n671 ) );
  INV3 U2895 ( .A(\u_decoder/fir_filter/n670 ), .Q(n2057) );
  AOI221 U2896 ( .A(\u_decoder/fir_filter/Q_data_add_6 [7]), .B(n839), .C(
        \u_decoder/fir_filter/Q_data_add_6_buff [7]), .D(n928), .Q(
        \u_decoder/fir_filter/n670 ) );
  INV3 U2897 ( .A(\u_decoder/fir_filter/n656 ), .Q(n2049) );
  AOI221 U2898 ( .A(\u_decoder/fir_filter/Q_data_add_5 [0]), .B(n840), .C(
        \u_decoder/fir_filter/Q_data_add_5_buff [0]), .D(n928), .Q(
        \u_decoder/fir_filter/n656 ) );
  XOR21 U2899 ( .A(\u_decoder/fir_filter/Q_data_mult_5_buff [0]), .B(
        \u_decoder/fir_filter/Q_data_add_6_buff [0]), .Q(
        \u_decoder/fir_filter/Q_data_add_5 [0]) );
  INV3 U2900 ( .A(\u_decoder/fir_filter/n655 ), .Q(n2048) );
  AOI221 U2901 ( .A(\u_decoder/fir_filter/Q_data_add_5 [1]), .B(n840), .C(
        \u_decoder/fir_filter/Q_data_add_5_buff [1]), .D(n930), .Q(
        \u_decoder/fir_filter/n655 ) );
  INV3 U2902 ( .A(\u_decoder/fir_filter/n654 ), .Q(n2047) );
  AOI221 U2903 ( .A(\u_decoder/fir_filter/Q_data_add_5 [2]), .B(n840), .C(
        \u_decoder/fir_filter/Q_data_add_5_buff [2]), .D(n927), .Q(
        \u_decoder/fir_filter/n654 ) );
  INV3 U2904 ( .A(\u_decoder/fir_filter/n653 ), .Q(n2046) );
  AOI221 U2905 ( .A(\u_decoder/fir_filter/Q_data_add_5 [3]), .B(n840), .C(
        \u_decoder/fir_filter/Q_data_add_5_buff [3]), .D(n924), .Q(
        \u_decoder/fir_filter/n653 ) );
  INV3 U2906 ( .A(\u_decoder/fir_filter/n652 ), .Q(n2045) );
  AOI221 U2907 ( .A(\u_decoder/fir_filter/Q_data_add_5 [4]), .B(n840), .C(
        \u_decoder/fir_filter/Q_data_add_5_buff [4]), .D(n922), .Q(
        \u_decoder/fir_filter/n652 ) );
  INV3 U2908 ( .A(\u_decoder/fir_filter/n651 ), .Q(n2044) );
  AOI221 U2909 ( .A(\u_decoder/fir_filter/Q_data_add_5 [5]), .B(n840), .C(
        \u_decoder/fir_filter/Q_data_add_5_buff [5]), .D(n925), .Q(
        \u_decoder/fir_filter/n651 ) );
  INV3 U2910 ( .A(\u_decoder/fir_filter/n650 ), .Q(n2043) );
  AOI221 U2911 ( .A(\u_decoder/fir_filter/Q_data_add_5 [6]), .B(n840), .C(
        \u_decoder/fir_filter/Q_data_add_5_buff [6]), .D(n926), .Q(
        \u_decoder/fir_filter/n650 ) );
  INV3 U2912 ( .A(\u_decoder/fir_filter/n649 ), .Q(n2042) );
  AOI221 U2913 ( .A(\u_decoder/fir_filter/Q_data_add_5 [7]), .B(n840), .C(
        \u_decoder/fir_filter/Q_data_add_5_buff [7]), .D(n928), .Q(
        \u_decoder/fir_filter/n649 ) );
  INV3 U2914 ( .A(\u_decoder/fir_filter/n629 ), .Q(n2028) );
  AOI221 U2915 ( .A(\u_decoder/fir_filter/Q_data_add_4 [6]), .B(n841), .C(
        \u_decoder/fir_filter/Q_data_add_4_buff [6]), .D(n926), .Q(
        \u_decoder/fir_filter/n629 ) );
  INV3 U2916 ( .A(\u_decoder/fir_filter/n628 ), .Q(n2027) );
  AOI221 U2917 ( .A(\u_decoder/fir_filter/Q_data_add_4 [7]), .B(n841), .C(
        \u_decoder/fir_filter/Q_data_add_4_buff [7]), .D(n926), .Q(
        \u_decoder/fir_filter/n628 ) );
  INV3 U2918 ( .A(\u_decoder/fir_filter/n608 ), .Q(n2013) );
  AOI221 U2919 ( .A(\u_decoder/fir_filter/Q_data_add_3 [6]), .B(n842), .C(
        \u_decoder/fir_filter/Q_data_add_3_buff [6]), .D(n926), .Q(
        \u_decoder/fir_filter/n608 ) );
  INV3 U2920 ( .A(\u_decoder/fir_filter/n607 ), .Q(n2012) );
  AOI221 U2921 ( .A(\u_decoder/fir_filter/Q_data_add_3 [7]), .B(n842), .C(
        \u_decoder/fir_filter/Q_data_add_3_buff [7]), .D(n926), .Q(
        \u_decoder/fir_filter/n607 ) );
  INV3 U2922 ( .A(\u_decoder/fir_filter/n587 ), .Q(n1998) );
  AOI221 U2923 ( .A(\u_decoder/fir_filter/Q_data_add_2 [6]), .B(n843), .C(
        \u_decoder/fir_filter/Q_data_add_2_buff [6]), .D(n925), .Q(
        \u_decoder/fir_filter/n587 ) );
  INV3 U2924 ( .A(\u_decoder/fir_filter/n586 ), .Q(n1997) );
  AOI221 U2925 ( .A(\u_decoder/fir_filter/Q_data_add_2 [7]), .B(n843), .C(
        \u_decoder/fir_filter/Q_data_add_2_buff [7]), .D(n925), .Q(
        \u_decoder/fir_filter/n586 ) );
  INV3 U2926 ( .A(\u_decoder/fir_filter/n566 ), .Q(n1978) );
  AOI221 U2927 ( .A(\u_decoder/fir_filter/Q_data_add_1 [6]), .B(n844), .C(
        \u_decoder/fir_filter/Q_data_add_1_buff [6]), .D(n929), .Q(
        \u_decoder/fir_filter/n566 ) );
  INV3 U2928 ( .A(\u_decoder/fir_filter/n565 ), .Q(n1977) );
  AOI221 U2929 ( .A(\u_decoder/fir_filter/Q_data_add_1 [7]), .B(n844), .C(
        \u_decoder/fir_filter/Q_data_add_1_buff [7]), .D(n931), .Q(
        \u_decoder/fir_filter/n565 ) );
  INV3 U2930 ( .A(\u_decoder/fir_filter/n885 ), .Q(n2118) );
  AOI221 U2931 ( .A(\u_decoder/fir_filter/I_data_add_2 [6]), .B(n850), .C(
        \u_decoder/fir_filter/I_data_add_2_buff [6]), .D(n932), .Q(
        \u_decoder/fir_filter/n885 ) );
  INV3 U2932 ( .A(\u_decoder/fir_filter/n884 ), .Q(n2117) );
  AOI221 U2933 ( .A(\u_decoder/fir_filter/I_data_add_2 [7]), .B(n850), .C(
        \u_decoder/fir_filter/I_data_add_2_buff [7]), .D(n922), .Q(
        \u_decoder/fir_filter/n884 ) );
  INV3 U2934 ( .A(\u_decoder/fir_filter/n864 ), .Q(n2098) );
  AOI221 U2935 ( .A(\u_decoder/fir_filter/I_data_add_1 [6]), .B(n851), .C(
        \u_decoder/fir_filter/I_data_add_1_buff [6]), .D(n924), .Q(
        \u_decoder/fir_filter/n864 ) );
  INV3 U2936 ( .A(\u_decoder/fir_filter/n863 ), .Q(n2097) );
  AOI221 U2937 ( .A(\u_decoder/fir_filter/I_data_add_1 [7]), .B(n851), .C(
        \u_decoder/fir_filter/I_data_add_1_buff [7]), .D(n930), .Q(
        \u_decoder/fir_filter/n863 ) );
  INV3 U2938 ( .A(\u_cordic/mycordic/n478 ), .Q(n1272) );
  AOI221 U2939 ( .A(\u_cordic/mycordic/N465 ), .B(n836), .C(
        \u_cordic/mycordic/N493 ), .D(n1581), .Q(\u_cordic/mycordic/n478 ) );
  XOR21 U2940 ( .A(\u_cordic/mycordic/present_ANGLE_table[3][9] ), .B(
        \u_cordic/mycordic/add_213/carry[9] ), .Q(\u_cordic/mycordic/N465 ) );
  XNR21 U2941 ( .A(\u_cordic/mycordic/present_ANGLE_table[3][9] ), .B(
        \u_cordic/mycordic/sub_218/carry[9] ), .Q(\u_cordic/mycordic/N493 ) );
  INV3 U2942 ( .A(\u_cordic/mycordic/n477 ), .Q(n1273) );
  AOI221 U2943 ( .A(\u_cordic/mycordic/N466 ), .B(n836), .C(
        \u_cordic/mycordic/N494 ), .D(n1581), .Q(\u_cordic/mycordic/n477 ) );
  XOR21 U2944 ( .A(\u_cordic/mycordic/present_ANGLE_table[3][10] ), .B(
        \u_cordic/mycordic/add_213/carry[10] ), .Q(\u_cordic/mycordic/N466 )
         );
  XNR21 U2945 ( .A(\u_cordic/mycordic/present_ANGLE_table[3][10] ), .B(
        \u_cordic/mycordic/sub_218/carry[10] ), .Q(\u_cordic/mycordic/N494 )
         );
  INV3 U2946 ( .A(\u_cordic/mycordic/n462 ), .Q(n1248) );
  AOI221 U2947 ( .A(\u_cordic/mycordic/N510 ), .B(n789), .C(
        \u_cordic/mycordic/N527 ), .D(n1580), .Q(\u_cordic/mycordic/n462 ) );
  XOR21 U2948 ( .A(\u_cordic/mycordic/present_ANGLE_table[4][9] ), .B(
        \u_cordic/mycordic/add_224/carry[9] ), .Q(\u_cordic/mycordic/N510 ) );
  XNR21 U2949 ( .A(\u_cordic/mycordic/present_ANGLE_table[4][9] ), .B(
        \u_cordic/mycordic/sub_229/carry[9] ), .Q(\u_cordic/mycordic/N527 ) );
  INV3 U2950 ( .A(\u_cordic/mycordic/n461 ), .Q(n1249) );
  AOI221 U2951 ( .A(\u_cordic/mycordic/N511 ), .B(n789), .C(
        \u_cordic/mycordic/N528 ), .D(n1580), .Q(\u_cordic/mycordic/n461 ) );
  XOR21 U2952 ( .A(\u_cordic/mycordic/present_ANGLE_table[4][10] ), .B(
        \u_cordic/mycordic/add_224/carry[10] ), .Q(\u_cordic/mycordic/N511 )
         );
  XNR21 U2953 ( .A(\u_cordic/mycordic/present_ANGLE_table[4][10] ), .B(
        \u_cordic/mycordic/sub_229/carry[10] ), .Q(\u_cordic/mycordic/N528 )
         );
  INV3 U2954 ( .A(\u_cordic/mycordic/n443 ), .Q(n1189) );
  AOI221 U2955 ( .A(\u_cordic/mycordic/N544 ), .B(n786), .C(
        \u_cordic/mycordic/N560 ), .D(n1577), .Q(\u_cordic/mycordic/n443 ) );
  XOR21 U2956 ( .A(\u_cordic/mycordic/present_ANGLE_table[5][10] ), .B(
        \u_cordic/mycordic/add_233/carry [10]), .Q(\u_cordic/mycordic/N544 )
         );
  XNR21 U2957 ( .A(\u_cordic/mycordic/present_ANGLE_table[5][10] ), .B(
        \u_cordic/mycordic/sub_236/carry [10]), .Q(\u_cordic/mycordic/N560 )
         );
  INV3 U2958 ( .A(\u_cordic/mycordic/n442 ), .Q(n1190) );
  AOI221 U2959 ( .A(\u_cordic/mycordic/N545 ), .B(n786), .C(
        \u_cordic/mycordic/N561 ), .D(n1577), .Q(\u_cordic/mycordic/n442 ) );
  XOR21 U2960 ( .A(\u_cordic/mycordic/present_ANGLE_table[5][11] ), .B(
        \u_cordic/mycordic/add_233/carry [11]), .Q(\u_cordic/mycordic/N545 )
         );
  XNR21 U2961 ( .A(\u_cordic/mycordic/present_ANGLE_table[5][11] ), .B(
        \u_cordic/mycordic/sub_236/carry [11]), .Q(\u_cordic/mycordic/N561 )
         );
  INV3 U2962 ( .A(n2630), .Q(n1491) );
  NAND22 U2963 ( .A(\u_cdr/phd1/cnt_phd/N59 ), .B(n976), .Q(n2630) );
  NOR31 U2964 ( .A(n1066), .B(n1065), .C(n1064), .Q(\u_cdr/phd1/cnt_phd/N59 )
         );
  INV3 U2965 ( .A(\u_cordic/mycordic/n404 ), .Q(n1547) );
  NAND22 U2966 ( .A(\u_cordic/mycordic/next_ANGLE_table[6][10] ), .B(n972), 
        .Q(\u_cordic/mycordic/n404 ) );
  INV3 U2967 ( .A(\u_cordic/mycordic/n403 ), .Q(n1546) );
  NAND22 U2968 ( .A(\u_cordic/mycordic/next_ANGLE_table[6][11] ), .B(n972), 
        .Q(\u_cordic/mycordic/n403 ) );
  NOR31 U2969 ( .A(\u_outFIFO/n195 ), .B(\u_outFIFO/n196 ), .C(
        \u_outFIFO/n544 ), .Q(\u_outFIFO/N178 ) );
  NAND41 U2970 ( .A(\u_coder/n329 ), .B(\u_coder/n330 ), .C(\u_coder/n331 ), 
        .D(\u_coder/n332 ), .Q(\u_coder/n275 ) );
  NOR40 U2971 ( .A(\u_coder/i [9]), .B(\u_coder/i [8]), .C(\u_coder/i [7]), 
        .D(\u_coder/i [6]), .Q(\u_coder/n332 ) );
  NOR40 U2972 ( .A(\u_coder/i [5]), .B(\u_coder/i [4]), .C(\u_coder/i [19]), 
        .D(\u_coder/i [18]), .Q(\u_coder/n331 ) );
  NOR40 U2973 ( .A(\u_coder/i [17]), .B(\u_coder/i [16]), .C(\u_coder/i [15]), 
        .D(\u_coder/i [14]), .Q(\u_coder/n330 ) );
  NAND41 U2974 ( .A(n2291), .B(n2290), .C(n2289), .D(n2288), .Q(\u_coder/N974 ) );
  NOR21 U2975 ( .A(\u_coder/j [10]), .B(n777), .Q(n2291) );
  NOR31 U2976 ( .A(\u_coder/j [11]), .B(\u_coder/j [13]), .C(\u_coder/j [12]), 
        .Q(n2290) );
  NOR40 U2977 ( .A(\u_coder/j [16]), .B(n1755), .C(\u_coder/j [15]), .D(
        \u_coder/j [14]), .Q(n2289) );
  NOR31 U2978 ( .A(\u_outFIFO/n531 ), .B(\u_outFIFO/n206 ), .C(n1468), .Q(
        \u_outFIFO/n527 ) );
  NOR40 U2979 ( .A(\u_outFIFO/outWriteCount[0] ), .B(
        \u_outFIFO/outWriteCount[1] ), .C(\u_outFIFO/n178 ), .D(
        \u_outFIFO/n532 ), .Q(\u_outFIFO/n531 ) );
  NAND31 U2980 ( .A(\u_outFIFO/n182 ), .B(\u_outFIFO/n180 ), .C(
        \u_outFIFO/n181 ), .Q(\u_outFIFO/n532 ) );
  NOR31 U2981 ( .A(\u_coder/n86 ), .B(\u_coder/n275 ), .C(\u_coder/n312 ), .Q(
        \u_coder/n266 ) );
  NAND31 U2982 ( .A(\u_coder/n89 ), .B(\u_coder/n85 ), .C(\u_coder/n88 ), .Q(
        \u_coder/n312 ) );
  NOR31 U2983 ( .A(\u_coder/n275 ), .B(n1720), .C(\u_coder/n89 ), .Q(
        \u_coder/n281 ) );
  NOR31 U2984 ( .A(\u_coder/n135 ), .B(\u_coder/n262 ), .C(\u_coder/n311 ), 
        .Q(\u_coder/n247 ) );
  NAND31 U2985 ( .A(\u_coder/n138 ), .B(\u_coder/n134 ), .C(\u_coder/n137 ), 
        .Q(\u_coder/n311 ) );
  AOI221 U2986 ( .A(\u_cordic/my_rotation/present_delta [7]), .B(n33), .C(
        \u_cordic/my_rotation/N48 ), .D(n748), .Q(\u_cordic/my_rotation/n63 )
         );
  XOR21 U2987 ( .A(\u_cordic/my_rotation/present_delta [7]), .B(
        \u_cordic/my_rotation/add_43/carry [7]), .Q(\u_cordic/my_rotation/N48 ) );
  AOI221 U2988 ( .A(\sig_MUX_inMUX4[0] ), .B(n1687), .C(in_MUX_inSEL3), .D(
        sig_DEMUX_outDEMUX1[1]), .Q(n2687) );
  NOR31 U2989 ( .A(\u_demux1/n4 ), .B(in_DEMUX_inSEL1[2]), .C(
        in_DEMUX_inSEL1[1]), .Q(sig_DEMUX_outDEMUX1[1]) );
  NAND41 U2990 ( .A(n976), .B(\u_cdr/div1/w_en_freq_synch ), .C(\u_cdr/w_sT ), 
        .D(\u_cdr/div1/n31 ), .Q(\u_cdr/div1/n30 ) );
  NOR40 U2991 ( .A(\u_coder/i [13]), .B(\u_coder/i [12]), .C(\u_coder/i [11]), 
        .D(\u_coder/i [10]), .Q(\u_coder/n329 ) );
  NOR21 U2992 ( .A(\u_outFIFO/n538 ), .B(\u_outFIFO/currentState [0]), .Q(
        \u_outFIFO/n206 ) );
  NAND31 U2993 ( .A(\u_coder/n89 ), .B(\u_coder/n85 ), .C(\u_coder/n165 ), .Q(
        \u_coder/n178 ) );
  NOR31 U2994 ( .A(\u_coder/j [2]), .B(\u_coder/j [4]), .C(n776), .Q(n2286) );
  AOI221 U2995 ( .A(n1724), .B(n1653), .C(\u_coder/isPositiveI ), .D(n1714), 
        .Q(\u_coder/n267 ) );
  AOI221 U2996 ( .A(\u_outFIFO/N136 ), .B(n1467), .C(\u_outFIFO/N118 ), .D(
        \u_outFIFO/n514 ), .Q(\u_outFIFO/n528 ) );
  XOR21 U2997 ( .A(\u_outFIFO/add_255/carry [5]), .B(
        \u_outFIFO/outWriteCount[5] ), .Q(\u_outFIFO/N118 ) );
  AOI221 U2998 ( .A(\u_outFIFO/N135 ), .B(n1467), .C(\u_outFIFO/N117 ), .D(
        \u_outFIFO/n514 ), .Q(\u_outFIFO/n513 ) );
  NOR21 U2999 ( .A(\u_coder/i [2]), .B(\u_coder/i [1]), .Q(\u_coder/n165 ) );
  NOR40 U3000 ( .A(n2287), .B(n1752), .C(\u_coder/j [1]), .D(\u_coder/j [19]), 
        .Q(n2288) );
  NAND22 U3001 ( .A(n2285), .B(n2284), .Q(n2287) );
  INV3 U3002 ( .A(n2286), .Q(n1752) );
  NOR21 U3003 ( .A(\u_coder/j [6]), .B(\u_coder/j [5]), .Q(n2285) );
  NAND22 U3004 ( .A(\u_coder/N974 ), .B(\u_coder/n144 ), .Q(\u_coder/n209 ) );
  NOR21 U3005 ( .A(\u_coder/j [2]), .B(\u_coder/j [1]), .Q(\u_coder/n208 ) );
  NAND22 U3006 ( .A(\u_outFIFO/currentState [2]), .B(\u_outFIFO/n173 ), .Q(
        \u_outFIFO/n538 ) );
  XNR21 U3007 ( .A(\u_coder/n140 ), .B(\u_coder/n175 ), .Q(\u_coder/n166 ) );
  OAI2111 U3008 ( .A(n1748), .B(n1712), .C(n1725), .D(\u_coder/n257 ), .Q(
        \u_coder/n344 ) );
  NAND31 U3009 ( .A(\u_coder/n254 ), .B(\u_coder/n186 ), .C(
        \sig_MUX_inMUX3[0] ), .Q(\u_coder/n257 ) );
  NAND22 U3010 ( .A(\u_inFIFO/n109 ), .B(\u_inFIFO/n76 ), .Q(\u_inFIFO/n200 )
         );
  NOR31 U3011 ( .A(\u_coder/j [7]), .B(\u_coder/j [9]), .C(\u_coder/j [8]), 
        .Q(n2284) );
  AOI221 U3012 ( .A(n1023), .B(n1111), .C(n1022), .D(n1014), .Q(n1015) );
  IMUX21 U3013 ( .A(n1022), .B(n1023), .S(n1109), .Q(n1024) );
  NOR40 U3014 ( .A(\u_cordic/my_rotation/n91 ), .B(n2225), .C(\u_cordic/dir ), 
        .D(n2224), .Q(\u_cordic/my_rotation/n90 ) );
  NAND22 U3015 ( .A(\u_cordic/my_rotation/n64 ), .B(\u_cordic/my_rotation/n63 ), .Q(\u_cordic/my_rotation/n91 ) );
  NAND22 U3016 ( .A(\u_outFIFO/outWriteCount[0] ), .B(n154), .Q(n2304) );
  NAND22 U3017 ( .A(\u_outFIFO/currentState [0]), .B(\u_outFIFO/n176 ), .Q(
        \u_outFIFO/n205 ) );
  NAND22 U3018 ( .A(\u_coder/n281 ), .B(\u_coder/i [3]), .Q(\u_coder/n261 ) );
  NOR21 U3019 ( .A(\u_inFIFO/n73 ), .B(\u_inFIFO/currentState [3]), .Q(
        \u_inFIFO/n109 ) );
  NAND22 U3020 ( .A(\u_coder/N974 ), .B(\u_coder/isPositiveQ ), .Q(
        \u_coder/n240 ) );
  NOR21 U3021 ( .A(n181), .B(\u_outFIFO/outWriteCount[2] ), .Q(n2314) );
  NAND22 U3022 ( .A(\u_decoder/fir_filter/I_data_mult_0_buff [1]), .B(n924), 
        .Q(\u_decoder/fir_filter/n1135 ) );
  NAND22 U3023 ( .A(\u_decoder/fir_filter/I_data_mult_1_buff [1]), .B(n920), 
        .Q(\u_decoder/fir_filter/n1119 ) );
  NAND22 U3024 ( .A(\u_decoder/fir_filter/I_data_mult_2_buff [2]), .B(n923), 
        .Q(\u_decoder/fir_filter/n1104 ) );
  NAND22 U3025 ( .A(\u_decoder/fir_filter/I_data_mult_6_buff [2]), .B(n920), 
        .Q(\u_decoder/fir_filter/n1039 ) );
  NAND22 U3026 ( .A(\u_decoder/fir_filter/I_data_mult_7_buff [1]), .B(n922), 
        .Q(\u_decoder/fir_filter/n1021 ) );
  NAND22 U3027 ( .A(\u_decoder/fir_filter/Q_data_mult_0_buff [1]), .B(n915), 
        .Q(\u_decoder/fir_filter/n838 ) );
  NAND22 U3028 ( .A(\u_decoder/fir_filter/Q_data_mult_1_buff [1]), .B(n915), 
        .Q(\u_decoder/fir_filter/n822 ) );
  NAND22 U3029 ( .A(\u_decoder/fir_filter/Q_data_mult_2_buff [2]), .B(n924), 
        .Q(\u_decoder/fir_filter/n807 ) );
  NAND22 U3030 ( .A(\u_decoder/fir_filter/Q_data_mult_6_buff [2]), .B(n917), 
        .Q(\u_decoder/fir_filter/n742 ) );
  NAND22 U3031 ( .A(\u_decoder/fir_filter/Q_data_mult_7_buff [1]), .B(n916), 
        .Q(\u_decoder/fir_filter/n724 ) );
  AOI221 U3032 ( .A(\u_outFIFO/N131 ), .B(n1467), .C(\u_outFIFO/n184 ), .D(
        \u_outFIFO/n514 ), .Q(\u_outFIFO/n518 ) );
  AOI221 U3033 ( .A(\u_outFIFO/N132 ), .B(n1467), .C(\u_outFIFO/N114 ), .D(
        \u_outFIFO/n514 ), .Q(\u_outFIFO/n517 ) );
  AOI221 U3034 ( .A(\u_outFIFO/N133 ), .B(n1467), .C(\u_outFIFO/N115 ), .D(
        \u_outFIFO/n514 ), .Q(\u_outFIFO/n516 ) );
  AOI221 U3035 ( .A(\u_outFIFO/N134 ), .B(n1467), .C(\u_outFIFO/N116 ), .D(
        \u_outFIFO/n514 ), .Q(\u_outFIFO/n515 ) );
  NAND22 U3036 ( .A(\u_decoder/fir_filter/I_data_mult_1_buff [5]), .B(n924), 
        .Q(\u_decoder/fir_filter/n1123 ) );
  NAND22 U3037 ( .A(\u_decoder/fir_filter/I_data_mult_7_buff [5]), .B(n919), 
        .Q(\u_decoder/fir_filter/n1025 ) );
  NAND22 U3038 ( .A(\u_decoder/fir_filter/Q_data_mult_1_buff [5]), .B(n915), 
        .Q(\u_decoder/fir_filter/n826 ) );
  NAND22 U3039 ( .A(\u_decoder/fir_filter/Q_data_mult_7_buff [5]), .B(n916), 
        .Q(\u_decoder/fir_filter/n728 ) );
  NAND22 U3040 ( .A(\u_decoder/fir_filter/I_data_mult_0_buff [4]), .B(n923), 
        .Q(\u_decoder/fir_filter/n1138 ) );
  NAND22 U3041 ( .A(\u_decoder/fir_filter/Q_data_mult_0_buff [4]), .B(n925), 
        .Q(\u_decoder/fir_filter/n841 ) );
  NAND22 U3042 ( .A(\u_decoder/fir_filter/I_data_mult_1_buff [6]), .B(n924), 
        .Q(\u_decoder/fir_filter/n1124 ) );
  NAND22 U3043 ( .A(\u_decoder/fir_filter/I_data_mult_7_buff [6]), .B(n919), 
        .Q(\u_decoder/fir_filter/n1026 ) );
  NAND22 U3044 ( .A(\u_decoder/fir_filter/Q_data_mult_1_buff [6]), .B(n915), 
        .Q(\u_decoder/fir_filter/n827 ) );
  NAND22 U3045 ( .A(\u_decoder/fir_filter/Q_data_mult_7_buff [6]), .B(n916), 
        .Q(\u_decoder/fir_filter/n729 ) );
  NAND22 U3046 ( .A(\u_decoder/fir_filter/I_data_mult_0_buff [5]), .B(n920), 
        .Q(\u_decoder/fir_filter/n1139 ) );
  NAND22 U3047 ( .A(\u_decoder/fir_filter/Q_data_mult_0_buff [5]), .B(n914), 
        .Q(\u_decoder/fir_filter/n842 ) );
  INV3 U3048 ( .A(\u_outFIFO/n499 ), .Q(n1458) );
  INV3 U3049 ( .A(\u_outFIFO/n494 ), .Q(n1456) );
  INV3 U3050 ( .A(\u_outFIFO/n490 ), .Q(n1454) );
  INV3 U3051 ( .A(\u_outFIFO/n486 ), .Q(n1452) );
  INV3 U3052 ( .A(\u_outFIFO/n482 ), .Q(n1450) );
  INV3 U3053 ( .A(\u_outFIFO/n478 ), .Q(n1448) );
  INV3 U3054 ( .A(\u_outFIFO/n474 ), .Q(n1446) );
  INV3 U3055 ( .A(\u_outFIFO/n470 ), .Q(n1444) );
  INV3 U3056 ( .A(\u_outFIFO/n466 ), .Q(n1442) );
  INV3 U3057 ( .A(\u_outFIFO/n462 ), .Q(n1440) );
  INV3 U3058 ( .A(\u_outFIFO/n458 ), .Q(n1438) );
  INV3 U3059 ( .A(\u_outFIFO/n454 ), .Q(n1436) );
  INV3 U3060 ( .A(\u_outFIFO/n450 ), .Q(n1434) );
  INV3 U3061 ( .A(\u_outFIFO/n446 ), .Q(n1432) );
  INV3 U3062 ( .A(\u_outFIFO/n440 ), .Q(n1430) );
  INV3 U3063 ( .A(\u_outFIFO/n434 ), .Q(n1428) );
  INV3 U3064 ( .A(\u_outFIFO/n430 ), .Q(n1426) );
  INV3 U3065 ( .A(\u_outFIFO/n425 ), .Q(n1424) );
  INV3 U3066 ( .A(\u_outFIFO/n421 ), .Q(n1422) );
  INV3 U3067 ( .A(\u_outFIFO/n234 ), .Q(n1338) );
  INV3 U3068 ( .A(\u_outFIFO/n223 ), .Q(n1334) );
  XOR21 U3069 ( .A(\u_cordic/mycordic/add_262/carry [10]), .B(
        \u_cordic/mycordic/present_ANGLE_table[6][10] ), .Q(
        \u_cordic/mycordic/N625 ) );
  XOR21 U3070 ( .A(\u_cordic/mycordic/add_262/carry [9]), .B(
        \u_cordic/mycordic/present_ANGLE_table[6][9] ), .Q(
        \u_cordic/mycordic/N624 ) );
  AOI221 U3071 ( .A(\u_inFIFO/N135 ), .B(\u_inFIFO/n211 ), .C(\u_inFIFO/N128 ), 
        .D(\u_inFIFO/n212 ), .Q(\u_inFIFO/n222 ) );
  XOR21 U3072 ( .A(\u_inFIFO/add_263/carry [5]), .B(
        \u_inFIFO/outWriteCount[5] ), .Q(\u_inFIFO/N135 ) );
  AOI221 U3073 ( .A(\u_inFIFO/N134 ), .B(\u_inFIFO/n211 ), .C(\u_inFIFO/N127 ), 
        .D(\u_inFIFO/n212 ), .Q(\u_inFIFO/n215 ) );
  NAND22 U3074 ( .A(\u_decoder/fir_filter/I_data_mult_1_buff [2]), .B(n921), 
        .Q(\u_decoder/fir_filter/n1120 ) );
  NAND22 U3075 ( .A(\u_decoder/fir_filter/I_data_mult_7_buff [2]), .B(n916), 
        .Q(\u_decoder/fir_filter/n1022 ) );
  NAND22 U3076 ( .A(\u_decoder/fir_filter/Q_data_mult_1_buff [2]), .B(n915), 
        .Q(\u_decoder/fir_filter/n823 ) );
  NAND22 U3077 ( .A(\u_decoder/fir_filter/Q_data_mult_7_buff [2]), .B(n916), 
        .Q(\u_decoder/fir_filter/n725 ) );
  NAND22 U3078 ( .A(\u_decoder/fir_filter/I_data_mult_0_buff [0]), .B(n924), 
        .Q(\u_decoder/fir_filter/n1134 ) );
  NAND22 U3079 ( .A(\u_decoder/fir_filter/I_data_mult_1_buff [0]), .B(n923), 
        .Q(\u_decoder/fir_filter/n1118 ) );
  NAND22 U3080 ( .A(\u_decoder/fir_filter/I_data_mult_2_buff [1]), .B(n923), 
        .Q(\u_decoder/fir_filter/n1103 ) );
  NAND22 U3081 ( .A(\u_decoder/fir_filter/I_data_mult_3_buff [0]), .B(n922), 
        .Q(\u_decoder/fir_filter/n1086 ) );
  NAND22 U3082 ( .A(\u_decoder/fir_filter/I_data_mult_5_buff [0]), .B(n921), 
        .Q(\u_decoder/fir_filter/n1054 ) );
  NAND22 U3083 ( .A(\u_decoder/fir_filter/I_data_mult_6_buff [1]), .B(n920), 
        .Q(\u_decoder/fir_filter/n1038 ) );
  NAND22 U3084 ( .A(\u_decoder/fir_filter/I_data_mult_7_buff [0]), .B(n922), 
        .Q(\u_decoder/fir_filter/n1020 ) );
  NAND22 U3085 ( .A(\u_decoder/fir_filter/Q_data_mult_0_buff [0]), .B(n915), 
        .Q(\u_decoder/fir_filter/n837 ) );
  NAND22 U3086 ( .A(\u_decoder/fir_filter/Q_data_mult_1_buff [0]), .B(n913), 
        .Q(\u_decoder/fir_filter/n821 ) );
  NAND22 U3087 ( .A(\u_decoder/fir_filter/Q_data_mult_2_buff [1]), .B(n922), 
        .Q(\u_decoder/fir_filter/n806 ) );
  NAND22 U3088 ( .A(\u_decoder/fir_filter/Q_data_mult_3_buff [0]), .B(n916), 
        .Q(\u_decoder/fir_filter/n789 ) );
  NAND22 U3089 ( .A(\u_decoder/fir_filter/Q_data_mult_5_buff [0]), .B(n918), 
        .Q(\u_decoder/fir_filter/n757 ) );
  NAND22 U3090 ( .A(\u_decoder/fir_filter/Q_data_mult_6_buff [1]), .B(n919), 
        .Q(\u_decoder/fir_filter/n741 ) );
  NAND22 U3091 ( .A(\u_decoder/fir_filter/Q_data_mult_7_buff [0]), .B(n916), 
        .Q(\u_decoder/fir_filter/n723 ) );
  INV3 U3092 ( .A(\u_outFIFO/n501 ), .Q(n1459) );
  INV3 U3093 ( .A(\u_outFIFO/n492 ), .Q(n1455) );
  INV3 U3094 ( .A(\u_outFIFO/n484 ), .Q(n1451) );
  INV3 U3095 ( .A(\u_outFIFO/n476 ), .Q(n1447) );
  INV3 U3096 ( .A(\u_outFIFO/n468 ), .Q(n1443) );
  INV3 U3097 ( .A(\u_outFIFO/n460 ), .Q(n1439) );
  INV3 U3098 ( .A(\u_outFIFO/n452 ), .Q(n1435) );
  INV3 U3099 ( .A(\u_outFIFO/n443 ), .Q(n1431) );
  INV3 U3100 ( .A(\u_outFIFO/n432 ), .Q(n1427) );
  INV3 U3101 ( .A(\u_outFIFO/n423 ), .Q(n1423) );
  INV3 U3102 ( .A(\u_outFIFO/n417 ), .Q(n1420) );
  INV3 U3103 ( .A(\u_outFIFO/n415 ), .Q(n1419) );
  INV3 U3104 ( .A(\u_outFIFO/n413 ), .Q(n1418) );
  INV3 U3105 ( .A(\u_outFIFO/n409 ), .Q(n1416) );
  INV3 U3106 ( .A(\u_outFIFO/n407 ), .Q(n1415) );
  INV3 U3107 ( .A(\u_outFIFO/n405 ), .Q(n1414) );
  INV3 U3108 ( .A(\u_outFIFO/n401 ), .Q(n1412) );
  INV3 U3109 ( .A(\u_outFIFO/n399 ), .Q(n1411) );
  INV3 U3110 ( .A(\u_outFIFO/n397 ), .Q(n1410) );
  INV3 U3111 ( .A(\u_outFIFO/n393 ), .Q(n1408) );
  INV3 U3112 ( .A(\u_outFIFO/n391 ), .Q(n1407) );
  INV3 U3113 ( .A(\u_outFIFO/n389 ), .Q(n1406) );
  INV3 U3114 ( .A(\u_outFIFO/n385 ), .Q(n1404) );
  INV3 U3115 ( .A(\u_outFIFO/n383 ), .Q(n1403) );
  INV3 U3116 ( .A(\u_outFIFO/n381 ), .Q(n1402) );
  INV3 U3117 ( .A(\u_outFIFO/n377 ), .Q(n1400) );
  INV3 U3118 ( .A(\u_outFIFO/n374 ), .Q(n1399) );
  INV3 U3119 ( .A(\u_outFIFO/n371 ), .Q(n1398) );
  INV3 U3120 ( .A(\u_outFIFO/n365 ), .Q(n1396) );
  INV3 U3121 ( .A(\u_outFIFO/n363 ), .Q(n1395) );
  INV3 U3122 ( .A(\u_outFIFO/n361 ), .Q(n1394) );
  INV3 U3123 ( .A(\u_outFIFO/n356 ), .Q(n1392) );
  INV3 U3124 ( .A(\u_outFIFO/n354 ), .Q(n1391) );
  INV3 U3125 ( .A(\u_outFIFO/n352 ), .Q(n1390) );
  INV3 U3126 ( .A(\u_outFIFO/n348 ), .Q(n1388) );
  INV3 U3127 ( .A(\u_outFIFO/n346 ), .Q(n1387) );
  INV3 U3128 ( .A(\u_outFIFO/n344 ), .Q(n1386) );
  INV3 U3129 ( .A(\u_outFIFO/n340 ), .Q(n1384) );
  INV3 U3130 ( .A(\u_outFIFO/n338 ), .Q(n1383) );
  INV3 U3131 ( .A(\u_outFIFO/n336 ), .Q(n1382) );
  INV3 U3132 ( .A(\u_outFIFO/n332 ), .Q(n1380) );
  INV3 U3133 ( .A(\u_outFIFO/n330 ), .Q(n1379) );
  INV3 U3134 ( .A(\u_outFIFO/n328 ), .Q(n1378) );
  INV3 U3135 ( .A(\u_outFIFO/n324 ), .Q(n1376) );
  INV3 U3136 ( .A(\u_outFIFO/n322 ), .Q(n1375) );
  INV3 U3137 ( .A(\u_outFIFO/n320 ), .Q(n1374) );
  INV3 U3138 ( .A(\u_outFIFO/n316 ), .Q(n1372) );
  INV3 U3139 ( .A(\u_outFIFO/n314 ), .Q(n1371) );
  INV3 U3140 ( .A(\u_outFIFO/n312 ), .Q(n1370) );
  INV3 U3141 ( .A(\u_outFIFO/n308 ), .Q(n1368) );
  INV3 U3142 ( .A(\u_outFIFO/n305 ), .Q(n1367) );
  INV3 U3143 ( .A(\u_outFIFO/n302 ), .Q(n1366) );
  INV3 U3144 ( .A(\u_outFIFO/n296 ), .Q(n1364) );
  INV3 U3145 ( .A(\u_outFIFO/n290 ), .Q(n1362) );
  INV3 U3146 ( .A(\u_outFIFO/n283 ), .Q(n1360) );
  INV3 U3147 ( .A(\u_outFIFO/n279 ), .Q(n1358) );
  INV3 U3148 ( .A(\u_outFIFO/n274 ), .Q(n1356) );
  INV3 U3149 ( .A(\u_outFIFO/n265 ), .Q(n1352) );
  INV3 U3150 ( .A(\u_outFIFO/n256 ), .Q(n1348) );
  INV3 U3151 ( .A(\u_outFIFO/n247 ), .Q(n1344) );
  INV3 U3152 ( .A(\u_cordic/mycordic/n512 ), .Q(n1202) );
  AOI221 U3153 ( .A(\u_cordic/mycordic/N339 ), .B(n833), .C(
        \u_cordic/mycordic/N371 ), .D(n1578), .Q(\u_cordic/mycordic/n512 ) );
  XNR21 U3154 ( .A(\u_cordic/mycordic/present_ANGLE_table[1][7] ), .B(
        \u_cordic/mycordic/sub_196/carry[7] ), .Q(\u_cordic/mycordic/N371 ) );
  XOR21 U3155 ( .A(\u_cordic/mycordic/present_ANGLE_table[1][7] ), .B(
        \u_cordic/mycordic/add_191/carry[7] ), .Q(\u_cordic/mycordic/N339 ) );
  INV3 U3156 ( .A(\u_outFIFO/n243 ), .Q(n1342) );
  INV3 U3157 ( .A(\u_outFIFO/n238 ), .Q(n1340) );
  INV3 U3158 ( .A(\u_outFIFO/n232 ), .Q(n1337) );
  INV3 U3159 ( .A(\u_outFIFO/n229 ), .Q(n1336) );
  INV3 U3160 ( .A(\u_outFIFO/n226 ), .Q(n1335) );
  INV3 U3161 ( .A(\u_outFIFO/n220 ), .Q(n1333) );
  INV3 U3162 ( .A(\u_outFIFO/n216 ), .Q(n1332) );
  NAND22 U3163 ( .A(\u_decoder/fir_filter/I_data_mult_8_buff [14]), .B(n919), 
        .Q(\u_decoder/fir_filter/n1011 ) );
  NAND22 U3164 ( .A(\u_decoder/fir_filter/I_data_mult_8_buff [13]), .B(n918), 
        .Q(\u_decoder/fir_filter/n1010 ) );
  NAND22 U3165 ( .A(\u_decoder/fir_filter/I_data_mult_8_buff [12]), .B(n917), 
        .Q(\u_decoder/fir_filter/n1009 ) );
  NAND22 U3166 ( .A(\u_decoder/fir_filter/Q_data_mult_8_buff [14]), .B(n914), 
        .Q(\u_decoder/fir_filter/n713 ) );
  NAND22 U3167 ( .A(\u_decoder/fir_filter/Q_data_mult_8_buff [13]), .B(n914), 
        .Q(\u_decoder/fir_filter/n712 ) );
  NAND22 U3168 ( .A(\u_decoder/fir_filter/Q_data_mult_8_buff [12]), .B(n914), 
        .Q(\u_decoder/fir_filter/n711 ) );
  NAND22 U3169 ( .A(\u_decoder/fir_filter/I_data_mult_1_buff [3]), .B(n922), 
        .Q(\u_decoder/fir_filter/n1121 ) );
  NAND22 U3170 ( .A(\u_decoder/fir_filter/I_data_mult_2_buff [3]), .B(n923), 
        .Q(\u_decoder/fir_filter/n1105 ) );
  NAND22 U3171 ( .A(\u_decoder/fir_filter/I_data_mult_3_buff [1]), .B(n922), 
        .Q(\u_decoder/fir_filter/n1087 ) );
  NAND22 U3172 ( .A(\u_decoder/fir_filter/I_data_mult_5_buff [1]), .B(n921), 
        .Q(\u_decoder/fir_filter/n1055 ) );
  NAND22 U3173 ( .A(\u_decoder/fir_filter/I_data_mult_6_buff [3]), .B(n920), 
        .Q(\u_decoder/fir_filter/n1040 ) );
  NAND22 U3174 ( .A(\u_decoder/fir_filter/I_data_mult_7_buff [3]), .B(n919), 
        .Q(\u_decoder/fir_filter/n1023 ) );
  NAND22 U3175 ( .A(\u_decoder/fir_filter/Q_data_mult_1_buff [3]), .B(n915), 
        .Q(\u_decoder/fir_filter/n824 ) );
  NAND22 U3176 ( .A(\u_decoder/fir_filter/Q_data_mult_2_buff [3]), .B(n923), 
        .Q(\u_decoder/fir_filter/n808 ) );
  NAND22 U3177 ( .A(\u_decoder/fir_filter/Q_data_mult_3_buff [1]), .B(n916), 
        .Q(\u_decoder/fir_filter/n790 ) );
  NAND22 U3178 ( .A(\u_decoder/fir_filter/Q_data_mult_5_buff [1]), .B(n918), 
        .Q(\u_decoder/fir_filter/n758 ) );
  NAND22 U3179 ( .A(\u_decoder/fir_filter/Q_data_mult_6_buff [3]), .B(n917), 
        .Q(\u_decoder/fir_filter/n743 ) );
  NAND22 U3180 ( .A(\u_decoder/fir_filter/Q_data_mult_7_buff [3]), .B(n916), 
        .Q(\u_decoder/fir_filter/n726 ) );
  NAND22 U3181 ( .A(\u_decoder/fir_filter/I_data_mult_0_buff [2]), .B(n924), 
        .Q(\u_decoder/fir_filter/n1136 ) );
  NAND22 U3182 ( .A(\u_decoder/fir_filter/Q_data_mult_0_buff [2]), .B(n927), 
        .Q(\u_decoder/fir_filter/n839 ) );
  NAND22 U3183 ( .A(\u_decoder/fir_filter/I_data_mult_8_buff [11]), .B(n916), 
        .Q(\u_decoder/fir_filter/n1008 ) );
  NAND22 U3184 ( .A(\u_decoder/fir_filter/I_data_mult_8_buff [10]), .B(n927), 
        .Q(\u_decoder/fir_filter/n1007 ) );
  NAND22 U3185 ( .A(\u_decoder/fir_filter/I_data_mult_8_buff [9]), .B(n926), 
        .Q(\u_decoder/fir_filter/n1006 ) );
  NAND22 U3186 ( .A(\u_decoder/fir_filter/I_data_mult_8_buff [8]), .B(n925), 
        .Q(\u_decoder/fir_filter/n1005 ) );
  NAND22 U3187 ( .A(\u_decoder/fir_filter/I_data_mult_8_buff [7]), .B(n915), 
        .Q(\u_decoder/fir_filter/n1004 ) );
  NAND22 U3188 ( .A(\u_decoder/fir_filter/I_data_mult_8_buff [6]), .B(n913), 
        .Q(\u_decoder/fir_filter/n1003 ) );
  NAND22 U3189 ( .A(\u_decoder/fir_filter/I_data_mult_8_buff [5]), .B(n913), 
        .Q(\u_decoder/fir_filter/n1002 ) );
  NAND22 U3190 ( .A(\u_decoder/fir_filter/I_data_mult_8_buff [4]), .B(n913), 
        .Q(\u_decoder/fir_filter/n1001 ) );
  NAND22 U3191 ( .A(\u_decoder/fir_filter/I_data_mult_8_buff [3]), .B(n913), 
        .Q(\u_decoder/fir_filter/n1000 ) );
  NAND22 U3192 ( .A(\u_decoder/fir_filter/I_data_mult_8_buff [2]), .B(n913), 
        .Q(\u_decoder/fir_filter/n999 ) );
  NAND22 U3193 ( .A(\u_decoder/fir_filter/I_data_mult_8_buff [1]), .B(n913), 
        .Q(\u_decoder/fir_filter/n998 ) );
  NAND22 U3194 ( .A(\u_decoder/fir_filter/I_data_mult_8_buff [0]), .B(n913), 
        .Q(\u_decoder/fir_filter/n997 ) );
  NAND22 U3195 ( .A(\u_decoder/fir_filter/Q_data_mult_8_buff [11]), .B(n914), 
        .Q(\u_decoder/fir_filter/n710 ) );
  NAND22 U3196 ( .A(\u_decoder/fir_filter/Q_data_mult_8_buff [10]), .B(n914), 
        .Q(\u_decoder/fir_filter/n709 ) );
  NAND22 U3197 ( .A(\u_decoder/fir_filter/Q_data_mult_8_buff [9]), .B(n914), 
        .Q(\u_decoder/fir_filter/n708 ) );
  NAND22 U3198 ( .A(\u_decoder/fir_filter/Q_data_mult_8_buff [8]), .B(n914), 
        .Q(\u_decoder/fir_filter/n707 ) );
  NAND22 U3199 ( .A(\u_decoder/fir_filter/Q_data_mult_8_buff [7]), .B(n914), 
        .Q(\u_decoder/fir_filter/n706 ) );
  NAND22 U3200 ( .A(\u_decoder/fir_filter/Q_data_mult_8_buff [6]), .B(n914), 
        .Q(\u_decoder/fir_filter/n705 ) );
  NAND22 U3201 ( .A(\u_decoder/fir_filter/Q_data_mult_8_buff [5]), .B(n914), 
        .Q(\u_decoder/fir_filter/n704 ) );
  NAND22 U3202 ( .A(\u_decoder/fir_filter/Q_data_mult_8_buff [4]), .B(n913), 
        .Q(\u_decoder/fir_filter/n703 ) );
  NAND22 U3203 ( .A(\u_decoder/fir_filter/Q_data_mult_8_buff [3]), .B(n913), 
        .Q(\u_decoder/fir_filter/n702 ) );
  NAND22 U3204 ( .A(\u_decoder/fir_filter/Q_data_mult_8_buff [2]), .B(n913), 
        .Q(\u_decoder/fir_filter/n701 ) );
  NAND22 U3205 ( .A(\u_decoder/fir_filter/Q_data_mult_8_buff [1]), .B(n913), 
        .Q(\u_decoder/fir_filter/n700 ) );
  NAND22 U3206 ( .A(\u_decoder/fir_filter/Q_data_mult_8_buff [0]), .B(n913), 
        .Q(\u_decoder/fir_filter/n699 ) );
  NAND22 U3207 ( .A(\u_decoder/fir_filter/I_data_mult_2_buff [4]), .B(n923), 
        .Q(\u_decoder/fir_filter/n1106 ) );
  NAND22 U3208 ( .A(\u_decoder/fir_filter/I_data_mult_6_buff [4]), .B(n920), 
        .Q(\u_decoder/fir_filter/n1041 ) );
  NAND22 U3209 ( .A(\u_decoder/fir_filter/Q_data_mult_2_buff [4]), .B(n913), 
        .Q(\u_decoder/fir_filter/n809 ) );
  NAND22 U3210 ( .A(\u_decoder/fir_filter/Q_data_mult_6_buff [4]), .B(n918), 
        .Q(\u_decoder/fir_filter/n744 ) );
  NAND22 U3211 ( .A(\u_decoder/fir_filter/I_data_mult_1_buff [4]), .B(n920), 
        .Q(\u_decoder/fir_filter/n1122 ) );
  NAND22 U3212 ( .A(\u_decoder/fir_filter/I_data_mult_3_buff [5]), .B(n922), 
        .Q(\u_decoder/fir_filter/n1091 ) );
  NAND22 U3213 ( .A(\u_decoder/fir_filter/I_data_mult_3_buff [4]), .B(n922), 
        .Q(\u_decoder/fir_filter/n1090 ) );
  NAND22 U3214 ( .A(\u_decoder/fir_filter/I_data_mult_5_buff [5]), .B(n921), 
        .Q(\u_decoder/fir_filter/n1059 ) );
  NAND22 U3215 ( .A(\u_decoder/fir_filter/I_data_mult_5_buff [4]), .B(n921), 
        .Q(\u_decoder/fir_filter/n1058 ) );
  NAND22 U3216 ( .A(\u_decoder/fir_filter/I_data_mult_7_buff [4]), .B(n919), 
        .Q(\u_decoder/fir_filter/n1024 ) );
  NAND22 U3217 ( .A(\u_decoder/fir_filter/Q_data_mult_1_buff [4]), .B(n915), 
        .Q(\u_decoder/fir_filter/n825 ) );
  NAND22 U3218 ( .A(\u_decoder/fir_filter/Q_data_mult_3_buff [5]), .B(n916), 
        .Q(\u_decoder/fir_filter/n794 ) );
  NAND22 U3219 ( .A(\u_decoder/fir_filter/Q_data_mult_3_buff [4]), .B(n916), 
        .Q(\u_decoder/fir_filter/n793 ) );
  NAND22 U3220 ( .A(\u_decoder/fir_filter/Q_data_mult_5_buff [5]), .B(n918), 
        .Q(\u_decoder/fir_filter/n762 ) );
  NAND22 U3221 ( .A(\u_decoder/fir_filter/Q_data_mult_5_buff [4]), .B(n918), 
        .Q(\u_decoder/fir_filter/n761 ) );
  NAND22 U3222 ( .A(\u_decoder/fir_filter/Q_data_mult_7_buff [4]), .B(n916), 
        .Q(\u_decoder/fir_filter/n727 ) );
  NAND22 U3223 ( .A(\u_decoder/fir_filter/I_data_mult_2_buff [6]), .B(n923), 
        .Q(\u_decoder/fir_filter/n1108 ) );
  NAND22 U3224 ( .A(\u_decoder/fir_filter/I_data_mult_2_buff [5]), .B(n923), 
        .Q(\u_decoder/fir_filter/n1107 ) );
  NAND22 U3225 ( .A(\u_decoder/fir_filter/I_data_mult_6_buff [6]), .B(n920), 
        .Q(\u_decoder/fir_filter/n1043 ) );
  NAND22 U3226 ( .A(\u_decoder/fir_filter/I_data_mult_6_buff [5]), .B(n920), 
        .Q(\u_decoder/fir_filter/n1042 ) );
  NAND22 U3227 ( .A(\u_decoder/fir_filter/Q_data_mult_2_buff [6]), .B(n913), 
        .Q(\u_decoder/fir_filter/n811 ) );
  NAND22 U3228 ( .A(\u_decoder/fir_filter/Q_data_mult_2_buff [5]), .B(n913), 
        .Q(\u_decoder/fir_filter/n810 ) );
  NAND22 U3229 ( .A(\u_decoder/fir_filter/Q_data_mult_6_buff [6]), .B(n917), 
        .Q(\u_decoder/fir_filter/n746 ) );
  NAND22 U3230 ( .A(\u_decoder/fir_filter/Q_data_mult_6_buff [5]), .B(n916), 
        .Q(\u_decoder/fir_filter/n745 ) );
  NAND22 U3231 ( .A(\u_decoder/fir_filter/I_data_mult_3_buff [3]), .B(n922), 
        .Q(\u_decoder/fir_filter/n1089 ) );
  NAND22 U3232 ( .A(\u_decoder/fir_filter/I_data_mult_3_buff [2]), .B(n922), 
        .Q(\u_decoder/fir_filter/n1088 ) );
  NAND22 U3233 ( .A(\u_decoder/fir_filter/I_data_mult_5_buff [3]), .B(n921), 
        .Q(\u_decoder/fir_filter/n1057 ) );
  NAND22 U3234 ( .A(\u_decoder/fir_filter/I_data_mult_5_buff [2]), .B(n921), 
        .Q(\u_decoder/fir_filter/n1056 ) );
  NAND22 U3235 ( .A(\u_decoder/fir_filter/Q_data_mult_3_buff [3]), .B(n916), 
        .Q(\u_decoder/fir_filter/n792 ) );
  NAND22 U3236 ( .A(\u_decoder/fir_filter/Q_data_mult_3_buff [2]), .B(n916), 
        .Q(\u_decoder/fir_filter/n791 ) );
  NAND22 U3237 ( .A(\u_decoder/fir_filter/Q_data_mult_5_buff [3]), .B(n918), 
        .Q(\u_decoder/fir_filter/n760 ) );
  NAND22 U3238 ( .A(\u_decoder/fir_filter/Q_data_mult_5_buff [2]), .B(n918), 
        .Q(\u_decoder/fir_filter/n759 ) );
  NAND22 U3239 ( .A(\u_decoder/fir_filter/I_data_mult_0_buff [3]), .B(n919), 
        .Q(\u_decoder/fir_filter/n1137 ) );
  NAND22 U3240 ( .A(\u_decoder/fir_filter/Q_data_mult_0_buff [3]), .B(n914), 
        .Q(\u_decoder/fir_filter/n840 ) );
  INV3 U3241 ( .A(\u_cordic/mycordic/n406 ), .Q(n1549) );
  NAND22 U3242 ( .A(\u_cordic/mycordic/next_ANGLE_table[6][8] ), .B(n972), .Q(
        \u_cordic/mycordic/n406 ) );
  XNR21 U3243 ( .A(\u_cordic/mycordic/add_262/carry [8]), .B(
        \u_cordic/mycordic/present_ANGLE_table[6][8] ), .Q(
        \u_cordic/mycordic/N623 ) );
  INV3 U3244 ( .A(n2309), .Q(n1792) );
  AOI311 U3245 ( .A(n2312), .B(n2313), .C(n2307), .D(
        \u_outFIFO/outWriteCount[5] ), .Q(n2308) );
  OAI2111 U3246 ( .A(\u_outFIFO/outReadCount[3] ), .B(\u_outFIFO/n181 ), .C(
        n1794), .D(n2306), .Q(n2307) );
  INV3 U3247 ( .A(\u_cordic/my_rotation/n93 ), .Q(n2225) );
  AOI221 U3248 ( .A(\u_cordic/my_rotation/present_delta [8]), .B(n33), .C(
        \u_cordic/my_rotation/N49 ), .D(n748), .Q(\u_cordic/my_rotation/n93 )
         );
  XNR21 U3249 ( .A(\u_cordic/my_rotation/present_delta [8]), .B(
        \u_cordic/my_rotation/add_43/carry [8]), .Q(\u_cordic/my_rotation/N49 ) );
  INV3 U3250 ( .A(\u_outFIFO/n293 ), .Q(n1363) );
  INV3 U3251 ( .A(\u_outFIFO/n287 ), .Q(n1361) );
  INV3 U3252 ( .A(\u_outFIFO/n281 ), .Q(n1359) );
  INV3 U3253 ( .A(\u_outFIFO/n277 ), .Q(n1357) );
  INV3 U3254 ( .A(\u_outFIFO/n272 ), .Q(n1355) );
  INV3 U3255 ( .A(\u_outFIFO/n270 ), .Q(n1354) );
  INV3 U3256 ( .A(\u_outFIFO/n268 ), .Q(n1353) );
  INV3 U3257 ( .A(\u_outFIFO/n263 ), .Q(n1351) );
  INV3 U3258 ( .A(\u_outFIFO/n261 ), .Q(n1350) );
  INV3 U3259 ( .A(\u_outFIFO/n259 ), .Q(n1349) );
  INV3 U3260 ( .A(\u_outFIFO/n254 ), .Q(n1347) );
  INV3 U3261 ( .A(\u_outFIFO/n252 ), .Q(n1346) );
  INV3 U3262 ( .A(\u_outFIFO/n250 ), .Q(n1345) );
  INV3 U3263 ( .A(\u_outFIFO/n245 ), .Q(n1343) );
  INV3 U3264 ( .A(\u_outFIFO/n241 ), .Q(n1341) );
  INV3 U3265 ( .A(\u_outFIFO/n236 ), .Q(n1339) );
  INV3 U3266 ( .A(\u_outFIFO/n497 ), .Q(n1457) );
  INV3 U3267 ( .A(\u_outFIFO/n488 ), .Q(n1453) );
  INV3 U3268 ( .A(\u_outFIFO/n480 ), .Q(n1449) );
  INV3 U3269 ( .A(\u_outFIFO/n472 ), .Q(n1445) );
  INV3 U3270 ( .A(\u_outFIFO/n464 ), .Q(n1441) );
  INV3 U3271 ( .A(\u_outFIFO/n456 ), .Q(n1437) );
  INV3 U3272 ( .A(\u_outFIFO/n448 ), .Q(n1433) );
  INV3 U3273 ( .A(\u_outFIFO/n437 ), .Q(n1429) );
  INV3 U3274 ( .A(\u_outFIFO/n428 ), .Q(n1425) );
  INV3 U3275 ( .A(\u_outFIFO/n419 ), .Q(n1421) );
  INV3 U3276 ( .A(\u_outFIFO/n411 ), .Q(n1417) );
  INV3 U3277 ( .A(\u_outFIFO/n403 ), .Q(n1413) );
  INV3 U3278 ( .A(\u_outFIFO/n395 ), .Q(n1409) );
  INV3 U3279 ( .A(\u_outFIFO/n387 ), .Q(n1405) );
  INV3 U3280 ( .A(\u_outFIFO/n379 ), .Q(n1401) );
  INV3 U3281 ( .A(\u_outFIFO/n368 ), .Q(n1397) );
  INV3 U3282 ( .A(\u_outFIFO/n359 ), .Q(n1393) );
  INV3 U3283 ( .A(\u_outFIFO/n350 ), .Q(n1389) );
  INV3 U3284 ( .A(\u_outFIFO/n342 ), .Q(n1385) );
  INV3 U3285 ( .A(\u_outFIFO/n334 ), .Q(n1381) );
  INV3 U3286 ( .A(\u_outFIFO/n326 ), .Q(n1377) );
  INV3 U3287 ( .A(\u_outFIFO/n318 ), .Q(n1373) );
  INV3 U3288 ( .A(\u_outFIFO/n310 ), .Q(n1369) );
  INV3 U3289 ( .A(\u_outFIFO/n299 ), .Q(n1365) );
  XNR21 U3290 ( .A(n375), .B(n2687), .Q(\u_coder/n175 ) );
  NOR40 U3291 ( .A(\u_coder/i [16]), .B(n1723), .C(\u_coder/i [15]), .D(
        \u_coder/i [14]), .Q(n2298) );
  INV3 U3292 ( .A(n2292), .Q(n1723) );
  NOR21 U3293 ( .A(\u_coder/i [18]), .B(\u_coder/i [17]), .Q(n2292) );
  INV3 U3294 ( .A(n2283), .Q(n1755) );
  NOR21 U3295 ( .A(\u_coder/j [18]), .B(\u_coder/j [17]), .Q(n2283) );
  INV3 U3296 ( .A(n2305), .Q(n1794) );
  AOI2111 U3297 ( .A(n2304), .B(\u_outFIFO/outReadCount[1] ), .C(n1795), .D(
        n2314), .Q(n2305) );
  INV3 U3298 ( .A(n2303), .Q(n1795) );
  XNR21 U3299 ( .A(\u_cordic/mycordic/r173/carry [7]), .B(n377), .Q(n376) );
  INV3 U3300 ( .A(\u_cordic/mycordic/n344 ), .Q(n1237) );
  AOI221 U3301 ( .A(n1579), .B(\u_cordic/mycordic/N259 ), .C(n787), .D(
        \u_cordic/mycordic/N267 ), .Q(\u_cordic/mycordic/n344 ) );
  INV3 U3302 ( .A(\u_cordic/mycordic/n383 ), .Q(n1232) );
  AOI221 U3303 ( .A(n1579), .B(\u_cordic/mycordic/N291 ), .C(n787), .D(
        \u_cordic/mycordic/N259 ), .Q(\u_cordic/mycordic/n383 ) );
  INV3 U3304 ( .A(\u_decoder/fir_filter/n1071 ), .Q(n1861) );
  AOI221 U3305 ( .A(\u_decoder/I_prefilter [1]), .B(n845), .C(
        \u_decoder/fir_filter/I_data_mult_4_buff [1]), .D(n930), .Q(
        \u_decoder/fir_filter/n1071 ) );
  XNR21 U3306 ( .A(\u_cordic/mycordic/r173/carry [9]), .B(
        \u_cordic/mycordic/present_ANGLE_table[6][9] ), .Q(n378) );
  XNR21 U3307 ( .A(\u_cordic/mycordic/r173/carry [8]), .B(
        \u_cordic/mycordic/present_ANGLE_table[6][8] ), .Q(n379) );
  INV3 U3308 ( .A(\u_inFIFO/n199 ), .Q(n1615) );
  AOI221 U3309 ( .A(\u_inFIFO/n101 ), .B(\u_inFIFO/n195 ), .C(n968), .D(
        \u_inFIFO/j_FIFO [0]), .Q(\u_inFIFO/n199 ) );
  INV3 U3310 ( .A(\u_inFIFO/n198 ), .Q(n1616) );
  AOI221 U3311 ( .A(\u_inFIFO/N192 ), .B(\u_inFIFO/n195 ), .C(n968), .D(
        \u_inFIFO/j_FIFO [1]), .Q(\u_inFIFO/n198 ) );
  INV3 U3312 ( .A(\u_inFIFO/n197 ), .Q(n1617) );
  AOI221 U3313 ( .A(\u_inFIFO/N193 ), .B(\u_inFIFO/n195 ), .C(n968), .D(
        \u_inFIFO/j_FIFO [2]), .Q(\u_inFIFO/n197 ) );
  INV3 U3314 ( .A(\u_inFIFO/n196 ), .Q(n1618) );
  AOI221 U3315 ( .A(\u_inFIFO/N194 ), .B(\u_inFIFO/n195 ), .C(n968), .D(
        \u_inFIFO/j_FIFO [3]), .Q(\u_inFIFO/n196 ) );
  INV3 U3316 ( .A(\u_inFIFO/n194 ), .Q(n1619) );
  AOI221 U3317 ( .A(\u_inFIFO/N195 ), .B(\u_inFIFO/n195 ), .C(n968), .D(
        \u_inFIFO/j_FIFO [4]), .Q(\u_inFIFO/n194 ) );
  XOR21 U3318 ( .A(\u_inFIFO/add_357/carry [4]), .B(\u_inFIFO/j_FIFO [4]), .Q(
        \u_inFIFO/N195 ) );
  INV3 U3319 ( .A(\u_decoder/fir_filter/n1070 ), .Q(n1818) );
  AOI221 U3320 ( .A(n773), .B(n845), .C(
        \u_decoder/fir_filter/I_data_mult_4_buff [0]), .D(n930), .Q(
        \u_decoder/fir_filter/n1070 ) );
  INV3 U3321 ( .A(\u_cordic/mycordic/n495 ), .Q(n1296) );
  AOI221 U3322 ( .A(\u_cordic/mycordic/N404 ), .B(n832), .C(
        \u_cordic/mycordic/N436 ), .D(n1582), .Q(\u_cordic/mycordic/n495 ) );
  XNR21 U3323 ( .A(\u_cordic/mycordic/present_ANGLE_table[2][8] ), .B(
        \u_cordic/mycordic/sub_207/carry [8]), .Q(\u_cordic/mycordic/N436 ) );
  XOR21 U3324 ( .A(\u_cordic/mycordic/present_ANGLE_table[2][8] ), .B(
        \u_cordic/mycordic/add_202/carry [8]), .Q(\u_cordic/mycordic/N404 ) );
  INV3 U3325 ( .A(\u_cordic/mycordic/n494 ), .Q(n1297) );
  AOI221 U3326 ( .A(\u_cordic/mycordic/N405 ), .B(\u_cordic/mycordic/n332 ), 
        .C(\u_cordic/mycordic/N437 ), .D(n1582), .Q(\u_cordic/mycordic/n494 )
         );
  XOR21 U3327 ( .A(\u_cordic/mycordic/present_ANGLE_table[2][9] ), .B(
        \u_cordic/mycordic/add_202/carry [9]), .Q(\u_cordic/mycordic/N405 ) );
  XNR21 U3328 ( .A(\u_cordic/mycordic/present_ANGLE_table[2][9] ), .B(
        \u_cordic/mycordic/sub_207/carry [9]), .Q(\u_cordic/mycordic/N437 ) );
  INV3 U3329 ( .A(\u_cordic/mycordic/n511 ), .Q(n1203) );
  AOI221 U3330 ( .A(\u_cordic/mycordic/N340 ), .B(n833), .C(
        \u_cordic/mycordic/N372 ), .D(n1578), .Q(\u_cordic/mycordic/n511 ) );
  XNR21 U3331 ( .A(\u_cordic/mycordic/present_ANGLE_table[1][8] ), .B(
        \u_cordic/mycordic/sub_196/carry[8] ), .Q(\u_cordic/mycordic/N372 ) );
  XOR21 U3332 ( .A(\u_cordic/mycordic/present_ANGLE_table[1][8] ), .B(
        \u_cordic/mycordic/add_191/carry[8] ), .Q(\u_cordic/mycordic/N340 ) );
  INV3 U3333 ( .A(\u_decoder/fir_filter/n1072 ), .Q(n1863) );
  AOI221 U3334 ( .A(n770), .B(n845), .C(
        \u_decoder/fir_filter/I_data_mult_4_buff [2]), .D(n930), .Q(
        \u_decoder/fir_filter/n1072 ) );
  INV3 U3335 ( .A(\u_decoder/fir_filter/n1076 ), .Q(n1833) );
  AOI221 U3336 ( .A(\u_decoder/fir_filter/I_data_mult_4 [6]), .B(n845), .C(
        \u_decoder/fir_filter/I_data_mult_4_buff [6]), .D(n930), .Q(
        \u_decoder/fir_filter/n1076 ) );
  INV3 U3337 ( .A(\u_decoder/fir_filter/n1075 ), .Q(n1834) );
  AOI221 U3338 ( .A(\u_decoder/fir_filter/I_data_mult_4 [5]), .B(n845), .C(
        \u_decoder/fir_filter/I_data_mult_4_buff [5]), .D(n930), .Q(
        \u_decoder/fir_filter/n1075 ) );
  INV3 U3339 ( .A(\u_decoder/fir_filter/n1074 ), .Q(n1835) );
  AOI221 U3340 ( .A(\u_decoder/fir_filter/I_data_mult_4 [4]), .B(n845), .C(
        \u_decoder/fir_filter/I_data_mult_4_buff [4]), .D(n930), .Q(
        \u_decoder/fir_filter/n1074 ) );
  INV3 U3341 ( .A(\u_decoder/fir_filter/n1073 ), .Q(n1836) );
  AOI221 U3342 ( .A(\u_decoder/fir_filter/I_data_mult_4 [3]), .B(n845), .C(
        \u_decoder/fir_filter/I_data_mult_4_buff [3]), .D(n930), .Q(
        \u_decoder/fir_filter/n1073 ) );
  XOR21 U3343 ( .A(n768), .B(n773), .Q(\u_decoder/fir_filter/I_data_mult_4 [3]) );
  INV3 U3344 ( .A(\u_decoder/fir_filter/n996 ), .Q(n2199) );
  AOI221 U3345 ( .A(\u_decoder/fir_filter/I_data_add_7 [0]), .B(n845), .C(
        \u_decoder/fir_filter/I_data_add_7_buff [0]), .D(n930), .Q(
        \u_decoder/fir_filter/n996 ) );
  XOR21 U3346 ( .A(\u_decoder/fir_filter/I_data_mult_7_buff [0]), .B(
        \u_decoder/fir_filter/I_data_mult_8_buff [0]), .Q(
        \u_decoder/fir_filter/I_data_add_7 [0]) );
  INV3 U3347 ( .A(\u_decoder/fir_filter/n995 ), .Q(n2198) );
  AOI221 U3348 ( .A(\u_decoder/fir_filter/I_data_add_7 [1]), .B(n845), .C(
        \u_decoder/fir_filter/I_data_add_7_buff [1]), .D(n930), .Q(
        \u_decoder/fir_filter/n995 ) );
  INV3 U3349 ( .A(\u_decoder/fir_filter/n994 ), .Q(n2197) );
  AOI221 U3350 ( .A(\u_decoder/fir_filter/I_data_add_7 [2]), .B(n845), .C(
        \u_decoder/fir_filter/I_data_add_7_buff [2]), .D(n930), .Q(
        \u_decoder/fir_filter/n994 ) );
  INV3 U3351 ( .A(\u_decoder/fir_filter/n993 ), .Q(n2196) );
  AOI221 U3352 ( .A(\u_decoder/fir_filter/I_data_add_7 [3]), .B(n845), .C(
        \u_decoder/fir_filter/I_data_add_7_buff [3]), .D(n930), .Q(
        \u_decoder/fir_filter/n993 ) );
  INV3 U3353 ( .A(\u_decoder/fir_filter/n992 ), .Q(n2195) );
  AOI221 U3354 ( .A(\u_decoder/fir_filter/I_data_add_7 [4]), .B(n845), .C(
        \u_decoder/fir_filter/I_data_add_7_buff [4]), .D(n930), .Q(
        \u_decoder/fir_filter/n992 ) );
  INV3 U3355 ( .A(\u_decoder/fir_filter/n991 ), .Q(n2194) );
  AOI221 U3356 ( .A(\u_decoder/fir_filter/I_data_add_7 [5]), .B(n845), .C(
        \u_decoder/fir_filter/I_data_add_7_buff [5]), .D(n930), .Q(
        \u_decoder/fir_filter/n991 ) );
  INV3 U3357 ( .A(\u_decoder/fir_filter/n975 ), .Q(n2184) );
  AOI221 U3358 ( .A(\u_decoder/fir_filter/I_data_add_6 [0]), .B(n846), .C(
        \u_decoder/fir_filter/I_data_add_6_buff [0]), .D(n931), .Q(
        \u_decoder/fir_filter/n975 ) );
  XOR21 U3359 ( .A(\u_decoder/fir_filter/I_data_mult_6_buff [0]), .B(
        \u_decoder/fir_filter/I_data_add_7_buff [0]), .Q(
        \u_decoder/fir_filter/I_data_add_6 [0]) );
  INV3 U3360 ( .A(\u_decoder/fir_filter/n974 ), .Q(n2183) );
  AOI221 U3361 ( .A(\u_decoder/fir_filter/I_data_add_6 [1]), .B(n846), .C(
        \u_decoder/fir_filter/I_data_add_6_buff [1]), .D(n931), .Q(
        \u_decoder/fir_filter/n974 ) );
  INV3 U3362 ( .A(\u_decoder/fir_filter/n973 ), .Q(n2182) );
  AOI221 U3363 ( .A(\u_decoder/fir_filter/I_data_add_6 [2]), .B(n846), .C(
        \u_decoder/fir_filter/I_data_add_6_buff [2]), .D(n931), .Q(
        \u_decoder/fir_filter/n973 ) );
  INV3 U3364 ( .A(\u_decoder/fir_filter/n972 ), .Q(n2181) );
  AOI221 U3365 ( .A(\u_decoder/fir_filter/I_data_add_6 [3]), .B(n846), .C(
        \u_decoder/fir_filter/I_data_add_6_buff [3]), .D(n931), .Q(
        \u_decoder/fir_filter/n972 ) );
  INV3 U3366 ( .A(\u_decoder/fir_filter/n971 ), .Q(n2180) );
  AOI221 U3367 ( .A(\u_decoder/fir_filter/I_data_add_6 [4]), .B(n846), .C(
        \u_decoder/fir_filter/I_data_add_6_buff [4]), .D(n931), .Q(
        \u_decoder/fir_filter/n971 ) );
  INV3 U3368 ( .A(\u_decoder/fir_filter/n970 ), .Q(n2179) );
  AOI221 U3369 ( .A(\u_decoder/fir_filter/I_data_add_6 [5]), .B(n846), .C(
        \u_decoder/fir_filter/I_data_add_6_buff [5]), .D(n931), .Q(
        \u_decoder/fir_filter/n970 ) );
  INV3 U3370 ( .A(\u_decoder/fir_filter/n954 ), .Q(n2169) );
  AOI221 U3371 ( .A(\u_decoder/fir_filter/I_data_add_5 [0]), .B(n847), .C(
        \u_decoder/fir_filter/I_data_add_5_buff [0]), .D(n928), .Q(
        \u_decoder/fir_filter/n954 ) );
  XOR21 U3372 ( .A(\u_decoder/fir_filter/I_data_mult_5_buff [0]), .B(
        \u_decoder/fir_filter/I_data_add_6_buff [0]), .Q(
        \u_decoder/fir_filter/I_data_add_5 [0]) );
  INV3 U3373 ( .A(\u_decoder/fir_filter/n953 ), .Q(n2168) );
  AOI221 U3374 ( .A(\u_decoder/fir_filter/I_data_add_5 [1]), .B(n847), .C(
        \u_decoder/fir_filter/I_data_add_5_buff [1]), .D(n929), .Q(
        \u_decoder/fir_filter/n953 ) );
  INV3 U3375 ( .A(\u_decoder/fir_filter/n952 ), .Q(n2167) );
  AOI221 U3376 ( .A(\u_decoder/fir_filter/I_data_add_5 [2]), .B(n847), .C(
        \u_decoder/fir_filter/I_data_add_5_buff [2]), .D(n926), .Q(
        \u_decoder/fir_filter/n952 ) );
  INV3 U3377 ( .A(\u_decoder/fir_filter/n951 ), .Q(n2166) );
  AOI221 U3378 ( .A(\u_decoder/fir_filter/I_data_add_5 [3]), .B(n847), .C(
        \u_decoder/fir_filter/I_data_add_5_buff [3]), .D(n925), .Q(
        \u_decoder/fir_filter/n951 ) );
  INV3 U3379 ( .A(\u_decoder/fir_filter/n950 ), .Q(n2165) );
  AOI221 U3380 ( .A(\u_decoder/fir_filter/I_data_add_5 [4]), .B(n847), .C(
        \u_decoder/fir_filter/I_data_add_5_buff [4]), .D(n930), .Q(
        \u_decoder/fir_filter/n950 ) );
  INV3 U3381 ( .A(\u_decoder/fir_filter/n949 ), .Q(n2164) );
  AOI221 U3382 ( .A(\u_decoder/fir_filter/I_data_add_5 [5]), .B(n847), .C(
        \u_decoder/fir_filter/I_data_add_5_buff [5]), .D(n931), .Q(
        \u_decoder/fir_filter/n949 ) );
  INV3 U3383 ( .A(\u_decoder/fir_filter/n933 ), .Q(n2154) );
  AOI221 U3384 ( .A(\u_decoder/fir_filter/I_data_add_4 [0]), .B(n848), .C(
        \u_decoder/fir_filter/I_data_add_4_buff [0]), .D(n920), .Q(
        \u_decoder/fir_filter/n933 ) );
  XOR21 U3385 ( .A(\u_decoder/fir_filter/I_data_mult_4_buff [0]), .B(
        \u_decoder/fir_filter/I_data_add_5_buff [0]), .Q(
        \u_decoder/fir_filter/I_data_add_4 [0]) );
  INV3 U3386 ( .A(\u_decoder/fir_filter/n932 ), .Q(n2153) );
  AOI221 U3387 ( .A(\u_decoder/fir_filter/I_data_add_4 [1]), .B(n848), .C(
        \u_decoder/fir_filter/I_data_add_4_buff [1]), .D(n921), .Q(
        \u_decoder/fir_filter/n932 ) );
  INV3 U3388 ( .A(\u_decoder/fir_filter/n931 ), .Q(n2152) );
  AOI221 U3389 ( .A(\u_decoder/fir_filter/I_data_add_4 [2]), .B(n848), .C(
        \u_decoder/fir_filter/I_data_add_4_buff [2]), .D(n932), .Q(
        \u_decoder/fir_filter/n931 ) );
  INV3 U3390 ( .A(\u_decoder/fir_filter/n930 ), .Q(n2151) );
  AOI221 U3391 ( .A(\u_decoder/fir_filter/I_data_add_4 [3]), .B(n848), .C(
        \u_decoder/fir_filter/I_data_add_4_buff [3]), .D(n932), .Q(
        \u_decoder/fir_filter/n930 ) );
  INV3 U3392 ( .A(\u_decoder/fir_filter/n929 ), .Q(n2150) );
  AOI221 U3393 ( .A(\u_decoder/fir_filter/I_data_add_4 [4]), .B(n848), .C(
        \u_decoder/fir_filter/I_data_add_4_buff [4]), .D(n932), .Q(
        \u_decoder/fir_filter/n929 ) );
  INV3 U3394 ( .A(\u_decoder/fir_filter/n928 ), .Q(n2149) );
  AOI221 U3395 ( .A(\u_decoder/fir_filter/I_data_add_4 [5]), .B(n848), .C(
        \u_decoder/fir_filter/I_data_add_4_buff [5]), .D(n932), .Q(
        \u_decoder/fir_filter/n928 ) );
  INV3 U3396 ( .A(\u_decoder/fir_filter/n912 ), .Q(n2139) );
  AOI221 U3397 ( .A(\u_decoder/fir_filter/I_data_add_3 [0]), .B(n849), .C(
        \u_decoder/fir_filter/I_data_add_3_buff [0]), .D(n932), .Q(
        \u_decoder/fir_filter/n912 ) );
  XOR21 U3398 ( .A(\u_decoder/fir_filter/I_data_mult_3_buff [0]), .B(
        \u_decoder/fir_filter/I_data_add_4_buff [0]), .Q(
        \u_decoder/fir_filter/I_data_add_3 [0]) );
  INV3 U3399 ( .A(\u_decoder/fir_filter/n911 ), .Q(n2138) );
  AOI221 U3400 ( .A(\u_decoder/fir_filter/I_data_add_3 [1]), .B(n849), .C(
        \u_decoder/fir_filter/I_data_add_3_buff [1]), .D(n932), .Q(
        \u_decoder/fir_filter/n911 ) );
  INV3 U3401 ( .A(\u_decoder/fir_filter/n910 ), .Q(n2137) );
  AOI221 U3402 ( .A(\u_decoder/fir_filter/I_data_add_3 [2]), .B(n849), .C(
        \u_decoder/fir_filter/I_data_add_3_buff [2]), .D(n932), .Q(
        \u_decoder/fir_filter/n910 ) );
  INV3 U3403 ( .A(\u_decoder/fir_filter/n909 ), .Q(n2136) );
  AOI221 U3404 ( .A(\u_decoder/fir_filter/I_data_add_3 [3]), .B(n849), .C(
        \u_decoder/fir_filter/I_data_add_3_buff [3]), .D(n932), .Q(
        \u_decoder/fir_filter/n909 ) );
  INV3 U3405 ( .A(\u_decoder/fir_filter/n908 ), .Q(n2135) );
  AOI221 U3406 ( .A(\u_decoder/fir_filter/I_data_add_3 [4]), .B(n849), .C(
        \u_decoder/fir_filter/I_data_add_3_buff [4]), .D(n930), .Q(
        \u_decoder/fir_filter/n908 ) );
  INV3 U3407 ( .A(\u_decoder/fir_filter/n907 ), .Q(n2134) );
  AOI221 U3408 ( .A(\u_decoder/fir_filter/I_data_add_3 [5]), .B(n849), .C(
        \u_decoder/fir_filter/I_data_add_3_buff [5]), .D(n931), .Q(
        \u_decoder/fir_filter/n907 ) );
  INV3 U3409 ( .A(\u_decoder/fir_filter/n635 ), .Q(n2034) );
  AOI221 U3410 ( .A(\u_decoder/fir_filter/Q_data_add_4 [0]), .B(n841), .C(
        \u_decoder/fir_filter/Q_data_add_4_buff [0]), .D(n927), .Q(
        \u_decoder/fir_filter/n635 ) );
  XOR21 U3411 ( .A(\u_decoder/fir_filter/Q_data_mult_4_buff [0]), .B(
        \u_decoder/fir_filter/Q_data_add_5_buff [0]), .Q(
        \u_decoder/fir_filter/Q_data_add_4 [0]) );
  INV3 U3412 ( .A(\u_decoder/fir_filter/n634 ), .Q(n2033) );
  AOI221 U3413 ( .A(\u_decoder/fir_filter/Q_data_add_4 [1]), .B(n841), .C(
        \u_decoder/fir_filter/Q_data_add_4_buff [1]), .D(n927), .Q(
        \u_decoder/fir_filter/n634 ) );
  INV3 U3414 ( .A(\u_decoder/fir_filter/n633 ), .Q(n2032) );
  AOI221 U3415 ( .A(\u_decoder/fir_filter/Q_data_add_4 [2]), .B(n841), .C(
        \u_decoder/fir_filter/Q_data_add_4_buff [2]), .D(n927), .Q(
        \u_decoder/fir_filter/n633 ) );
  INV3 U3416 ( .A(\u_decoder/fir_filter/n632 ), .Q(n2031) );
  AOI221 U3417 ( .A(\u_decoder/fir_filter/Q_data_add_4 [3]), .B(n841), .C(
        \u_decoder/fir_filter/Q_data_add_4_buff [3]), .D(n927), .Q(
        \u_decoder/fir_filter/n632 ) );
  INV3 U3418 ( .A(\u_decoder/fir_filter/n631 ), .Q(n2030) );
  AOI221 U3419 ( .A(\u_decoder/fir_filter/Q_data_add_4 [4]), .B(n841), .C(
        \u_decoder/fir_filter/Q_data_add_4_buff [4]), .D(n927), .Q(
        \u_decoder/fir_filter/n631 ) );
  INV3 U3420 ( .A(\u_decoder/fir_filter/n630 ), .Q(n2029) );
  AOI221 U3421 ( .A(\u_decoder/fir_filter/Q_data_add_4 [5]), .B(n841), .C(
        \u_decoder/fir_filter/Q_data_add_4_buff [5]), .D(n926), .Q(
        \u_decoder/fir_filter/n630 ) );
  INV3 U3422 ( .A(\u_decoder/fir_filter/n614 ), .Q(n2019) );
  AOI221 U3423 ( .A(\u_decoder/fir_filter/Q_data_add_3 [0]), .B(n841), .C(
        \u_decoder/fir_filter/Q_data_add_3_buff [0]), .D(n926), .Q(
        \u_decoder/fir_filter/n614 ) );
  XOR21 U3424 ( .A(\u_decoder/fir_filter/Q_data_mult_3_buff [0]), .B(
        \u_decoder/fir_filter/Q_data_add_4_buff [0]), .Q(
        \u_decoder/fir_filter/Q_data_add_3 [0]) );
  INV3 U3425 ( .A(\u_decoder/fir_filter/n613 ), .Q(n2018) );
  AOI221 U3426 ( .A(\u_decoder/fir_filter/Q_data_add_3 [1]), .B(n842), .C(
        \u_decoder/fir_filter/Q_data_add_3_buff [1]), .D(n926), .Q(
        \u_decoder/fir_filter/n613 ) );
  INV3 U3427 ( .A(\u_decoder/fir_filter/n612 ), .Q(n2017) );
  AOI221 U3428 ( .A(\u_decoder/fir_filter/Q_data_add_3 [2]), .B(n842), .C(
        \u_decoder/fir_filter/Q_data_add_3_buff [2]), .D(n926), .Q(
        \u_decoder/fir_filter/n612 ) );
  INV3 U3429 ( .A(\u_decoder/fir_filter/n611 ), .Q(n2016) );
  AOI221 U3430 ( .A(\u_decoder/fir_filter/Q_data_add_3 [3]), .B(n842), .C(
        \u_decoder/fir_filter/Q_data_add_3_buff [3]), .D(n926), .Q(
        \u_decoder/fir_filter/n611 ) );
  INV3 U3431 ( .A(\u_decoder/fir_filter/n610 ), .Q(n2015) );
  AOI221 U3432 ( .A(\u_decoder/fir_filter/Q_data_add_3 [4]), .B(n842), .C(
        \u_decoder/fir_filter/Q_data_add_3_buff [4]), .D(n926), .Q(
        \u_decoder/fir_filter/n610 ) );
  INV3 U3433 ( .A(\u_decoder/fir_filter/n609 ), .Q(n2014) );
  AOI221 U3434 ( .A(\u_decoder/fir_filter/Q_data_add_3 [5]), .B(n842), .C(
        \u_decoder/fir_filter/Q_data_add_3_buff [5]), .D(n926), .Q(
        \u_decoder/fir_filter/n609 ) );
  INV3 U3435 ( .A(\u_decoder/fir_filter/n593 ), .Q(n2004) );
  AOI221 U3436 ( .A(\u_decoder/fir_filter/Q_data_add_2 [0]), .B(n842), .C(
        \u_decoder/fir_filter/Q_data_add_2_buff [0]), .D(n925), .Q(
        \u_decoder/fir_filter/n593 ) );
  XOR21 U3437 ( .A(\u_decoder/fir_filter/Q_data_mult_2_buff [0]), .B(
        \u_decoder/fir_filter/Q_data_add_3_buff [0]), .Q(
        \u_decoder/fir_filter/Q_data_add_2 [0]) );
  INV3 U3438 ( .A(\u_decoder/fir_filter/n592 ), .Q(n2003) );
  AOI221 U3439 ( .A(\u_decoder/fir_filter/Q_data_add_2 [1]), .B(n842), .C(
        \u_decoder/fir_filter/Q_data_add_2_buff [1]), .D(n925), .Q(
        \u_decoder/fir_filter/n592 ) );
  INV3 U3440 ( .A(\u_decoder/fir_filter/n591 ), .Q(n2002) );
  AOI221 U3441 ( .A(\u_decoder/fir_filter/Q_data_add_2 [2]), .B(n842), .C(
        \u_decoder/fir_filter/Q_data_add_2_buff [2]), .D(n925), .Q(
        \u_decoder/fir_filter/n591 ) );
  INV3 U3442 ( .A(\u_decoder/fir_filter/n590 ), .Q(n2001) );
  AOI221 U3443 ( .A(\u_decoder/fir_filter/Q_data_add_2 [3]), .B(n843), .C(
        \u_decoder/fir_filter/Q_data_add_2_buff [3]), .D(n925), .Q(
        \u_decoder/fir_filter/n590 ) );
  INV3 U3444 ( .A(\u_decoder/fir_filter/n589 ), .Q(n2000) );
  AOI221 U3445 ( .A(\u_decoder/fir_filter/Q_data_add_2 [4]), .B(n843), .C(
        \u_decoder/fir_filter/Q_data_add_2_buff [4]), .D(n925), .Q(
        \u_decoder/fir_filter/n589 ) );
  INV3 U3446 ( .A(\u_decoder/fir_filter/n588 ), .Q(n1999) );
  AOI221 U3447 ( .A(\u_decoder/fir_filter/Q_data_add_2 [5]), .B(n843), .C(
        \u_decoder/fir_filter/Q_data_add_2_buff [5]), .D(n925), .Q(
        \u_decoder/fir_filter/n588 ) );
  INV3 U3448 ( .A(\u_decoder/fir_filter/n572 ), .Q(n1989) );
  AOI221 U3449 ( .A(\u_decoder/fir_filter/Q_data_add_1 [0]), .B(n843), .C(
        \u_decoder/fir_filter/Q_data_add_1_buff [0]), .D(n927), .Q(
        \u_decoder/fir_filter/n572 ) );
  XOR21 U3450 ( .A(\u_decoder/fir_filter/Q_data_mult_1_buff [0]), .B(
        \u_decoder/fir_filter/Q_data_add_2_buff [0]), .Q(
        \u_decoder/fir_filter/Q_data_add_1 [0]) );
  INV3 U3451 ( .A(\u_decoder/fir_filter/n571 ), .Q(n1988) );
  AOI221 U3452 ( .A(\u_decoder/fir_filter/Q_data_add_1 [1]), .B(n843), .C(
        \u_decoder/fir_filter/Q_data_add_1_buff [1]), .D(n926), .Q(
        \u_decoder/fir_filter/n571 ) );
  INV3 U3453 ( .A(\u_decoder/fir_filter/n570 ), .Q(n1986) );
  AOI221 U3454 ( .A(\u_decoder/fir_filter/Q_data_add_1 [2]), .B(n843), .C(
        \u_decoder/fir_filter/Q_data_add_1_buff [2]), .D(n925), .Q(
        \u_decoder/fir_filter/n570 ) );
  INV3 U3455 ( .A(\u_decoder/fir_filter/n569 ), .Q(n1984) );
  AOI221 U3456 ( .A(\u_decoder/fir_filter/Q_data_add_1 [3]), .B(n843), .C(
        \u_decoder/fir_filter/Q_data_add_1_buff [3]), .D(n924), .Q(
        \u_decoder/fir_filter/n569 ) );
  INV3 U3457 ( .A(\u_decoder/fir_filter/n568 ), .Q(n1982) );
  AOI221 U3458 ( .A(\u_decoder/fir_filter/Q_data_add_1 [4]), .B(n843), .C(
        \u_decoder/fir_filter/Q_data_add_1_buff [4]), .D(n929), .Q(
        \u_decoder/fir_filter/n568 ) );
  INV3 U3459 ( .A(\u_decoder/fir_filter/n567 ), .Q(n1980) );
  AOI221 U3460 ( .A(\u_decoder/fir_filter/Q_data_add_1 [5]), .B(n844), .C(
        \u_decoder/fir_filter/Q_data_add_1_buff [5]), .D(n930), .Q(
        \u_decoder/fir_filter/n567 ) );
  INV3 U3461 ( .A(\u_decoder/fir_filter/n891 ), .Q(n2124) );
  AOI221 U3462 ( .A(\u_decoder/fir_filter/I_data_add_2 [0]), .B(n850), .C(
        \u_decoder/fir_filter/I_data_add_2_buff [0]), .D(n928), .Q(
        \u_decoder/fir_filter/n891 ) );
  XOR21 U3463 ( .A(\u_decoder/fir_filter/I_data_mult_2_buff [0]), .B(
        \u_decoder/fir_filter/I_data_add_3_buff [0]), .Q(
        \u_decoder/fir_filter/I_data_add_2 [0]) );
  INV3 U3464 ( .A(\u_decoder/fir_filter/n890 ), .Q(n2123) );
  AOI221 U3465 ( .A(\u_decoder/fir_filter/I_data_add_2 [1]), .B(n850), .C(
        \u_decoder/fir_filter/I_data_add_2_buff [1]), .D(n928), .Q(
        \u_decoder/fir_filter/n890 ) );
  INV3 U3466 ( .A(\u_decoder/fir_filter/n889 ), .Q(n2122) );
  AOI221 U3467 ( .A(\u_decoder/fir_filter/I_data_add_2 [2]), .B(n850), .C(
        \u_decoder/fir_filter/I_data_add_2_buff [2]), .D(n929), .Q(
        \u_decoder/fir_filter/n889 ) );
  INV3 U3468 ( .A(\u_decoder/fir_filter/n888 ), .Q(n2121) );
  AOI221 U3469 ( .A(\u_decoder/fir_filter/I_data_add_2 [3]), .B(n850), .C(
        \u_decoder/fir_filter/I_data_add_2_buff [3]), .D(n919), .Q(
        \u_decoder/fir_filter/n888 ) );
  INV3 U3470 ( .A(\u_decoder/fir_filter/n887 ), .Q(n2120) );
  AOI221 U3471 ( .A(\u_decoder/fir_filter/I_data_add_2 [4]), .B(n850), .C(
        \u_decoder/fir_filter/I_data_add_2_buff [4]), .D(n918), .Q(
        \u_decoder/fir_filter/n887 ) );
  INV3 U3472 ( .A(\u_decoder/fir_filter/n886 ), .Q(n2119) );
  AOI221 U3473 ( .A(\u_decoder/fir_filter/I_data_add_2 [5]), .B(n850), .C(
        \u_decoder/fir_filter/I_data_add_2_buff [5]), .D(n917), .Q(
        \u_decoder/fir_filter/n886 ) );
  INV3 U3474 ( .A(\u_decoder/fir_filter/n870 ), .Q(n2109) );
  AOI221 U3475 ( .A(\u_decoder/fir_filter/I_data_add_1 [0]), .B(n850), .C(
        \u_decoder/fir_filter/I_data_add_1_buff [0]), .D(n929), .Q(
        \u_decoder/fir_filter/n870 ) );
  XOR21 U3476 ( .A(\u_decoder/fir_filter/I_data_mult_1_buff [0]), .B(
        \u_decoder/fir_filter/I_data_add_2_buff [0]), .Q(
        \u_decoder/fir_filter/I_data_add_1 [0]) );
  INV3 U3477 ( .A(\u_decoder/fir_filter/n869 ), .Q(n2108) );
  AOI221 U3478 ( .A(\u_decoder/fir_filter/I_data_add_1 [1]), .B(n851), .C(
        \u_decoder/fir_filter/I_data_add_1_buff [1]), .D(n928), .Q(
        \u_decoder/fir_filter/n869 ) );
  INV3 U3479 ( .A(\u_decoder/fir_filter/n868 ), .Q(n2106) );
  AOI221 U3480 ( .A(\u_decoder/fir_filter/I_data_add_1 [2]), .B(n851), .C(
        \u_decoder/fir_filter/I_data_add_1_buff [2]), .D(n929), .Q(
        \u_decoder/fir_filter/n868 ) );
  INV3 U3481 ( .A(\u_decoder/fir_filter/n867 ), .Q(n2104) );
  AOI221 U3482 ( .A(\u_decoder/fir_filter/I_data_add_1 [3]), .B(n851), .C(
        \u_decoder/fir_filter/I_data_add_1_buff [3]), .D(n931), .Q(
        \u_decoder/fir_filter/n867 ) );
  INV3 U3483 ( .A(\u_decoder/fir_filter/n866 ), .Q(n2102) );
  AOI221 U3484 ( .A(\u_decoder/fir_filter/I_data_add_1 [4]), .B(n851), .C(
        \u_decoder/fir_filter/I_data_add_1_buff [4]), .D(n926), .Q(
        \u_decoder/fir_filter/n866 ) );
  INV3 U3485 ( .A(\u_decoder/fir_filter/n865 ), .Q(n2100) );
  AOI221 U3486 ( .A(\u_decoder/fir_filter/I_data_add_1 [5]), .B(n851), .C(
        \u_decoder/fir_filter/I_data_add_1_buff [5]), .D(n925), .Q(
        \u_decoder/fir_filter/n865 ) );
  INV3 U3487 ( .A(\u_cordic/mycordic/n480 ), .Q(n1270) );
  AOI221 U3488 ( .A(\u_cordic/mycordic/N463 ), .B(n836), .C(
        \u_cordic/mycordic/N491 ), .D(n1581), .Q(\u_cordic/mycordic/n480 ) );
  XNR21 U3489 ( .A(\u_cordic/mycordic/present_ANGLE_table[3][7] ), .B(
        \u_cordic/mycordic/sub_218/carry[7] ), .Q(\u_cordic/mycordic/N491 ) );
  XOR21 U3490 ( .A(\u_cordic/mycordic/present_ANGLE_table[3][7] ), .B(
        \u_cordic/mycordic/add_213/carry[7] ), .Q(\u_cordic/mycordic/N463 ) );
  INV3 U3491 ( .A(\u_cordic/mycordic/n479 ), .Q(n1271) );
  AOI221 U3492 ( .A(\u_cordic/mycordic/N464 ), .B(n836), .C(
        \u_cordic/mycordic/N492 ), .D(n1581), .Q(\u_cordic/mycordic/n479 ) );
  XOR21 U3493 ( .A(\u_cordic/mycordic/present_ANGLE_table[3][8] ), .B(
        \u_cordic/mycordic/add_213/carry[8] ), .Q(\u_cordic/mycordic/N464 ) );
  XNR21 U3494 ( .A(\u_cordic/mycordic/present_ANGLE_table[3][8] ), .B(
        \u_cordic/mycordic/sub_218/carry[8] ), .Q(\u_cordic/mycordic/N492 ) );
  INV3 U3495 ( .A(\u_cordic/mycordic/n464 ), .Q(n1246) );
  AOI221 U3496 ( .A(\u_cordic/mycordic/N508 ), .B(n788), .C(
        \u_cordic/mycordic/N525 ), .D(n1580), .Q(\u_cordic/mycordic/n464 ) );
  XOR21 U3497 ( .A(\u_cordic/mycordic/present_ANGLE_table[4][7] ), .B(
        \u_cordic/mycordic/add_224/carry[7] ), .Q(\u_cordic/mycordic/N508 ) );
  XNR21 U3498 ( .A(\u_cordic/mycordic/present_ANGLE_table[4][7] ), .B(
        \u_cordic/mycordic/sub_229/carry[7] ), .Q(\u_cordic/mycordic/N525 ) );
  INV3 U3499 ( .A(\u_cordic/mycordic/n463 ), .Q(n1247) );
  AOI221 U3500 ( .A(\u_cordic/mycordic/N509 ), .B(n789), .C(
        \u_cordic/mycordic/N526 ), .D(n1580), .Q(\u_cordic/mycordic/n463 ) );
  XOR21 U3501 ( .A(\u_cordic/mycordic/present_ANGLE_table[4][8] ), .B(
        \u_cordic/mycordic/add_224/carry[8] ), .Q(\u_cordic/mycordic/N509 ) );
  XNR21 U3502 ( .A(\u_cordic/mycordic/present_ANGLE_table[4][8] ), .B(
        \u_cordic/mycordic/sub_229/carry[8] ), .Q(\u_cordic/mycordic/N526 ) );
  INV3 U3503 ( .A(\u_cordic/mycordic/n445 ), .Q(n1187) );
  AOI221 U3504 ( .A(\u_cordic/mycordic/N542 ), .B(n786), .C(
        \u_cordic/mycordic/N558 ), .D(n1577), .Q(\u_cordic/mycordic/n445 ) );
  XOR21 U3505 ( .A(\u_cordic/mycordic/present_ANGLE_table[5][8] ), .B(
        \u_cordic/mycordic/add_233/carry [8]), .Q(\u_cordic/mycordic/N542 ) );
  XNR21 U3506 ( .A(\u_cordic/mycordic/present_ANGLE_table[5][8] ), .B(
        \u_cordic/mycordic/sub_236/carry [8]), .Q(\u_cordic/mycordic/N558 ) );
  INV3 U3507 ( .A(\u_cordic/mycordic/n444 ), .Q(n1188) );
  AOI221 U3508 ( .A(\u_cordic/mycordic/N543 ), .B(n786), .C(
        \u_cordic/mycordic/N559 ), .D(n1577), .Q(\u_cordic/mycordic/n444 ) );
  XOR21 U3509 ( .A(\u_cordic/mycordic/present_ANGLE_table[5][9] ), .B(
        \u_cordic/mycordic/add_233/carry [9]), .Q(\u_cordic/mycordic/N543 ) );
  XNR21 U3510 ( .A(\u_cordic/mycordic/present_ANGLE_table[5][9] ), .B(
        \u_cordic/mycordic/sub_236/carry [9]), .Q(\u_cordic/mycordic/N559 ) );
  INV3 U3511 ( .A(n2631), .Q(n1492) );
  NAND22 U3512 ( .A(\u_cdr/phd1/cnt_phd/N51 ), .B(n976), .Q(n2631) );
  NOR31 U3513 ( .A(n1080), .B(n1079), .C(n1078), .Q(\u_cdr/phd1/cnt_phd/N51 )
         );
  INV3 U3514 ( .A(\u_cordic/mycordic/n407 ), .Q(n1550) );
  NAND22 U3515 ( .A(\u_cordic/mycordic/next_ANGLE_table[6][7] ), .B(n972), .Q(
        \u_cordic/mycordic/n407 ) );
  INV3 U3516 ( .A(\u_cordic/mycordic/n405 ), .Q(n1548) );
  NAND22 U3517 ( .A(\u_cordic/mycordic/next_ANGLE_table[6][9] ), .B(n972), .Q(
        \u_cordic/mycordic/n405 ) );
  NOR31 U3518 ( .A(n1778), .B(\u_cordic/n18 ), .C(\u_cordic/n12 ), .Q(
        \u_cordic/n20 ) );
  NAND41 U3519 ( .A(\u_cdr/cnt_in [0]), .B(\u_cdr/cnt_in [2]), .C(n3), .D(n36), 
        .Q(\u_cdr/N100 ) );
  AOI211 U3520 ( .A(\u_outFIFO/currentState [1]), .B(\u_outFIFO/n206 ), .C(
        n982), .Q(\u_outFIFO/n209 ) );
  OAI311 U3521 ( .A(\u_inFIFO/n225 ), .B(\u_inFIFO/sigEnableCounter ), .C(
        n1702), .D(\u_inFIFO/n226 ), .Q(\u_inFIFO/n218 ) );
  XNR21 U3522 ( .A(\u_coder/n175 ), .B(\u_coder/sin_was_positiveQ ), .Q(
        \u_coder/n212 ) );
  NAND22 U3523 ( .A(\u_coder/my_clk_10M ), .B(\u_coder/stateI[0] ), .Q(
        \u_coder/n161 ) );
  NAND41 U3524 ( .A(n2281), .B(n2280), .C(n2279), .D(n2278), .Q(n2282) );
  NOR40 U3525 ( .A(\u_coder/i [4]), .B(\u_coder/i [19]), .C(\u_coder/i [18]), 
        .D(\u_coder/i [17]), .Q(n2279) );
  NOR40 U3526 ( .A(\u_coder/i [16]), .B(\u_coder/i [15]), .C(\u_coder/i [14]), 
        .D(\u_coder/i [13]), .Q(n2280) );
  NOR40 U3527 ( .A(\u_coder/i [7]), .B(n1722), .C(\u_coder/i [6]), .D(
        \u_coder/i [5]), .Q(n2278) );
  AOI221 U3528 ( .A(\sig_MUX_inMUX11[0] ), .B(n1692), .C(in_MUX_inSEL11), .D(
        sig_DEMUX_outDEMUX1[3]), .Q(n2689) );
  NOR31 U3529 ( .A(n1682), .B(in_DEMUX_inSEL1[2]), .C(\u_demux1/n4 ), .Q(
        sig_DEMUX_outDEMUX1[3]) );
  NAND41 U3530 ( .A(n2274), .B(n2273), .C(n2272), .D(n2271), .Q(n2275) );
  NOR40 U3531 ( .A(\u_coder/j [4]), .B(\u_coder/j [19]), .C(\u_coder/j [18]), 
        .D(\u_coder/j [17]), .Q(n2272) );
  NOR40 U3532 ( .A(\u_coder/j [16]), .B(\u_coder/j [15]), .C(\u_coder/j [14]), 
        .D(\u_coder/j [13]), .Q(n2273) );
  NOR40 U3533 ( .A(\u_coder/j [7]), .B(n1754), .C(\u_coder/j [6]), .D(
        \u_coder/j [5]), .Q(n2271) );
  OAI2111 U3534 ( .A(n777), .B(\u_coder/n134 ), .C(\u_coder/n222 ), .D(
        \u_coder/n223 ), .Q(\u_coder/n219 ) );
  AOI311 U3535 ( .A(n777), .B(\u_coder/n135 ), .C(\u_coder/j [1]), .D(
        \u_coder/n224 ), .Q(\u_coder/n223 ) );
  NOR31 U3536 ( .A(\u_coder/n138 ), .B(n776), .C(\u_coder/j [1]), .Q(
        \u_coder/n224 ) );
  OAI2111 U3537 ( .A(n778), .B(\u_coder/n85 ), .C(\u_coder/n179 ), .D(
        \u_coder/n180 ), .Q(\u_coder/n177 ) );
  AOI311 U3538 ( .A(n778), .B(\u_coder/n86 ), .C(\u_coder/i [1]), .D(
        \u_coder/n181 ), .Q(\u_coder/n180 ) );
  NOR31 U3539 ( .A(\u_coder/n89 ), .B(\u_coder/i [3]), .C(\u_coder/i [1]), .Q(
        \u_coder/n181 ) );
  NAND22 U3540 ( .A(\u_coder/stateQ[0] ), .B(\u_coder/my_clk_10M ), .Q(
        \u_coder/n200 ) );
  NOR31 U3541 ( .A(\u_coder/n262 ), .B(n1751), .C(\u_coder/n138 ), .Q(
        \u_coder/n280 ) );
  XNR21 U3542 ( .A(\u_coder/sin_was_positiveI ), .B(\u_coder/n175 ), .Q(
        \u_coder/n195 ) );
  NOR31 U3543 ( .A(\u_cordic/n12 ), .B(\u_cordic/present_state [0]), .C(
        \u_cordic/n11 ), .Q(\sig_MUX_inMUX11[0] ) );
  NAND22 U3544 ( .A(n978), .B(\u_coder/old_i_data ), .Q(\u_coder/n277 ) );
  INV3 U3545 ( .A(\u_coder/n276 ), .Q(n1713) );
  NOR21 U3546 ( .A(\u_coder/n141 ), .B(\u_coder/n145 ), .Q(\u_coder/n168 ) );
  AOI221 U3547 ( .A(\u_inFIFO/n86 ), .B(\u_inFIFO/n211 ), .C(\u_inFIFO/N123 ), 
        .D(\u_inFIFO/n212 ), .Q(\u_inFIFO/n216 ) );
  AOI221 U3548 ( .A(\u_inFIFO/N131 ), .B(\u_inFIFO/n211 ), .C(\u_inFIFO/N124 ), 
        .D(\u_inFIFO/n212 ), .Q(\u_inFIFO/n210 ) );
  AOI221 U3549 ( .A(\u_inFIFO/N132 ), .B(\u_inFIFO/n211 ), .C(\u_inFIFO/N125 ), 
        .D(\u_inFIFO/n212 ), .Q(\u_inFIFO/n213 ) );
  NOR40 U3550 ( .A(\u_coder/i [12]), .B(\u_coder/i [11]), .C(\u_coder/i [10]), 
        .D(n1717), .Q(n2281) );
  INV3 U3551 ( .A(n2276), .Q(n1717) );
  OAI311 U3552 ( .A(n778), .B(\u_coder/i [2]), .C(\u_coder/i [1]), .D(
        \u_coder/i [3]), .Q(n2276) );
  AOI2111 U3553 ( .A(n777), .B(n776), .C(\u_coder/n225 ), .D(\u_coder/j [1]), 
        .Q(\u_coder/n217 ) );
  NOR21 U3554 ( .A(\u_coder/n144 ), .B(\u_coder/n145 ), .Q(\u_coder/n218 ) );
  NOR21 U3555 ( .A(\u_coder/n145 ), .B(\u_coder/n168 ), .Q(\u_coder/n154 ) );
  AOI221 U3556 ( .A(\u_coder/isPositiveQ ), .B(n1726), .C(n1756), .D(n1655), 
        .Q(\u_coder/n248 ) );
  NOR40 U3557 ( .A(\u_coder/j [12]), .B(\u_coder/j [11]), .C(\u_coder/j [10]), 
        .D(n1747), .Q(n2274) );
  INV3 U3558 ( .A(n2269), .Q(n1747) );
  OAI311 U3559 ( .A(n777), .B(\u_coder/j [2]), .C(\u_coder/j [1]), .D(n776), 
        .Q(n2269) );
  XNR21 U3560 ( .A(\u_outFIFO/outWriteCount[0] ), .B(n154), .Q(
        \u_outFIFO/N131 ) );
  XNR21 U3561 ( .A(\u_cordic/n11 ), .B(\u_cordic/n13 ), .Q(\u_cordic/n29 ) );
  XNR21 U3562 ( .A(\u_inFIFO/outWriteCount[0] ), .B(n105), .Q(\u_inFIFO/N123 )
         );
  NAND22 U3563 ( .A(\u_cdr/cnt_in [0]), .B(\u_cdr/N100 ), .Q(
        \u_cdr/dp_cluster_0/mult_add_59_aco/PROD_not[0] ) );
  AOI221 U3564 ( .A(\u_cordic/my_rotation/present_delta [6]), .B(n33), .C(
        \u_cordic/my_rotation/N47 ), .D(n748), .Q(\u_cordic/my_rotation/n64 )
         );
  XNR21 U3565 ( .A(\u_cordic/my_rotation/present_delta [6]), .B(
        \u_cordic/my_rotation/add_43/carry [6]), .Q(\u_cordic/my_rotation/N47 ) );
  OAI2111 U3566 ( .A(\u_coder/n76 ), .B(n1712), .C(n1725), .D(\u_coder/n243 ), 
        .Q(\u_coder/n338 ) );
  NAND41 U3567 ( .A(n976), .B(\u_coder/is9 ), .C(\u_coder/stateQ[0] ), .D(
        \u_coder/stateI[0] ), .Q(\u_coder/n243 ) );
  NAND41 U3568 ( .A(\u_inFIFO/n86 ), .B(\u_inFIFO/n85 ), .C(
        \u_inFIFO/outWriteCount[5] ), .D(\u_inFIFO/n229 ), .Q(\u_inFIFO/n224 )
         );
  NOR31 U3569 ( .A(\u_inFIFO/outWriteCount[2] ), .B(
        \u_inFIFO/outWriteCount[4] ), .C(\u_inFIFO/outWriteCount[3] ), .Q(
        \u_inFIFO/n229 ) );
  NOR21 U3570 ( .A(\u_coder/n145 ), .B(\u_coder/n218 ), .Q(\u_coder/n220 ) );
  AOI211 U3571 ( .A(\u_cdr/cnt_d [1]), .B(n978), .C(\u_cdr/n26 ), .Q(
        \u_cdr/n41 ) );
  NOR21 U3572 ( .A(n983), .B(\u_outFIFO/sigEnableCounter ), .Q(
        \u_outFIFO/n530 ) );
  INV3 U3573 ( .A(\u_outFIFO/N122 ), .Q(n1797) );
  XNR21 U3574 ( .A(\u_outFIFO/add_256/carry [4]), .B(\u_outFIFO/i_FIFO [4]), 
        .Q(n380) );
  NAND31 U3575 ( .A(n1756), .B(\u_coder/n134 ), .C(\u_coder/n280 ), .Q(
        \u_coder/n279 ) );
  OAI311 U3576 ( .A(n3), .B(\u_cdr/cnt_in [0]), .C(\u_cdr/n29 ), .D(n978), .Q(
        \u_cdr/n27 ) );
  OAI311 U3577 ( .A(n294), .B(\u_cdr/cnt_in [1]), .C(\u_cdr/n29 ), .D(n978), 
        .Q(\u_cdr/n30 ) );
  OAI311 U3578 ( .A(n295), .B(\u_cdr/n22 ), .C(\u_cdr/n23 ), .D(\u_cdr/n24 ), 
        .Q(\u_cdr/n49 ) );
  MAJ31 U3579 ( .A(\u_cdr/n19 ), .B(\u_cdr/n18 ), .C(\u_cdr/n3 ), .Q(
        \u_cdr/n22 ) );
  NOR21 U3580 ( .A(\u_cdr/cnt_in [2]), .B(n982), .Q(\u_cdr/n25 ) );
  NAND22 U3581 ( .A(\u_outFIFO/outReadCount[4] ), .B(\u_outFIFO/n180 ), .Q(
        n2312) );
  AOI221 U3582 ( .A(\u_inFIFO/N133 ), .B(\u_inFIFO/n211 ), .C(\u_inFIFO/N126 ), 
        .D(\u_inFIFO/n212 ), .Q(\u_inFIFO/n214 ) );
  AOI2111 U3583 ( .A(\u_cdr/n38 ), .B(\u_cdr/n39 ), .C(n985), .D(\u_cdr/n40 ), 
        .Q(\u_cdr/n52 ) );
  NOR31 U3584 ( .A(\u_cdr/n16 ), .B(\u_cdr/cnt [1]), .C(\u_cdr/cnt [0]), .Q(
        \u_cdr/n40 ) );
  NAND22 U3585 ( .A(\u_cdr/flag ), .B(n2689), .Q(\u_cdr/n39 ) );
  NAND41 U3586 ( .A(n976), .B(\u_coder/IorQ ), .C(\u_coder/n309 ), .D(
        \u_coder/n310 ), .Q(\u_coder/n308 ) );
  NOR21 U3587 ( .A(n1714), .B(n1726), .Q(\u_coder/n307 ) );
  NAND22 U3588 ( .A(\u_outFIFO/outReadCount[3] ), .B(\u_outFIFO/n181 ), .Q(
        n2313) );
  INV3 U3589 ( .A(\u_cordic/mycordic/n514 ), .Q(n1200) );
  AOI221 U3590 ( .A(\u_cordic/mycordic/N337 ), .B(n833), .C(
        \u_cordic/mycordic/N369 ), .D(n1578), .Q(\u_cordic/mycordic/n514 ) );
  XNR21 U3591 ( .A(\u_cordic/mycordic/present_ANGLE_table[1][5] ), .B(
        \u_cordic/mycordic/sub_196/carry[5] ), .Q(\u_cordic/mycordic/N369 ) );
  XOR21 U3592 ( .A(\u_cordic/mycordic/present_ANGLE_table[1][5] ), .B(
        \u_cordic/mycordic/add_191/carry[5] ), .Q(\u_cordic/mycordic/N337 ) );
  INV3 U3593 ( .A(\u_cordic/mycordic/n513 ), .Q(n1201) );
  AOI221 U3594 ( .A(\u_cordic/mycordic/N338 ), .B(n833), .C(
        \u_cordic/mycordic/N370 ), .D(n1578), .Q(\u_cordic/mycordic/n513 ) );
  XNR21 U3595 ( .A(\u_cordic/mycordic/present_ANGLE_table[1][6] ), .B(
        \u_cordic/mycordic/sub_196/carry[6] ), .Q(\u_cordic/mycordic/N370 ) );
  XOR21 U3596 ( .A(\u_cordic/mycordic/present_ANGLE_table[1][6] ), .B(
        \u_cordic/mycordic/add_191/carry[6] ), .Q(\u_cordic/mycordic/N338 ) );
  BUF2 U3597 ( .A(\u_cordic/my_rotation/N39 ), .Q(n748) );
  BUF2 U3598 ( .A(\u_cordic/my_rotation/N39 ), .Q(n747) );
  XNR21 U3599 ( .A(\u_cordic/mycordic/add_262/carry [6]), .B(
        \u_cordic/mycordic/present_ANGLE_table[6][6] ), .Q(
        \u_cordic/mycordic/N621 ) );
  BUF2 U3600 ( .A(\u_outFIFO/n213 ), .Q(n805) );
  NAND31 U3601 ( .A(n978), .B(n958), .C(n1664), .Q(\u_outFIFO/n213 ) );
  INV3 U3602 ( .A(n2691), .Q(n1664) );
  AOI221 U3603 ( .A(\sig_MUX_inMUX13[0] ), .B(n1693), .C(in_MUX_inSEL12), .D(
        sig_DEMUX_outDEMUX2[4]), .Q(n2691) );
  NAND22 U3604 ( .A(\u_coder/n281 ), .B(\u_coder/n85 ), .Q(\u_coder/n278 ) );
  INV3 U3605 ( .A(\u_cdr/dp_cluster_0/mult_add_59_aco/PROD_not[1] ), .Q(n1786)
         );
  NAND22 U3606 ( .A(\u_cdr/cnt_in [1]), .B(\u_cdr/N100 ), .Q(
        \u_cdr/dp_cluster_0/mult_add_59_aco/PROD_not[1] ) );
  INV3 U3607 ( .A(\u_cordic/my_rotation/n95 ), .Q(n2227) );
  AOI221 U3608 ( .A(\u_cordic/my_rotation/present_delta [3]), .B(n33), .C(n266), .D(n748), .Q(\u_cordic/my_rotation/n95 ) );
  INV3 U3609 ( .A(\u_cordic/my_rotation/n97 ), .Q(n2229) );
  AOI221 U3610 ( .A(\u_cordic/my_rotation/present_delta [5]), .B(n33), .C(
        \u_cordic/my_rotation/N46 ), .D(n748), .Q(\u_cordic/my_rotation/n97 )
         );
  XNR21 U3611 ( .A(\u_cordic/my_rotation/present_delta [5]), .B(
        \u_cordic/my_rotation/add_43/carry [5]), .Q(\u_cordic/my_rotation/N46 ) );
  XOR21 U3612 ( .A(\u_cordic/mycordic/add_262/carry [7]), .B(
        \u_cordic/mycordic/present_ANGLE_table[6][7] ), .Q(
        \u_cordic/mycordic/N622 ) );
  NAND22 U3613 ( .A(\u_outFIFO/outWriteCount[2] ), .B(n181), .Q(n2306) );
  INV3 U3614 ( .A(\u_cordic/my_rotation/n94 ), .Q(n2226) );
  AOI221 U3615 ( .A(\u_cordic/my_rotation/present_delta [2]), .B(n33), .C(
        \u_cordic/my_rotation/present_delta [2]), .D(n748), .Q(
        \u_cordic/my_rotation/n94 ) );
  INV3 U3616 ( .A(\u_cordic/my_rotation/n96 ), .Q(n2228) );
  AOI221 U3617 ( .A(\u_cordic/my_rotation/present_delta [4]), .B(n33), .C(
        \u_cordic/my_rotation/N45 ), .D(n748), .Q(\u_cordic/my_rotation/n96 )
         );
  XOR21 U3618 ( .A(\u_cordic/my_rotation/present_delta [4]), .B(
        \u_cordic/my_rotation/present_delta [3]), .Q(
        \u_cordic/my_rotation/N45 ) );
  INV3 U3619 ( .A(\u_cordic/n28 ), .Q(n1673) );
  AOI221 U3620 ( .A(sig_MUX_outMUX7[3]), .B(\u_cordic/n20 ), .C(
        \u_cordic/Q [3]), .D(\u_cordic/n21 ), .Q(\u_cordic/n28 ) );
  NAND22 U3621 ( .A(sig_DEMUX_outDEMUX18[7]), .B(n1689), .Q(n2685) );
  INV3 U3622 ( .A(\u_cordic/n27 ), .Q(n1675) );
  AOI221 U3623 ( .A(sig_MUX_outMUX7[2]), .B(\u_cordic/n20 ), .C(
        \u_cordic/Q [2]), .D(\u_cordic/n21 ), .Q(\u_cordic/n27 ) );
  NAND22 U3624 ( .A(sig_DEMUX_outDEMUX18[6]), .B(n1689), .Q(n2683) );
  INV3 U3625 ( .A(\u_cordic/n26 ), .Q(n1677) );
  AOI221 U3626 ( .A(sig_MUX_outMUX7[1]), .B(\u_cordic/n20 ), .C(
        \u_cordic/Q [1]), .D(\u_cordic/n21 ), .Q(\u_cordic/n26 ) );
  NAND22 U3627 ( .A(sig_DEMUX_outDEMUX18[5]), .B(n1689), .Q(n2681) );
  INV3 U3628 ( .A(\u_cordic/n25 ), .Q(n1679) );
  AOI221 U3629 ( .A(sig_MUX_outMUX7[0]), .B(\u_cordic/n20 ), .C(
        \u_cordic/Q [0]), .D(\u_cordic/n21 ), .Q(\u_cordic/n25 ) );
  NAND22 U3630 ( .A(sig_DEMUX_outDEMUX18[4]), .B(n1689), .Q(n2679) );
  INV3 U3631 ( .A(\u_cordic/n24 ), .Q(n1665) );
  AOI221 U3632 ( .A(sig_MUX_outMUX6[3]), .B(\u_cordic/n20 ), .C(
        \u_cordic/I [3]), .D(\u_cordic/n21 ), .Q(\u_cordic/n24 ) );
  NAND22 U3633 ( .A(sig_DEMUX_outDEMUX17[7]), .B(n1689), .Q(n2677) );
  INV3 U3634 ( .A(\u_cordic/n23 ), .Q(n1667) );
  AOI221 U3635 ( .A(sig_MUX_outMUX6[2]), .B(\u_cordic/n20 ), .C(
        \u_cordic/I [2]), .D(\u_cordic/n21 ), .Q(\u_cordic/n23 ) );
  NAND22 U3636 ( .A(sig_DEMUX_outDEMUX17[6]), .B(n1689), .Q(n2675) );
  INV3 U3637 ( .A(\u_cordic/n22 ), .Q(n1669) );
  AOI221 U3638 ( .A(sig_MUX_outMUX6[1]), .B(\u_cordic/n20 ), .C(
        \u_cordic/I [1]), .D(\u_cordic/n21 ), .Q(\u_cordic/n22 ) );
  NAND22 U3639 ( .A(sig_DEMUX_outDEMUX17[5]), .B(n1689), .Q(n2673) );
  INV3 U3640 ( .A(\u_cordic/n19 ), .Q(n1671) );
  AOI221 U3641 ( .A(sig_MUX_outMUX6[0]), .B(\u_cordic/n20 ), .C(
        \u_cordic/I [0]), .D(\u_cordic/n21 ), .Q(\u_cordic/n19 ) );
  NAND22 U3642 ( .A(sig_DEMUX_outDEMUX17[4]), .B(n1689), .Q(n2671) );
  INV3 U3643 ( .A(n2277), .Q(n1722) );
  NOR21 U3644 ( .A(\u_coder/i [9]), .B(\u_coder/i [8]), .Q(n2277) );
  INV3 U3645 ( .A(\u_outFIFO/n503 ), .Q(n1331) );
  AOI221 U3646 ( .A(\u_outFIFO/n504 ), .B(\u_outFIFO/N39 ), .C(
        \u_outFIFO/n505 ), .D(\u_outFIFO/N199 ), .Q(\u_outFIFO/n503 ) );
  XOR21 U3647 ( .A(\u_outFIFO/add_360/carry [4]), .B(\u_outFIFO/N39 ), .Q(
        \u_outFIFO/N199 ) );
  INV3 U3648 ( .A(\u_inFIFO/n201 ), .Q(n1479) );
  AOI221 U3649 ( .A(\u_inFIFO/n202 ), .B(\u_inFIFO/N37 ), .C(\u_inFIFO/n203 ), 
        .D(\u_inFIFO/N121 ), .Q(\u_inFIFO/n201 ) );
  XOR21 U3650 ( .A(\u_inFIFO/add_253/carry [4]), .B(\u_inFIFO/N37 ), .Q(
        \u_inFIFO/N121 ) );
  XNR21 U3651 ( .A(\u_cordic/mycordic/r173/carry [5]), .B(n382), .Q(n381) );
  INV3 U3652 ( .A(\u_outFIFO/n207 ), .Q(n1326) );
  AOI221 U3653 ( .A(\u_outFIFO/N182 ), .B(\u_outFIFO/n208 ), .C(
        sig_outFIFO_outData[3]), .D(\u_outFIFO/n209 ), .Q(\u_outFIFO/n207 ) );
  INV3 U3654 ( .A(\u_outFIFO/n210 ), .Q(n1325) );
  AOI221 U3655 ( .A(\u_outFIFO/N183 ), .B(\u_outFIFO/n208 ), .C(
        sig_outFIFO_outData[2]), .D(\u_outFIFO/n209 ), .Q(\u_outFIFO/n210 ) );
  INV3 U3656 ( .A(\u_outFIFO/n211 ), .Q(n1324) );
  AOI221 U3657 ( .A(\u_outFIFO/N184 ), .B(\u_outFIFO/n208 ), .C(
        sig_outFIFO_outData[1]), .D(\u_outFIFO/n209 ), .Q(\u_outFIFO/n211 ) );
  INV3 U3658 ( .A(\u_outFIFO/n212 ), .Q(n1323) );
  AOI221 U3659 ( .A(\u_outFIFO/N185 ), .B(\u_outFIFO/n208 ), .C(
        sig_outFIFO_outData[0]), .D(\u_outFIFO/n209 ), .Q(\u_outFIFO/n212 ) );
  INV3 U3660 ( .A(\u_inFIFO/n228 ), .Q(n1480) );
  AOI221 U3661 ( .A(\u_inFIFO/N116 ), .B(n1652), .C(\u_inFIFO/outReadCount[4] ), .D(\u_inFIFO/n218 ), .Q(\u_inFIFO/n228 ) );
  XOR21 U3662 ( .A(\u_inFIFO/add_252/carry [4]), .B(\u_inFIFO/outReadCount[4] ), .Q(\u_inFIFO/N116 ) );
  INV3 U3663 ( .A(\u_inFIFO/n221 ), .Q(n1481) );
  AOI221 U3664 ( .A(n105), .B(n1652), .C(\u_inFIFO/outReadCount[0] ), .D(
        \u_inFIFO/n218 ), .Q(\u_inFIFO/n221 ) );
  INV3 U3665 ( .A(\u_inFIFO/n220 ), .Q(n1482) );
  AOI221 U3666 ( .A(\u_inFIFO/N113 ), .B(n1652), .C(\u_inFIFO/outReadCount[1] ), .D(\u_inFIFO/n218 ), .Q(\u_inFIFO/n220 ) );
  INV3 U3667 ( .A(\u_inFIFO/n219 ), .Q(n1483) );
  AOI221 U3668 ( .A(\u_inFIFO/N114 ), .B(n1652), .C(\u_inFIFO/outReadCount[2] ), .D(\u_inFIFO/n218 ), .Q(\u_inFIFO/n219 ) );
  INV3 U3669 ( .A(\u_inFIFO/n217 ), .Q(n1484) );
  AOI221 U3670 ( .A(\u_inFIFO/N115 ), .B(n1652), .C(\u_inFIFO/outReadCount[3] ), .D(\u_inFIFO/n218 ), .Q(\u_inFIFO/n217 ) );
  XNR21 U3671 ( .A(\u_cordic/mycordic/r173/carry [6]), .B(
        \u_cordic/mycordic/present_ANGLE_table[6][6] ), .Q(n383) );
  INV3 U3672 ( .A(\u_outFIFO/n524 ), .Q(n1465) );
  AOI221 U3673 ( .A(n154), .B(\u_outFIFO/n520 ), .C(
        \u_outFIFO/outReadCount[0] ), .D(n1466), .Q(\u_outFIFO/n524 ) );
  INV3 U3674 ( .A(\u_outFIFO/n523 ), .Q(n1464) );
  AOI221 U3675 ( .A(\u_outFIFO/N126 ), .B(\u_outFIFO/n520 ), .C(
        \u_outFIFO/outReadCount[1] ), .D(n1466), .Q(\u_outFIFO/n523 ) );
  INV3 U3676 ( .A(\u_outFIFO/n522 ), .Q(n1463) );
  AOI221 U3677 ( .A(\u_outFIFO/N127 ), .B(\u_outFIFO/n520 ), .C(
        \u_outFIFO/outReadCount[2] ), .D(n1466), .Q(\u_outFIFO/n522 ) );
  INV3 U3678 ( .A(\u_outFIFO/n521 ), .Q(n1462) );
  AOI221 U3679 ( .A(\u_outFIFO/N128 ), .B(\u_outFIFO/n520 ), .C(
        \u_outFIFO/outReadCount[3] ), .D(n1466), .Q(\u_outFIFO/n521 ) );
  INV3 U3680 ( .A(\u_outFIFO/n519 ), .Q(n1461) );
  AOI221 U3681 ( .A(\u_outFIFO/N129 ), .B(\u_outFIFO/n520 ), .C(
        \u_outFIFO/outReadCount[4] ), .D(n1466), .Q(\u_outFIFO/n519 ) );
  XOR21 U3682 ( .A(\u_outFIFO/add_260/carry [4]), .B(
        \u_outFIFO/outReadCount[4] ), .Q(\u_outFIFO/N129 ) );
  INV3 U3683 ( .A(\u_cordic/mycordic/n497 ), .Q(n1294) );
  AOI221 U3684 ( .A(\u_cordic/mycordic/N402 ), .B(n831), .C(
        \u_cordic/mycordic/N434 ), .D(n1582), .Q(\u_cordic/mycordic/n497 ) );
  XNR21 U3685 ( .A(\u_cordic/mycordic/present_ANGLE_table[2][6] ), .B(
        \u_cordic/mycordic/sub_207/carry [6]), .Q(\u_cordic/mycordic/N434 ) );
  XOR21 U3686 ( .A(\u_cordic/mycordic/present_ANGLE_table[2][6] ), .B(
        \u_cordic/mycordic/add_202/carry [6]), .Q(\u_cordic/mycordic/N402 ) );
  INV3 U3687 ( .A(\u_cordic/mycordic/n496 ), .Q(n1295) );
  AOI221 U3688 ( .A(\u_cordic/mycordic/N403 ), .B(n831), .C(
        \u_cordic/mycordic/N435 ), .D(n1582), .Q(\u_cordic/mycordic/n496 ) );
  XNR21 U3689 ( .A(\u_cordic/mycordic/present_ANGLE_table[2][7] ), .B(
        \u_cordic/mycordic/sub_207/carry [7]), .Q(\u_cordic/mycordic/N435 ) );
  XOR21 U3690 ( .A(\u_cordic/mycordic/present_ANGLE_table[2][7] ), .B(
        \u_cordic/mycordic/add_202/carry [7]), .Q(\u_cordic/mycordic/N403 ) );
  INV3 U3691 ( .A(\u_cordic/mycordic/n482 ), .Q(n1268) );
  AOI221 U3692 ( .A(\u_cordic/mycordic/N461 ), .B(n835), .C(
        \u_cordic/mycordic/N489 ), .D(n1581), .Q(\u_cordic/mycordic/n482 ) );
  XNR21 U3693 ( .A(\u_cordic/mycordic/present_ANGLE_table[3][5] ), .B(
        \u_cordic/mycordic/sub_218/carry[5] ), .Q(\u_cordic/mycordic/N489 ) );
  XOR21 U3694 ( .A(\u_cordic/mycordic/present_ANGLE_table[3][5] ), .B(
        \u_cordic/mycordic/add_213/carry[5] ), .Q(\u_cordic/mycordic/N461 ) );
  INV3 U3695 ( .A(\u_cordic/mycordic/n481 ), .Q(n1269) );
  AOI221 U3696 ( .A(\u_cordic/mycordic/N462 ), .B(n836), .C(
        \u_cordic/mycordic/N490 ), .D(n1581), .Q(\u_cordic/mycordic/n481 ) );
  XNR21 U3697 ( .A(\u_cordic/mycordic/present_ANGLE_table[3][6] ), .B(
        \u_cordic/mycordic/sub_218/carry[6] ), .Q(\u_cordic/mycordic/N490 ) );
  XOR21 U3698 ( .A(\u_cordic/mycordic/present_ANGLE_table[3][6] ), .B(
        \u_cordic/mycordic/add_213/carry[6] ), .Q(\u_cordic/mycordic/N462 ) );
  INV3 U3699 ( .A(\u_cordic/mycordic/n466 ), .Q(n1244) );
  AOI221 U3700 ( .A(\u_cordic/mycordic/N506 ), .B(n788), .C(
        \u_cordic/mycordic/N523 ), .D(n1580), .Q(\u_cordic/mycordic/n466 ) );
  XNR21 U3701 ( .A(\u_cordic/mycordic/present_ANGLE_table[4][5] ), .B(
        \u_cordic/mycordic/sub_229/carry[5] ), .Q(\u_cordic/mycordic/N523 ) );
  XOR21 U3702 ( .A(\u_cordic/mycordic/present_ANGLE_table[4][5] ), .B(
        \u_cordic/mycordic/add_224/carry[5] ), .Q(\u_cordic/mycordic/N506 ) );
  INV3 U3703 ( .A(\u_cordic/mycordic/n465 ), .Q(n1245) );
  AOI221 U3704 ( .A(\u_cordic/mycordic/N507 ), .B(n788), .C(
        \u_cordic/mycordic/N524 ), .D(n1580), .Q(\u_cordic/mycordic/n465 ) );
  XOR21 U3705 ( .A(\u_cordic/mycordic/present_ANGLE_table[4][6] ), .B(
        \u_cordic/mycordic/add_224/carry[6] ), .Q(\u_cordic/mycordic/N507 ) );
  XNR21 U3706 ( .A(\u_cordic/mycordic/present_ANGLE_table[4][6] ), .B(
        \u_cordic/mycordic/sub_229/carry[6] ), .Q(\u_cordic/mycordic/N524 ) );
  INV3 U3707 ( .A(\u_cordic/mycordic/n447 ), .Q(n1185) );
  AOI221 U3708 ( .A(\u_cordic/mycordic/N540 ), .B(n785), .C(
        \u_cordic/mycordic/N556 ), .D(n1577), .Q(\u_cordic/mycordic/n447 ) );
  XOR21 U3709 ( .A(\u_cordic/mycordic/present_ANGLE_table[5][6] ), .B(
        \u_cordic/mycordic/add_233/carry [6]), .Q(\u_cordic/mycordic/N540 ) );
  XNR21 U3710 ( .A(\u_cordic/mycordic/present_ANGLE_table[5][6] ), .B(
        \u_cordic/mycordic/sub_236/carry [6]), .Q(\u_cordic/mycordic/N556 ) );
  INV3 U3711 ( .A(\u_cordic/mycordic/n446 ), .Q(n1186) );
  AOI221 U3712 ( .A(\u_cordic/mycordic/N541 ), .B(n785), .C(
        \u_cordic/mycordic/N557 ), .D(n1577), .Q(\u_cordic/mycordic/n446 ) );
  XOR21 U3713 ( .A(\u_cordic/mycordic/present_ANGLE_table[5][7] ), .B(
        \u_cordic/mycordic/add_233/carry [7]), .Q(\u_cordic/mycordic/N541 ) );
  XNR21 U3714 ( .A(\u_cordic/mycordic/present_ANGLE_table[5][7] ), .B(
        \u_cordic/mycordic/sub_236/carry [7]), .Q(\u_cordic/mycordic/N557 ) );
  INV3 U3715 ( .A(\u_cordic/mycordic/n436 ), .Q(n1576) );
  NAND22 U3716 ( .A(\u_cordic/mycordic/next_ANGLE_table[6][0] ), .B(n970), .Q(
        \u_cordic/mycordic/n436 ) );
  INV3 U3717 ( .A(\u_cordic/mycordic/n424 ), .Q(n1567) );
  NAND22 U3718 ( .A(\u_cordic/mycordic/next_ANGLE_table[6][1] ), .B(n971), .Q(
        \u_cordic/mycordic/n424 ) );
  INV3 U3719 ( .A(\u_cordic/mycordic/n413 ), .Q(n1556) );
  NAND22 U3720 ( .A(\u_cordic/mycordic/next_ANGLE_table[6][2] ), .B(n971), .Q(
        \u_cordic/mycordic/n413 ) );
  INV3 U3721 ( .A(\u_cordic/mycordic/n411 ), .Q(n1554) );
  NAND22 U3722 ( .A(\u_cordic/mycordic/next_ANGLE_table[6][3] ), .B(n972), .Q(
        \u_cordic/mycordic/n411 ) );
  INV3 U3723 ( .A(\u_cordic/mycordic/n410 ), .Q(n1553) );
  NAND22 U3724 ( .A(\u_cordic/mycordic/next_ANGLE_table[6][4] ), .B(n972), .Q(
        \u_cordic/mycordic/n410 ) );
  INV3 U3725 ( .A(\u_cordic/mycordic/n409 ), .Q(n1552) );
  NAND22 U3726 ( .A(\u_cordic/mycordic/next_ANGLE_table[6][5] ), .B(n972), .Q(
        \u_cordic/mycordic/n409 ) );
  INV3 U3727 ( .A(\u_cordic/mycordic/n408 ), .Q(n1551) );
  NAND22 U3728 ( .A(\u_cordic/mycordic/next_ANGLE_table[6][6] ), .B(n972), .Q(
        \u_cordic/mycordic/n408 ) );
  NAND41 U3729 ( .A(\u_coder/n316 ), .B(\u_coder/n317 ), .C(\u_coder/n318 ), 
        .D(\u_coder/n319 ), .Q(\u_coder/n314 ) );
  NOR21 U3730 ( .A(\u_coder/c [14]), .B(\u_coder/c [13]), .Q(\u_coder/n316 )
         );
  NOR31 U3731 ( .A(\u_coder/c [15]), .B(\u_coder/c [17]), .C(\u_coder/c [16]), 
        .Q(\u_coder/n317 ) );
  NOR40 U3732 ( .A(\u_coder/n324 ), .B(\u_coder/c [10]), .C(\u_coder/c [12]), 
        .D(\u_coder/c [11]), .Q(\u_coder/n318 ) );
  NAND22 U3733 ( .A(\u_inFIFO/n98 ), .B(\u_inFIFO/n97 ), .Q(\u_inFIFO/n121 )
         );
  NAND22 U3734 ( .A(\u_inFIFO/j_FIFO [4]), .B(\u_inFIFO/j_FIFO [3]), .Q(
        \u_inFIFO/n179 ) );
  NAND22 U3735 ( .A(\u_inFIFO/j_FIFO [3]), .B(\u_inFIFO/n97 ), .Q(
        \u_inFIFO/n145 ) );
  NAND22 U3736 ( .A(\u_inFIFO/j_FIFO [4]), .B(\u_inFIFO/n98 ), .Q(
        \u_inFIFO/n162 ) );
  OAI2111 U3737 ( .A(\u_coder/i [2]), .B(n778), .C(\u_coder/i [1]), .D(
        \u_coder/n197 ), .Q(\u_coder/n194 ) );
  AOI211 U3738 ( .A(n778), .B(\u_coder/i [2]), .C(\u_coder/i [3]), .Q(
        \u_coder/n197 ) );
  OAI2111 U3739 ( .A(\u_coder/j [2]), .B(n777), .C(\u_coder/j [1]), .D(
        \u_coder/n242 ), .Q(\u_coder/n239 ) );
  AOI211 U3740 ( .A(n777), .B(\u_coder/j [2]), .C(n776), .Q(\u_coder/n242 ) );
  NAND31 U3741 ( .A(n746), .B(\u_decoder/iq_demod/cossin_dig/n23 ), .C(n976), 
        .Q(\u_decoder/iq_demod/cossin_dig/n44 ) );
  INV6 U3742 ( .A(\u_cordic/mycordic/n554 ), .Q(n1582) );
  NAND22 U3743 ( .A(\u_cordic/mycordic/present_Q_table[3][7] ), .B(n969), .Q(
        \u_cordic/mycordic/n554 ) );
  INV6 U3744 ( .A(\u_cordic/mycordic/n520 ), .Q(n1578) );
  NAND22 U3745 ( .A(\u_cordic/mycordic/present_Q_table[2][7] ), .B(n970), .Q(
        \u_cordic/mycordic/n520 ) );
  NOR40 U3746 ( .A(\u_cordic/mycordic/present_Q_table[0][3] ), .B(
        \u_cordic/mycordic/present_Q_table[0][4] ), .C(n2221), .D(n1169), .Q(
        \u_cordic/mycordic/N212 ) );
  INV3 U3747 ( .A(n784), .Q(n1169) );
  INV3 U3748 ( .A(\u_cordic/mycordic/n435 ), .Q(n2221) );
  NOR31 U3749 ( .A(\u_cordic/mycordic/present_Q_table[0][5] ), .B(
        \u_cordic/mycordic/present_Q_table[0][7] ), .C(
        \u_cordic/mycordic/present_Q_table[0][6] ), .Q(
        \u_cordic/mycordic/n435 ) );
  OAI2111 U3750 ( .A(\u_coder/n89 ), .B(\u_coder/n85 ), .C(\u_coder/n178 ), 
        .D(\u_coder/n88 ), .Q(\u_coder/n173 ) );
  NOR31 U3751 ( .A(\u_outFIFO/n176 ), .B(\u_outFIFO/currentState [0]), .C(
        \u_outFIFO/n546 ), .Q(\u_outFIFO/n539 ) );
  NOR21 U3752 ( .A(\u_outFIFO/n195 ), .B(\u_outFIFO/k_FIFO [0]), .Q(
        \u_outFIFO/n288 ) );
  NOR21 U3753 ( .A(\u_outFIFO/n196 ), .B(\u_outFIFO/k_FIFO [1]), .Q(
        \u_outFIFO/n291 ) );
  NAND22 U3754 ( .A(sig_DEMUX_outDEMUX2[2]), .B(n1689), .Q(\u_mux8/n3 ) );
  AOI221 U3755 ( .A(\sig_MUX_inMUX8[0] ), .B(n1689), .C(in_MUX_inSEL6[0]), .D(
        sig_DEMUX_outDEMUX2[2]), .Q(\u_mux8/n4 ) );
  NOR31 U3756 ( .A(n2693), .B(in_DEMUX_inSEL2[2]), .C(n1685), .Q(
        sig_DEMUX_outDEMUX2[2]) );
  NOR21 U3757 ( .A(n984), .B(\u_cordic/mycordic/present_Q_table[3][7] ), .Q(
        \u_cordic/mycordic/n332 ) );
  XNR21 U3758 ( .A(\u_decoder/iq_demod/cossin_dig/n19 ), .B(
        \u_decoder/iq_demod/cossin_dig/n21 ), .Q(
        \u_decoder/iq_demod/cossin_dig/n54 ) );
  NOR21 U3759 ( .A(\u_decoder/iq_demod/cossin_dig/n23 ), .B(n746), .Q(
        \u_decoder/iq_demod/cossin_dig/n26 ) );
  NOR21 U3760 ( .A(\u_outFIFO/i_FIFO [4]), .B(\u_outFIFO/i_FIFO [3]), .Q(
        \u_outFIFO/n285 ) );
  NOR31 U3761 ( .A(\u_cdr/cnt_in [1]), .B(\u_cdr/cnt_in [3]), .C(
        \u_cdr/cnt_in [0]), .Q(\u_cdr/n42 ) );
  INV3 U3762 ( .A(\u_cdr/n32 ), .Q(n1470) );
  NOR31 U3763 ( .A(\u_outFIFO/n177 ), .B(\u_outFIFO/n176 ), .C(
        \u_outFIFO/n546 ), .Q(\u_outFIFO/n537 ) );
  NOR21 U3764 ( .A(\u_outFIFO/k_FIFO [0]), .B(\u_outFIFO/k_FIFO [1]), .Q(
        \u_outFIFO/n294 ) );
  NAND31 U3765 ( .A(\u_cdr/cnt_d [1]), .B(\u_cdr/cnt_d [0]), .C(\u_cdr/flag ), 
        .Q(\u_cdr/n37 ) );
  NOR21 U3766 ( .A(n154), .B(\u_outFIFO/outWriteCount[0] ), .Q(n2310) );
  NAND22 U3767 ( .A(\u_outFIFO/n173 ), .B(\u_outFIFO/n174 ), .Q(
        \u_outFIFO/n546 ) );
  NOR21 U3768 ( .A(n981), .B(\u_cordic/mycordic/present_Q_table[2][7] ), .Q(
        \u_cordic/mycordic/n336 ) );
  NAND31 U3769 ( .A(\u_inFIFO/currentState [0]), .B(\u_inFIFO/n76 ), .C(n1698), 
        .Q(\u_inFIFO/n236 ) );
  NOR21 U3770 ( .A(\u_cordic/n11 ), .B(\u_cordic/n13 ), .Q(\u_cordic/n18 ) );
  NAND22 U3771 ( .A(\u_cdr/cnt_in [2]), .B(\u_cdr/N100 ), .Q(
        \u_cdr/dp_cluster_0/mult_add_59_aco/PROD_not[2] ) );
  BUF6 U3772 ( .A(\u_decoder/iq_demod/n42 ), .Q(n790) );
  NOR21 U3773 ( .A(\u_decoder/iq_demod/n30 ), .B(n752), .Q(
        \u_decoder/iq_demod/n42 ) );
  NAND31 U3774 ( .A(\u_outFIFO/i_FIFO [1]), .B(\u_outFIFO/i_FIFO [0]), .C(
        \u_outFIFO/i_FIFO [2]), .Q(\u_outFIFO/n284 ) );
  NAND31 U3775 ( .A(\u_outFIFO/i_FIFO [1]), .B(\u_outFIFO/n194 ), .C(
        \u_outFIFO/i_FIFO [2]), .Q(\u_outFIFO/n275 ) );
  NAND31 U3776 ( .A(\u_outFIFO/i_FIFO [0]), .B(\u_outFIFO/n193 ), .C(
        \u_outFIFO/i_FIFO [2]), .Q(\u_outFIFO/n266 ) );
  NAND31 U3777 ( .A(\u_outFIFO/n194 ), .B(\u_outFIFO/n193 ), .C(
        \u_outFIFO/i_FIFO [2]), .Q(\u_outFIFO/n257 ) );
  NOR21 U3778 ( .A(\u_outFIFO/n191 ), .B(\u_outFIFO/i_FIFO [4]), .Q(
        \u_outFIFO/n357 ) );
  NAND31 U3779 ( .A(\u_outFIFO/n193 ), .B(\u_outFIFO/n192 ), .C(
        \u_outFIFO/i_FIFO [0]), .Q(\u_outFIFO/n230 ) );
  NOR21 U3780 ( .A(\u_outFIFO/n185 ), .B(\u_outFIFO/i_FIFO [3]), .Q(
        \u_outFIFO/n426 ) );
  NOR21 U3781 ( .A(\u_outFIFO/n185 ), .B(\u_outFIFO/n191 ), .Q(
        \u_outFIFO/n495 ) );
  NAND31 U3782 ( .A(\u_outFIFO/i_FIFO [0]), .B(\u_outFIFO/n192 ), .C(
        \u_outFIFO/i_FIFO [1]), .Q(\u_outFIFO/n248 ) );
  NAND31 U3783 ( .A(\u_outFIFO/n194 ), .B(\u_outFIFO/n192 ), .C(
        \u_outFIFO/i_FIFO [1]), .Q(\u_outFIFO/n239 ) );
  OAI2111 U3784 ( .A(\u_cordic/mycordic/present_Q_table[0][7] ), .B(
        \u_cordic/mycordic/n391 ), .C(\u_cordic/mycordic/n432 ), .D(n1167), 
        .Q(\u_cordic/mycordic/N211 ) );
  NAND22 U3785 ( .A(\u_cordic/mycordic/present_Q_table[0][7] ), .B(n784), .Q(
        \u_cordic/mycordic/n432 ) );
  INV3 U3786 ( .A(\u_cordic/mycordic/N212 ), .Q(n1167) );
  NAND31 U3787 ( .A(\u_outFIFO/n193 ), .B(\u_outFIFO/n192 ), .C(
        \u_outFIFO/n194 ), .Q(\u_outFIFO/n217 ) );
  NOR21 U3788 ( .A(\u_decoder/iq_demod/cossin_dig/n44 ), .B(
        \u_decoder/iq_demod/cossin_dig/counter [0]), .Q(
        \u_decoder/iq_demod/cossin_dig/N20 ) );
  NOR40 U3789 ( .A(\u_coder/n320 ), .B(n1773), .C(\u_coder/c [19]), .D(
        \u_coder/c [18]), .Q(\u_coder/n319 ) );
  INV3 U3790 ( .A(\u_coder/n321 ), .Q(n1773) );
  NAND22 U3791 ( .A(\u_coder/n322 ), .B(\u_coder/n323 ), .Q(\u_coder/n320 ) );
  NOR31 U3792 ( .A(\u_coder/c [1]), .B(\u_coder/c [4]), .C(\u_coder/c [3]), 
        .Q(\u_coder/n321 ) );
  NOR31 U3793 ( .A(\u_coder/c [7]), .B(\u_coder/c [9]), .C(\u_coder/c [8]), 
        .Q(\u_coder/n323 ) );
  INV3 U3794 ( .A(\u_decoder/iq_demod/cossin_dig/n39 ), .Q(n1504) );
  INV3 U3795 ( .A(\u_cordic/mycordic/n355 ), .Q(n1177) );
  AOI221 U3796 ( .A(n1575), .B(\u_cordic/mycordic/N246 ), .C(n784), .D(
        \u_cordic/mycordic/present_Q_table[0][6] ), .Q(
        \u_cordic/mycordic/n355 ) );
  XOR21 U3797 ( .A(\u_cordic/mycordic/sub_add_151_b0/carry [6]), .B(n41), .Q(
        \u_cordic/mycordic/N246 ) );
  NAND22 U3798 ( .A(\u_cdr/N100 ), .B(\u_cdr/cnt_in [3]), .Q(
        \u_cdr/dp_cluster_0/mult_add_59_aco/PROD_not[3] ) );
  NAND31 U3799 ( .A(n978), .B(\u_cdr/n37 ), .C(\u_cdr/flag ), .Q(\u_cdr/n34 )
         );
  INV3 U3800 ( .A(\u_outFIFO/N120 ), .Q(n1799) );
  INV3 U3801 ( .A(\u_outFIFO/N121 ), .Q(n1798) );
  NOR21 U3802 ( .A(\u_outFIFO/n288 ), .B(\u_outFIFO/n291 ), .Q(
        \u_outFIFO/n510 ) );
  NOR21 U3803 ( .A(\u_inFIFO/n76 ), .B(\u_inFIFO/currentState [0]), .Q(
        \u_inFIFO/n106 ) );
  NAND22 U3804 ( .A(\u_cordic/n16 ), .B(\u_cordic/n17 ), .Q(\u_cordic/n37 ) );
  NAND31 U3805 ( .A(\u_cordic/n18 ), .B(\u_cordic/n12 ), .C(\u_cordic/dir ), 
        .Q(\u_cordic/n17 ) );
  XNR21 U3806 ( .A(\u_inFIFO/n93 ), .B(\u_inFIFO/n94 ), .Q(\u_inFIFO/n208 ) );
  NAND22 U3807 ( .A(\u_inFIFO/sigEnableCounter ), .B(n969), .Q(\u_inFIFO/n227 ) );
  OAI311 U3808 ( .A(\u_decoder/fir_filter/n1150 ), .B(
        \u_decoder/fir_filter/n1149 ), .C(\u_decoder/fir_filter/n1151 ), .D(
        \u_decoder/fir_filter/n1152 ), .Q(\u_decoder/fir_filter/n1451 ) );
  NAND22 U3809 ( .A(\sig_MUX_inMUX8[0] ), .B(\u_decoder/fir_filter/n1150 ), 
        .Q(\u_decoder/fir_filter/n1152 ) );
  NOR21 U3810 ( .A(n933), .B(\u_decoder/fir_filter/n1151 ), .Q(
        \u_decoder/fir_filter/n1150 ) );
  OAI311 U3811 ( .A(\u_decoder/iq_demod/cossin_dig/n43 ), .B(
        \u_decoder/iq_demod/cossin_dig/counter [2]), .C(
        \u_decoder/iq_demod/cossin_dig/n44 ), .D(
        \u_decoder/iq_demod/cossin_dig/n46 ), .Q(
        \u_decoder/iq_demod/cossin_dig/N22 ) );
  NOR21 U3812 ( .A(\u_decoder/iq_demod/cossin_dig/counter [1]), .B(
        \u_decoder/iq_demod/cossin_dig/n44 ), .Q(
        \u_decoder/iq_demod/cossin_dig/n47 ) );
  NOR21 U3813 ( .A(n814), .B(\u_coder/c [0]), .Q(\u_coder/N503 ) );
  BUF2 U3814 ( .A(\u_cordic/mycordic/n108 ), .Q(n751) );
  NAND22 U3815 ( .A(n1720), .B(\u_coder/n85 ), .Q(\u_coder/n163 ) );
  NAND22 U3816 ( .A(\u_inFIFO/n26 ), .B(\u_inFIFO/n73 ), .Q(\u_inFIFO/n241 )
         );
  AOI311 U3817 ( .A(\u_inFIFO/n240 ), .B(\u_inFIFO/n26 ), .C(\u_inFIFO/n230 ), 
        .D(\u_inFIFO/n233 ), .Q(\u_inFIFO/n238 ) );
  XOR21 U3818 ( .A(\u_inFIFO/sig_fsm_start_R ), .B(\u_inFIFO/sig_fsm_start_W ), 
        .Q(\u_inFIFO/n240 ) );
  NOR21 U3819 ( .A(\u_inFIFO/os2/sigQout2 ), .B(n290), .Q(
        \u_inFIFO/sig_fsm_start_W ) );
  AOI311 U3820 ( .A(n1790), .B(\u_outFIFO/n173 ), .C(
        \u_outFIFO/sig_fsm_start_R ), .D(\u_outFIFO/n539 ), .Q(
        \u_outFIFO/n548 ) );
  INV3 U3821 ( .A(\u_outFIFO/n534 ), .Q(n1790) );
  NAND41 U3822 ( .A(\u_cdr/cnt [1]), .B(\u_cdr/cnt [0]), .C(\u_cdr/n32 ), .D(
        \u_cdr/n16 ), .Q(\u_cdr/n36 ) );
  AOI211 U3823 ( .A(\u_cdr/n32 ), .B(\u_cdr/n17 ), .C(\u_cdr/n33 ), .Q(
        \u_cdr/n35 ) );
  BUF2 U3824 ( .A(\u_decoder/iq_demod/cossin_dig/state[0] ), .Q(n746) );
  NAND31 U3825 ( .A(\u_cdr/n32 ), .B(\u_cdr/n17 ), .C(\u_cdr/cnt [0]), .Q(
        \u_cdr/n31 ) );
  INV3 U3826 ( .A(\u_cdr/n33 ), .Q(n1469) );
  NOR21 U3827 ( .A(\u_decoder/iq_demod/cossin_dig/n56 ), .B(
        \u_decoder/iq_demod/cossin_dig/n31 ), .Q(
        \u_decoder/iq_demod/cossin_dig/n34 ) );
  AOI211 U3828 ( .A(\u_cordic/n32 ), .B(\u_cordic/n33 ), .C(n986), .Q(
        \u_cordic/N16 ) );
  OAI2111 U3829 ( .A(sig_MUX_outMUX8), .B(\u_cordic/n11 ), .C(\u_cordic/n13 ), 
        .D(\u_cordic/present_state [1]), .Q(\u_cordic/n33 ) );
  NAND22 U3830 ( .A(\u_cordic/n34 ), .B(\u_cordic/n12 ), .Q(\u_cordic/n32 ) );
  BUF2 U3831 ( .A(\u_cordic/mycordic/n354 ), .Q(n784) );
  NOR21 U3832 ( .A(n983), .B(\u_cordic/mycordic/present_I_table[0][7] ), .Q(
        \u_cordic/mycordic/n354 ) );
  BUF2 U3833 ( .A(\u_decoder/iq_demod/state [1]), .Q(n752) );
  INV3 U3834 ( .A(\u_cordic/mycordic/n516 ), .Q(n1198) );
  AOI221 U3835 ( .A(\u_cordic/mycordic/N335 ), .B(n833), .C(
        \u_cordic/mycordic/N367 ), .D(n1578), .Q(\u_cordic/mycordic/n516 ) );
  XOR21 U3836 ( .A(\u_cordic/mycordic/present_ANGLE_table[1][3] ), .B(
        \u_cordic/mycordic/sub_196/carry[3] ), .Q(\u_cordic/mycordic/N367 ) );
  XNR21 U3837 ( .A(\u_cordic/mycordic/present_ANGLE_table[1][3] ), .B(
        \u_cordic/mycordic/add_191/carry[3] ), .Q(\u_cordic/mycordic/N335 ) );
  NOR21 U3838 ( .A(\u_cordic/mycordic/n391 ), .B(n39), .Q(
        \u_cordic/mycordic/N44 ) );
  BUF2 U3839 ( .A(\u_outFIFO/N37 ), .Q(n774) );
  BUF2 U3840 ( .A(\u_inFIFO/N35 ), .Q(n779) );
  XOR21 U3841 ( .A(\u_cordic/mycordic/present_ANGLE_table[6][3] ), .B(
        \u_cordic/mycordic/present_ANGLE_table[6][4] ), .Q(
        \u_cordic/mycordic/N619 ) );
  XNR21 U3842 ( .A(\u_cordic/mycordic/add_262/carry [5]), .B(
        \u_cordic/mycordic/present_ANGLE_table[6][5] ), .Q(
        \u_cordic/mycordic/N620 ) );
  NOR21 U3843 ( .A(\u_outFIFO/os2/sigQout2 ), .B(n291), .Q(
        \u_outFIFO/sig_fsm_start_W ) );
  NAND22 U3844 ( .A(\u_coder/c [2]), .B(\u_coder/n33 ), .Q(\u_coder/n324 ) );
  NOR21 U3845 ( .A(\u_coder/c [6]), .B(\u_coder/c [5]), .Q(\u_coder/n322 ) );
  INV3 U3846 ( .A(\u_inFIFO/n239 ), .Q(n1486) );
  INV3 U3847 ( .A(n2270), .Q(n1754) );
  NOR21 U3848 ( .A(\u_coder/j [9]), .B(\u_coder/j [8]), .Q(n2270) );
  INV3 U3849 ( .A(\u_outFIFO/n549 ), .Q(n1585) );
  NOR21 U3850 ( .A(\u_outFIFO/os1/sigQout2 ), .B(n292), .Q(
        \u_outFIFO/sig_fsm_start_R ) );
  XNR21 U3851 ( .A(\u_cordic/mycordic/r173/carry [4]), .B(n385), .Q(n384) );
  XNR21 U3852 ( .A(\u_cordic/mycordic/present_ANGLE_table[6][2] ), .B(
        \u_cordic/mycordic/present_ANGLE_table[6][3] ), .Q(n386) );
  INV3 U3853 ( .A(\u_cordic/mycordic/n433 ), .Q(n1168) );
  AOI211 U3854 ( .A(n978), .B(\u_cordic/mycordic/present_Q_table[0][7] ), .C(
        \u_cordic/mycordic/N212 ), .Q(\u_cordic/mycordic/n433 ) );
  INV3 U3855 ( .A(\u_decoder/iq_demod/cossin_dig/n36 ), .Q(n2247) );
  AOI221 U3856 ( .A(\u_decoder/iq_demod/cossin_dig/N60 ), .B(n2248), .C(
        \u_decoder/iq_demod/sin_out [3]), .D(n746), .Q(
        \u_decoder/iq_demod/cossin_dig/n36 ) );
  INV3 U3857 ( .A(\u_decoder/iq_demod/cossin_dig/n31 ), .Q(n2248) );
  INV3 U3858 ( .A(\u_decoder/iq_demod/cossin_dig/n35 ), .Q(n2246) );
  AOI211 U3859 ( .A(\u_decoder/iq_demod/sin_out [2]), .B(n746), .C(
        \u_decoder/iq_demod/cossin_dig/n34 ), .Q(
        \u_decoder/iq_demod/cossin_dig/n35 ) );
  INV3 U3860 ( .A(\u_decoder/iq_demod/cossin_dig/n33 ), .Q(n2245) );
  AOI211 U3861 ( .A(\u_decoder/iq_demod/sin_out [1]), .B(n746), .C(
        \u_decoder/iq_demod/cossin_dig/n34 ), .Q(
        \u_decoder/iq_demod/cossin_dig/n33 ) );
  INV3 U3862 ( .A(\u_cordic/mycordic/n334 ), .Q(n1312) );
  AOI221 U3863 ( .A(\u_cordic/mycordic/N388 ), .B(n832), .C(
        \u_cordic/mycordic/N420 ), .D(n1582), .Q(\u_cordic/mycordic/n334 ) );
  XOR21 U3864 ( .A(\u_cordic/mycordic/present_Q_table[3][0] ), .B(
        \u_cordic/mycordic/present_I_table[3][2] ), .Q(
        \u_cordic/mycordic/N420 ) );
  XNR21 U3865 ( .A(\u_cordic/mycordic/present_Q_table[3][0] ), .B(n157), .Q(
        \u_cordic/mycordic/N388 ) );
  INV3 U3866 ( .A(\u_cordic/mycordic/n374 ), .Q(n1304) );
  AOI221 U3867 ( .A(\u_cordic/mycordic/N380 ), .B(\u_cordic/mycordic/n332 ), 
        .C(\u_cordic/mycordic/N412 ), .D(n1582), .Q(\u_cordic/mycordic/n374 )
         );
  XOR21 U3868 ( .A(\u_cordic/mycordic/present_I_table[3][0] ), .B(
        \u_cordic/mycordic/present_Q_table[3][2] ), .Q(
        \u_cordic/mycordic/N380 ) );
  XNR21 U3869 ( .A(\u_cordic/mycordic/present_I_table[3][0] ), .B(n158), .Q(
        \u_cordic/mycordic/N412 ) );
  INV3 U3870 ( .A(\u_cordic/mycordic/n503 ), .Q(n1288) );
  AOI221 U3871 ( .A(\u_cordic/mycordic/N428 ), .B(n831), .C(
        \u_cordic/mycordic/N428 ), .D(n1582), .Q(\u_cordic/mycordic/n503 ) );
  INV3 U3872 ( .A(\u_cordic/mycordic/n502 ), .Q(n1289) );
  AOI221 U3873 ( .A(n297), .B(n831), .C(n297), .D(n1582), .Q(
        \u_cordic/mycordic/n502 ) );
  INV3 U3874 ( .A(\u_cordic/mycordic/n501 ), .Q(n1290) );
  AOI221 U3875 ( .A(\u_cordic/mycordic/N398 ), .B(n831), .C(
        \u_cordic/mycordic/N430 ), .D(n1582), .Q(\u_cordic/mycordic/n501 ) );
  XOR21 U3876 ( .A(\u_cordic/mycordic/present_ANGLE_table[2][2] ), .B(
        \u_cordic/mycordic/present_ANGLE_table[2][1] ), .Q(
        \u_cordic/mycordic/N430 ) );
  XNR21 U3877 ( .A(\u_cordic/mycordic/present_ANGLE_table[2][2] ), .B(
        \u_cordic/mycordic/present_ANGLE_table[2][1] ), .Q(
        \u_cordic/mycordic/N398 ) );
  INV3 U3878 ( .A(\u_cordic/mycordic/n500 ), .Q(n1291) );
  AOI221 U3879 ( .A(\u_cordic/mycordic/N399 ), .B(n831), .C(
        \u_cordic/mycordic/N431 ), .D(n1582), .Q(\u_cordic/mycordic/n500 ) );
  XOR21 U3880 ( .A(\u_cordic/mycordic/present_ANGLE_table[2][3] ), .B(
        \u_cordic/mycordic/sub_207/carry [3]), .Q(\u_cordic/mycordic/N431 ) );
  XNR21 U3881 ( .A(\u_cordic/mycordic/present_ANGLE_table[2][3] ), .B(
        \u_cordic/mycordic/add_202/carry [3]), .Q(\u_cordic/mycordic/N399 ) );
  INV3 U3882 ( .A(\u_cordic/mycordic/n499 ), .Q(n1292) );
  AOI221 U3883 ( .A(\u_cordic/mycordic/N400 ), .B(n831), .C(
        \u_cordic/mycordic/N432 ), .D(n1582), .Q(\u_cordic/mycordic/n499 ) );
  XNR21 U3884 ( .A(\u_cordic/mycordic/present_ANGLE_table[2][4] ), .B(
        \u_cordic/mycordic/sub_207/carry [4]), .Q(\u_cordic/mycordic/N432 ) );
  XOR21 U3885 ( .A(\u_cordic/mycordic/present_ANGLE_table[2][4] ), .B(
        \u_cordic/mycordic/add_202/carry [4]), .Q(\u_cordic/mycordic/N400 ) );
  INV3 U3886 ( .A(\u_cordic/mycordic/n498 ), .Q(n1293) );
  AOI221 U3887 ( .A(\u_cordic/mycordic/N401 ), .B(n831), .C(
        \u_cordic/mycordic/N433 ), .D(n1582), .Q(\u_cordic/mycordic/n498 ) );
  XNR21 U3888 ( .A(\u_cordic/mycordic/present_ANGLE_table[2][5] ), .B(
        \u_cordic/mycordic/sub_207/carry [5]), .Q(\u_cordic/mycordic/N433 ) );
  XOR21 U3889 ( .A(\u_cordic/mycordic/present_ANGLE_table[2][5] ), .B(
        \u_cordic/mycordic/add_202/carry [5]), .Q(\u_cordic/mycordic/N401 ) );
  INV3 U3890 ( .A(\u_cordic/mycordic/n382 ), .Q(n1211) );
  AOI221 U3891 ( .A(\u_cordic/mycordic/N316 ), .B(\u_cordic/mycordic/n336 ), 
        .C(\u_cordic/mycordic/N348 ), .D(n1578), .Q(\u_cordic/mycordic/n382 )
         );
  XOR21 U3892 ( .A(\u_cordic/mycordic/present_I_table[2][0] ), .B(
        \u_cordic/mycordic/present_Q_table[2][1] ), .Q(
        \u_cordic/mycordic/N316 ) );
  XNR21 U3893 ( .A(\u_cordic/mycordic/present_I_table[2][0] ), .B(n159), .Q(
        \u_cordic/mycordic/N348 ) );
  INV3 U3894 ( .A(\u_cordic/mycordic/n343 ), .Q(n1219) );
  AOI221 U3895 ( .A(\u_cordic/mycordic/N324 ), .B(\u_cordic/mycordic/n336 ), 
        .C(\u_cordic/mycordic/N356 ), .D(n1578), .Q(\u_cordic/mycordic/n343 )
         );
  XOR21 U3896 ( .A(\u_cordic/mycordic/present_Q_table[2][0] ), .B(
        \u_cordic/mycordic/present_I_table[2][1] ), .Q(
        \u_cordic/mycordic/N356 ) );
  XNR21 U3897 ( .A(\u_cordic/mycordic/present_Q_table[2][0] ), .B(n160), .Q(
        \u_cordic/mycordic/N324 ) );
  INV3 U3898 ( .A(\u_cordic/mycordic/n519 ), .Q(n1195) );
  AOI221 U3899 ( .A(n298), .B(n833), .C(n298), .D(n1578), .Q(
        \u_cordic/mycordic/n519 ) );
  INV3 U3900 ( .A(\u_cordic/mycordic/n518 ), .Q(n1196) );
  AOI221 U3901 ( .A(\u_cordic/mycordic/N333 ), .B(n833), .C(
        \u_cordic/mycordic/N365 ), .D(n1578), .Q(\u_cordic/mycordic/n518 ) );
  XOR21 U3902 ( .A(\u_cordic/mycordic/present_ANGLE_table[1][1] ), .B(
        \u_cordic/mycordic/present_ANGLE_table[1][0] ), .Q(
        \u_cordic/mycordic/N365 ) );
  XNR21 U3903 ( .A(\u_cordic/mycordic/present_ANGLE_table[1][1] ), .B(
        \u_cordic/mycordic/present_ANGLE_table[1][0] ), .Q(
        \u_cordic/mycordic/N333 ) );
  INV3 U3904 ( .A(\u_cordic/mycordic/n517 ), .Q(n1197) );
  AOI221 U3905 ( .A(\u_cordic/mycordic/N334 ), .B(n833), .C(
        \u_cordic/mycordic/N366 ), .D(n1578), .Q(\u_cordic/mycordic/n517 ) );
  XNR21 U3906 ( .A(\u_cordic/mycordic/present_ANGLE_table[1][2] ), .B(
        \u_cordic/mycordic/sub_196/carry[2] ), .Q(\u_cordic/mycordic/N366 ) );
  XOR21 U3907 ( .A(\u_cordic/mycordic/present_ANGLE_table[1][2] ), .B(
        \u_cordic/mycordic/add_191/carry[2] ), .Q(\u_cordic/mycordic/N334 ) );
  INV3 U3908 ( .A(\u_cordic/mycordic/n515 ), .Q(n1199) );
  AOI221 U3909 ( .A(\u_cordic/mycordic/N336 ), .B(n833), .C(
        \u_cordic/mycordic/N368 ), .D(n1578), .Q(\u_cordic/mycordic/n515 ) );
  XOR21 U3910 ( .A(\u_cordic/mycordic/present_ANGLE_table[1][4] ), .B(
        \u_cordic/mycordic/sub_196/carry[4] ), .Q(\u_cordic/mycordic/N368 ) );
  XNR21 U3911 ( .A(\u_cordic/mycordic/present_ANGLE_table[1][4] ), .B(
        \u_cordic/mycordic/add_191/carry[4] ), .Q(\u_cordic/mycordic/N336 ) );
  XNR21 U3912 ( .A(\u_cordic/mycordic/present_Q_table[0][7] ), .B(
        \u_cordic/mycordic/sub_add_151_b0/carry [7]), .Q(
        \u_cordic/mycordic/N247 ) );
  INV3 U3913 ( .A(\u_cordic/mycordic/n484 ), .Q(n1266) );
  AOI221 U3914 ( .A(\u_cordic/mycordic/N459 ), .B(n835), .C(
        \u_cordic/mycordic/N487 ), .D(n1581), .Q(\u_cordic/mycordic/n484 ) );
  XNR21 U3915 ( .A(\u_cordic/mycordic/present_ANGLE_table[3][3] ), .B(
        \u_cordic/mycordic/sub_218/carry[3] ), .Q(\u_cordic/mycordic/N487 ) );
  XOR21 U3916 ( .A(\u_cordic/mycordic/present_ANGLE_table[3][3] ), .B(
        \u_cordic/mycordic/add_213/carry[3] ), .Q(\u_cordic/mycordic/N459 ) );
  INV3 U3917 ( .A(\u_cordic/mycordic/n483 ), .Q(n1267) );
  AOI221 U3918 ( .A(\u_cordic/mycordic/N460 ), .B(n835), .C(
        \u_cordic/mycordic/N488 ), .D(n1581), .Q(\u_cordic/mycordic/n483 ) );
  XNR21 U3919 ( .A(\u_cordic/mycordic/present_ANGLE_table[3][4] ), .B(
        \u_cordic/mycordic/sub_218/carry[4] ), .Q(\u_cordic/mycordic/N488 ) );
  XOR21 U3920 ( .A(\u_cordic/mycordic/present_ANGLE_table[3][4] ), .B(
        \u_cordic/mycordic/add_213/carry[4] ), .Q(\u_cordic/mycordic/N460 ) );
  INV3 U3921 ( .A(\u_cordic/mycordic/n468 ), .Q(n1242) );
  AOI221 U3922 ( .A(\u_cordic/mycordic/N504 ), .B(n788), .C(
        \u_cordic/mycordic/N521 ), .D(n1580), .Q(\u_cordic/mycordic/n468 ) );
  XNR21 U3923 ( .A(\u_cordic/mycordic/present_ANGLE_table[4][3] ), .B(
        \u_cordic/mycordic/sub_229/carry[3] ), .Q(\u_cordic/mycordic/N521 ) );
  XOR21 U3924 ( .A(\u_cordic/mycordic/present_ANGLE_table[4][3] ), .B(
        \u_cordic/mycordic/add_224/carry[3] ), .Q(\u_cordic/mycordic/N504 ) );
  INV3 U3925 ( .A(\u_cordic/mycordic/n467 ), .Q(n1243) );
  AOI221 U3926 ( .A(\u_cordic/mycordic/N505 ), .B(n788), .C(
        \u_cordic/mycordic/N522 ), .D(n1580), .Q(\u_cordic/mycordic/n467 ) );
  XNR21 U3927 ( .A(\u_cordic/mycordic/present_ANGLE_table[4][4] ), .B(
        \u_cordic/mycordic/sub_229/carry[4] ), .Q(\u_cordic/mycordic/N522 ) );
  XOR21 U3928 ( .A(\u_cordic/mycordic/present_ANGLE_table[4][4] ), .B(
        \u_cordic/mycordic/add_224/carry[4] ), .Q(\u_cordic/mycordic/N505 ) );
  INV3 U3929 ( .A(\u_cordic/mycordic/n449 ), .Q(n1183) );
  AOI221 U3930 ( .A(\u_cordic/mycordic/N538 ), .B(n785), .C(
        \u_cordic/mycordic/N554 ), .D(n1577), .Q(\u_cordic/mycordic/n449 ) );
  XOR21 U3931 ( .A(\u_cordic/mycordic/present_ANGLE_table[5][4] ), .B(
        \u_cordic/mycordic/add_233/carry [4]), .Q(\u_cordic/mycordic/N538 ) );
  XNR21 U3932 ( .A(\u_cordic/mycordic/present_ANGLE_table[5][4] ), .B(
        \u_cordic/mycordic/sub_236/carry [4]), .Q(\u_cordic/mycordic/N554 ) );
  INV3 U3933 ( .A(\u_cordic/mycordic/n448 ), .Q(n1184) );
  AOI221 U3934 ( .A(\u_cordic/mycordic/N539 ), .B(n785), .C(
        \u_cordic/mycordic/N555 ), .D(n1577), .Q(\u_cordic/mycordic/n448 ) );
  XOR21 U3935 ( .A(\u_cordic/mycordic/present_ANGLE_table[5][5] ), .B(
        \u_cordic/mycordic/add_233/carry [5]), .Q(\u_cordic/mycordic/N539 ) );
  XNR21 U3936 ( .A(\u_cordic/mycordic/present_ANGLE_table[5][5] ), .B(
        \u_cordic/mycordic/sub_236/carry [5]), .Q(\u_cordic/mycordic/N555 ) );
  INV3 U3937 ( .A(\u_cordic/mycordic/n392 ), .Q(n1173) );
  AOI221 U3938 ( .A(\u_cordic/mycordic/present_I_table[0][6] ), .B(n784), .C(
        \u_cordic/mycordic/N238 ), .D(n1575), .Q(\u_cordic/mycordic/n392 ) );
  XOR21 U3939 ( .A(\u_cordic/mycordic/sub_add_150_b0/carry [6]), .B(n44), .Q(
        \u_cordic/mycordic/N238 ) );
  BUF2 U3940 ( .A(\u_inFIFO/N34 ), .Q(n965) );
  BUF2 U3941 ( .A(\u_outFIFO/N36 ), .Q(n943) );
  INV3 U3942 ( .A(\u_decoder/fir_filter/n1037 ), .Q(n2200) );
  NAND22 U3943 ( .A(\u_decoder/fir_filter/I_data_mult_6_buff [0]), .B(n919), 
        .Q(\u_decoder/fir_filter/n1037 ) );
  INV3 U3944 ( .A(\u_decoder/fir_filter/n805 ), .Q(n2081) );
  NAND22 U3945 ( .A(\u_decoder/fir_filter/Q_data_mult_2_buff [0]), .B(n917), 
        .Q(\u_decoder/fir_filter/n805 ) );
  INV3 U3946 ( .A(\u_decoder/fir_filter/n740 ), .Q(n2080) );
  NAND22 U3947 ( .A(\u_decoder/fir_filter/Q_data_mult_6_buff [0]), .B(n919), 
        .Q(\u_decoder/fir_filter/n740 ) );
  INV3 U3948 ( .A(\u_decoder/fir_filter/n1102 ), .Q(n2201) );
  NAND22 U3949 ( .A(\u_decoder/fir_filter/I_data_mult_2_buff [0]), .B(n923), 
        .Q(\u_decoder/fir_filter/n1102 ) );
  INV3 U3950 ( .A(\u_decoder/iq_demod/cossin_dig/n38 ), .Q(n1505) );
  NAND22 U3951 ( .A(\u_decoder/iq_demod/cossin_dig/n39 ), .B(
        \u_decoder/iq_demod/cossin_dig/val_counter [2]), .Q(
        \u_decoder/iq_demod/cossin_dig/n38 ) );
  NOR31 U3952 ( .A(\u_inFIFO/n77 ), .B(\u_inFIFO/n76 ), .C(\u_inFIFO/n241 ), 
        .Q(\u_inFIFO/n233 ) );
  AOI211 U3953 ( .A(\u_decoder/iq_demod/cossin_dig/val_counter [1]), .B(
        \u_decoder/iq_demod/cossin_dig/N55 ), .C(
        \u_decoder/iq_demod/cossin_dig/val_counter [2]), .Q(
        \u_decoder/iq_demod/cossin_dig/n37 ) );
  NAND22 U3954 ( .A(\u_cordic/mycordic/present_I_table[0][7] ), .B(n970), .Q(
        \u_cordic/mycordic/n391 ) );
  NAND22 U3955 ( .A(\u_cordic/mycordic/present_Q_table[1][7] ), .B(n970), .Q(
        \u_cordic/mycordic/n537 ) );
  INV3 U3956 ( .A(\u_cordic/mycordic/n539 ), .Q(n1580) );
  NAND22 U3957 ( .A(\u_cordic/mycordic/present_Q_table[5][7] ), .B(n969), .Q(
        \u_cordic/mycordic/n539 ) );
  NAND31 U3958 ( .A(\u_cdr/div1/w_en_freq_synch ), .B(\u_cdr/w_sT ), .C(n976), 
        .Q(\u_cdr/div1/n26 ) );
  NOR21 U3959 ( .A(\u_decoder/fir_filter/n410 ), .B(
        \u_decoder/fir_filter/state [1]), .Q(\u_decoder/fir_filter/n1151 ) );
  NAND22 U3960 ( .A(\u_decoder/iq_demod/cossin_dig/counter [1]), .B(
        \u_decoder/iq_demod/cossin_dig/counter [0]), .Q(
        \u_decoder/iq_demod/cossin_dig/n43 ) );
  INV3 U3961 ( .A(\u_cordic/mycordic/n454 ), .Q(n1577) );
  NAND22 U3962 ( .A(\u_cordic/mycordic/present_Q_table[6][7] ), .B(n970), .Q(
        \u_cordic/mycordic/n454 ) );
  NOR40 U3963 ( .A(n2253), .B(n2620), .C(\u_cdr/phd1/cnt_phd/cnt [1]), .D(n984), .Q(\u_cdr/phd1/cnt_phd/N92 ) );
  INV3 U3964 ( .A(n2633), .Q(n2253) );
  NOR40 U3965 ( .A(\u_cdr/phd1/cnt_phd/cnt [2]), .B(
        \u_cdr/phd1/cnt_phd/cnt [3]), .C(\u_cdr/phd1/cnt_phd/cnt [4]), .D(
        \u_cdr/phd1/cnt_phd/cnt [5]), .Q(n2633) );
  NOR21 U3966 ( .A(n981), .B(\u_cordic/mycordic/present_Q_table[1][7] ), .Q(
        \u_cordic/mycordic/n345 ) );
  NOR40 U3967 ( .A(n984), .B(\u_inFIFO/n93 ), .C(\u_inFIFO/n94 ), .D(
        \u_inFIFO/n209 ), .Q(\u_inFIFO/N176 ) );
  XNR21 U3968 ( .A(\u_cdr/phd1/w_s4 ), .B(\u_cdr/phd1/w_s2 ), .Q(
        \u_cdr/phd1/n19 ) );
  XNR21 U3969 ( .A(\u_cdr/phd1/w_s2 ), .B(\u_cdr/phd1/w_s1 ), .Q(
        \u_cdr/phd1/n17 ) );
  AOI221 U3970 ( .A(sig_decod_outQ[3]), .B(n1689), .C(in_MUX_inSEL6[0]), .D(
        sig_coder_outSinQMasked[3]), .Q(n2686) );
  AOI221 U3971 ( .A(sig_decod_outQ[2]), .B(n1689), .C(in_MUX_inSEL6[0]), .D(
        sig_coder_outSinQMasked[2]), .Q(n2684) );
  AOI221 U3972 ( .A(sig_decod_outQ[1]), .B(n1689), .C(in_MUX_inSEL6[0]), .D(
        sig_coder_outSinQMasked[1]), .Q(n2682) );
  AOI221 U3973 ( .A(sig_decod_outQ[0]), .B(n1689), .C(in_MUX_inSEL6[0]), .D(
        sig_coder_outSinQMasked[0]), .Q(n2680) );
  AOI221 U3974 ( .A(sig_decod_outI[3]), .B(n1689), .C(in_MUX_inSEL6[0]), .D(
        sig_coder_outSinIMasked[3]), .Q(n2678) );
  AOI221 U3975 ( .A(sig_decod_outI[2]), .B(n1689), .C(in_MUX_inSEL6[0]), .D(
        sig_coder_outSinIMasked[2]), .Q(n2676) );
  AOI221 U3976 ( .A(sig_decod_outI[1]), .B(n1689), .C(in_MUX_inSEL6[0]), .D(
        sig_coder_outSinIMasked[1]), .Q(n2674) );
  AOI221 U3977 ( .A(sig_decod_outI[0]), .B(n1689), .C(in_MUX_inSEL6[0]), .D(
        sig_coder_outSinIMasked[0]), .Q(n2672) );
  AOI211 U3978 ( .A(\u_cordic/n35 ), .B(\u_cordic/n36 ), .C(n987), .Q(
        \u_cordic/N15 ) );
  OAI311 U3979 ( .A(n1663), .B(\u_cordic/n11 ), .C(\u_cordic/n12 ), .D(
        \u_cordic/n13 ), .Q(\u_cordic/n35 ) );
  NAND31 U3980 ( .A(\u_cordic/n12 ), .B(\u_cordic/n11 ), .C(n1663), .Q(
        \u_cordic/n36 ) );
  NAND22 U3981 ( .A(\u_outFIFO/n177 ), .B(\u_outFIFO/n176 ), .Q(
        \u_outFIFO/n534 ) );
  NOR21 U3982 ( .A(\u_inFIFO/currentState [0]), .B(\u_inFIFO/currentState [1]), 
        .Q(\u_inFIFO/n230 ) );
  NAND22 U3983 ( .A(\u_decoder/iq_demod/sin_out [0]), .B(n746), .Q(
        \u_decoder/iq_demod/cossin_dig/n32 ) );
  NOR21 U3984 ( .A(n981), .B(\u_cordic/mycordic/present_Q_table[5][7] ), .Q(
        \u_cordic/mycordic/n456 ) );
  NOR21 U3985 ( .A(\u_cdr/phd1/w_en_f ), .B(\u_cdr/phd1/w_en_d ), .Q(
        \u_cdr/phd1/n15 ) );
  AOI211 U3986 ( .A(\u_decoder/iq_demod/cossin_dig/n10 ), .B(
        \u_decoder/iq_demod/cossin_dig/n43 ), .C(
        \u_decoder/iq_demod/cossin_dig/n44 ), .Q(
        \u_decoder/iq_demod/cossin_dig/N42 ) );
  BUF2 U3987 ( .A(\u_cordic/mycordic/n108 ), .Q(n750) );
  INV3 U3988 ( .A(\u_cordic/mycordic/n393 ), .Q(n1172) );
  AOI221 U3989 ( .A(\u_cordic/mycordic/present_I_table[0][5] ), .B(n784), .C(
        \u_cordic/mycordic/N237 ), .D(n1575), .Q(\u_cordic/mycordic/n393 ) );
  XOR21 U3990 ( .A(\u_cordic/mycordic/sub_add_150_b0/carry [5]), .B(n45), .Q(
        \u_cordic/mycordic/N237 ) );
  NOR21 U3991 ( .A(\u_inFIFO/os1/sigQout2 ), .B(n293), .Q(
        \u_inFIFO/sig_fsm_start_R ) );
  NOR21 U3992 ( .A(n983), .B(\u_cordic/mycordic/present_Q_table[6][7] ), .Q(
        \u_cordic/mycordic/n438 ) );
  AOI211 U3993 ( .A(\u_cordic/n30 ), .B(\u_cordic/n31 ), .C(n982), .Q(
        \u_cordic/N17 ) );
  NAND22 U3994 ( .A(\u_cordic/present_state [2]), .B(\u_cordic/n12 ), .Q(
        \u_cordic/n30 ) );
  NAND31 U3995 ( .A(\u_cordic/present_state [0]), .B(\u_cordic/n11 ), .C(
        \u_cordic/present_state [1]), .Q(\u_cordic/n31 ) );
  NAND22 U3996 ( .A(\u_decoder/iq_demod/cossin_dig/n26 ), .B(n2249), .Q(
        \u_decoder/iq_demod/cossin_dig/n27 ) );
  INV3 U3997 ( .A(\u_decoder/iq_demod/cossin_dig/n55 ), .Q(n2249) );
  NAND22 U3998 ( .A(n753), .B(\u_decoder/iq_demod/n30 ), .Q(
        \u_decoder/iq_demod/n59 ) );
  BUF2 U3999 ( .A(\u_decoder/iq_demod/state [1]), .Q(n753) );
  NOR21 U4000 ( .A(\u_decoder/iq_demod/cossin_dig/n48 ), .B(
        \u_decoder/iq_demod/cossin_dig/n44 ), .Q(
        \u_decoder/iq_demod/cossin_dig/N21 ) );
  XNR21 U4001 ( .A(\u_decoder/iq_demod/cossin_dig/counter [1]), .B(
        \u_decoder/iq_demod/cossin_dig/counter [0]), .Q(
        \u_decoder/iq_demod/cossin_dig/n48 ) );
  AOI211 U4002 ( .A(\u_decoder/iq_demod/cossin_dig/state[0] ), .B(
        \u_decoder/iq_demod/cossin_dig/n45 ), .C(n987), .Q(
        \u_decoder/iq_demod/cossin_dig/N41 ) );
  NAND31 U4003 ( .A(\u_decoder/iq_demod/cossin_dig/n10 ), .B(
        \u_decoder/iq_demod/cossin_dig/n23 ), .C(
        \u_decoder/iq_demod/cossin_dig/n43 ), .Q(
        \u_decoder/iq_demod/cossin_dig/n45 ) );
  NAND22 U4004 ( .A(\u_decoder/iq_demod/cossin_dig/n27 ), .B(
        \u_decoder/iq_demod/cossin_dig/n29 ), .Q(
        \u_decoder/iq_demod/cossin_dig/n50 ) );
  NAND22 U4005 ( .A(\u_decoder/iq_demod/cos_out [2]), .B(n746), .Q(
        \u_decoder/iq_demod/cossin_dig/n29 ) );
  NAND22 U4006 ( .A(\u_decoder/iq_demod/cossin_dig/n27 ), .B(
        \u_decoder/iq_demod/cossin_dig/n28 ), .Q(
        \u_decoder/iq_demod/cossin_dig/n49 ) );
  NAND22 U4007 ( .A(\u_decoder/iq_demod/cos_out [1]), .B(n746), .Q(
        \u_decoder/iq_demod/cossin_dig/n28 ) );
  INV3 U4008 ( .A(\u_cdr/n28 ), .Q(n1586) );
  NAND22 U4009 ( .A(n1662), .B(n969), .Q(\u_cdr/n28 ) );
  INV3 U4010 ( .A(n2690), .Q(n1662) );
  AOI221 U4011 ( .A(\sig_MUX_inMUX14[0] ), .B(n1692), .C(in_MUX_inSEL11), .D(
        sig_DEMUX_outDEMUX2[3]), .Q(n2690) );
  INV3 U4012 ( .A(\u_cdr/dec1/n24 ), .Q(n1508) );
  OAI2111 U4013 ( .A(\u_cdr/cnt_d [0]), .B(\u_cdr/cnt_d [1]), .C(n978), .D(
        \u_cdr/dec1/n25 ), .Q(\u_cdr/dec1/n24 ) );
  INV3 U4014 ( .A(\u_decoder/iq_demod/cossin_dig/n25 ), .Q(n2243) );
  AOI221 U4015 ( .A(\u_decoder/iq_demod/cos_out [0]), .B(n746), .C(
        \u_decoder/iq_demod/cossin_dig/N55 ), .D(
        \u_decoder/iq_demod/cossin_dig/n26 ), .Q(
        \u_decoder/iq_demod/cossin_dig/n25 ) );
  INV3 U4016 ( .A(\u_decoder/iq_demod/cossin_dig/n30 ), .Q(n2244) );
  AOI221 U4017 ( .A(\u_decoder/iq_demod/cossin_dig/N52 ), .B(
        \u_decoder/iq_demod/cossin_dig/n26 ), .C(
        \u_decoder/iq_demod/cos_out [3]), .D(n746), .Q(
        \u_decoder/iq_demod/cossin_dig/n30 ) );
  INV3 U4018 ( .A(\u_cordic/mycordic/n358 ), .Q(n1174) );
  AOI221 U4019 ( .A(n1575), .B(\u_cordic/mycordic/present_Q_table[0][3] ), .C(
        n784), .D(\u_cordic/mycordic/present_Q_table[0][3] ), .Q(
        \u_cordic/mycordic/n358 ) );
  INV3 U4020 ( .A(\u_cordic/mycordic/n395 ), .Q(n1170) );
  AOI221 U4021 ( .A(\u_cordic/mycordic/present_I_table[0][3] ), .B(n784), .C(
        \u_cordic/mycordic/present_I_table[0][3] ), .D(n1575), .Q(
        \u_cordic/mycordic/n395 ) );
  INV3 U4022 ( .A(\u_cordic/mycordic/n547 ), .Q(n1255) );
  AOI221 U4023 ( .A(\u_cordic/mycordic/N448 ), .B(n835), .C(
        \u_cordic/mycordic/N476 ), .D(n1581), .Q(\u_cordic/mycordic/n547 ) );
  XOR21 U4024 ( .A(\u_cordic/mycordic/present_Q_table[4][0] ), .B(
        \u_cordic/mycordic/present_I_table[4][3] ), .Q(
        \u_cordic/mycordic/N476 ) );
  XNR21 U4025 ( .A(\u_cordic/mycordic/present_Q_table[4][0] ), .B(n155), .Q(
        \u_cordic/mycordic/N448 ) );
  INV3 U4026 ( .A(\u_cordic/mycordic/n487 ), .Q(n1263) );
  AOI221 U4027 ( .A(n299), .B(n835), .C(n299), .D(n1581), .Q(
        \u_cordic/mycordic/n487 ) );
  INV3 U4028 ( .A(\u_cordic/mycordic/n486 ), .Q(n1264) );
  AOI221 U4029 ( .A(\u_cordic/mycordic/N457 ), .B(n835), .C(
        \u_cordic/mycordic/N485 ), .D(n1581), .Q(\u_cordic/mycordic/n486 ) );
  XOR21 U4030 ( .A(\u_cordic/mycordic/present_ANGLE_table[3][1] ), .B(
        \u_cordic/mycordic/present_ANGLE_table[3][0] ), .Q(
        \u_cordic/mycordic/N485 ) );
  XNR21 U4031 ( .A(\u_cordic/mycordic/present_ANGLE_table[3][1] ), .B(
        \u_cordic/mycordic/present_ANGLE_table[3][0] ), .Q(
        \u_cordic/mycordic/N457 ) );
  INV3 U4032 ( .A(\u_cordic/mycordic/n485 ), .Q(n1265) );
  AOI221 U4033 ( .A(\u_cordic/mycordic/N458 ), .B(n835), .C(
        \u_cordic/mycordic/N486 ), .D(n1581), .Q(\u_cordic/mycordic/n485 ) );
  XOR21 U4034 ( .A(\u_cordic/mycordic/present_ANGLE_table[3][2] ), .B(
        \u_cordic/mycordic/sub_218/carry[2] ), .Q(\u_cordic/mycordic/N486 ) );
  XNR21 U4035 ( .A(\u_cordic/mycordic/present_ANGLE_table[3][2] ), .B(
        \u_cordic/mycordic/add_213/carry[2] ), .Q(\u_cordic/mycordic/N458 ) );
  INV3 U4036 ( .A(\u_cordic/mycordic/n469 ), .Q(n1241) );
  AOI221 U4037 ( .A(\u_cordic/mycordic/N503 ), .B(n788), .C(
        \u_cordic/mycordic/N520 ), .D(n1580), .Q(\u_cordic/mycordic/n469 ) );
  XNR21 U4038 ( .A(\u_cordic/mycordic/present_ANGLE_table[4][2] ), .B(
        \u_cordic/mycordic/sub_229/carry[2] ), .Q(\u_cordic/mycordic/N520 ) );
  XOR21 U4039 ( .A(\u_cordic/mycordic/present_ANGLE_table[4][2] ), .B(
        \u_cordic/mycordic/add_224/carry[2] ), .Q(\u_cordic/mycordic/N503 ) );
  INV3 U4040 ( .A(\u_cordic/mycordic/n451 ), .Q(n1181) );
  AOI221 U4041 ( .A(\u_cordic/mycordic/N536 ), .B(n785), .C(
        \u_cordic/mycordic/N552 ), .D(n1577), .Q(\u_cordic/mycordic/n451 ) );
  XOR21 U4042 ( .A(\u_cordic/mycordic/present_ANGLE_table[5][2] ), .B(
        \u_cordic/mycordic/present_ANGLE_table[5][1] ), .Q(
        \u_cordic/mycordic/N536 ) );
  XNR21 U4043 ( .A(\u_cordic/mycordic/present_ANGLE_table[5][2] ), .B(
        \u_cordic/mycordic/present_ANGLE_table[5][1] ), .Q(
        \u_cordic/mycordic/N552 ) );
  INV3 U4044 ( .A(\u_cordic/mycordic/n450 ), .Q(n1182) );
  AOI221 U4045 ( .A(\u_cordic/mycordic/N537 ), .B(n785), .C(
        \u_cordic/mycordic/N553 ), .D(n1577), .Q(\u_cordic/mycordic/n450 ) );
  XOR21 U4046 ( .A(\u_cordic/mycordic/present_ANGLE_table[5][3] ), .B(
        \u_cordic/mycordic/add_233/carry [3]), .Q(\u_cordic/mycordic/N537 ) );
  XNR21 U4047 ( .A(\u_cordic/mycordic/present_ANGLE_table[5][3] ), .B(
        \u_cordic/mycordic/sub_236/carry [3]), .Q(\u_cordic/mycordic/N553 ) );
  INV3 U4048 ( .A(\u_cordic/mycordic/n394 ), .Q(n1171) );
  AOI221 U4049 ( .A(\u_cordic/mycordic/present_I_table[0][4] ), .B(n784), .C(
        \u_cordic/mycordic/N236 ), .D(n1575), .Q(\u_cordic/mycordic/n394 ) );
  XOR21 U4050 ( .A(n257), .B(n46), .Q(\u_cordic/mycordic/N236 ) );
  INV3 U4051 ( .A(\u_cordic/mycordic/n357 ), .Q(n1175) );
  AOI221 U4052 ( .A(n1575), .B(\u_cordic/mycordic/N244 ), .C(n784), .D(
        \u_cordic/mycordic/present_Q_table[0][4] ), .Q(
        \u_cordic/mycordic/n357 ) );
  XOR21 U4053 ( .A(n254), .B(n43), .Q(\u_cordic/mycordic/N244 ) );
  INV3 U4054 ( .A(\u_cordic/mycordic/n356 ), .Q(n1176) );
  AOI221 U4055 ( .A(n1575), .B(\u_cordic/mycordic/N245 ), .C(n784), .D(
        \u_cordic/mycordic/present_Q_table[0][5] ), .Q(
        \u_cordic/mycordic/n356 ) );
  XOR21 U4056 ( .A(\u_cordic/mycordic/sub_add_151_b0/carry [5]), .B(n42), .Q(
        \u_cordic/mycordic/N245 ) );
  INV3 U4057 ( .A(\u_decoder/iq_demod/n58 ), .Q(n1942) );
  AOI311 U4058 ( .A(n752), .B(\u_decoder/iq_demod/n59 ), .C(
        \u_decoder/sample_ready ), .D(n790), .Q(\u_decoder/iq_demod/n58 ) );
  INV3 U4059 ( .A(\u_cordic/mycordic/n470 ), .Q(n1240) );
  AOI221 U4060 ( .A(\u_cordic/mycordic/N502 ), .B(n788), .C(
        \u_cordic/mycordic/N519 ), .D(n1580), .Q(\u_cordic/mycordic/n470 ) );
  XOR21 U4061 ( .A(\u_cordic/mycordic/present_ANGLE_table[4][1] ), .B(
        \u_cordic/mycordic/present_ANGLE_table[4][0] ), .Q(
        \u_cordic/mycordic/N519 ) );
  XNR21 U4062 ( .A(\u_cordic/mycordic/present_ANGLE_table[4][1] ), .B(
        \u_cordic/mycordic/present_ANGLE_table[4][0] ), .Q(
        \u_cordic/mycordic/N502 ) );
  INV3 U4063 ( .A(\u_cordic/mycordic/n453 ), .Q(n1179) );
  AOI221 U4064 ( .A(\u_cordic/mycordic/N550 ), .B(n785), .C(
        \u_cordic/mycordic/N550 ), .D(n1577), .Q(\u_cordic/mycordic/n453 ) );
  INV3 U4065 ( .A(\u_cordic/mycordic/n471 ), .Q(n1239) );
  AOI221 U4066 ( .A(n300), .B(n788), .C(n300), .D(n1580), .Q(
        \u_cordic/mycordic/n471 ) );
  INV3 U4067 ( .A(\u_cordic/mycordic/n452 ), .Q(n1180) );
  AOI221 U4068 ( .A(n301), .B(n785), .C(n301), .D(n1577), .Q(
        \u_cordic/mycordic/n452 ) );
  INV3 U4069 ( .A(n2617), .Q(n1487) );
  NAND22 U4070 ( .A(n977), .B(n2250), .Q(n2617) );
  INV3 U4071 ( .A(\u_cdr/phd1/n13 ), .Q(n2250) );
  AOI221 U4072 ( .A(\u_cdr/phd1/w_en_f ), .B(\u_cdr/phd1/w_s1 ), .C(n302), .D(
        \u_cdr/phd1/w_s2 ), .Q(\u_cdr/phd1/n13 ) );
  INV3 U4073 ( .A(n2618), .Q(n1488) );
  NAND22 U4074 ( .A(n977), .B(n1779), .Q(n2618) );
  INV3 U4075 ( .A(\u_cdr/phd1/n12 ), .Q(n1779) );
  AOI221 U4076 ( .A(n313), .B(\u_cdr/phd1/w_s3 ), .C(\u_cdr/dir ), .D(
        \u_cdr/phd1/w_en_m ), .Q(\u_cdr/phd1/n12 ) );
  INV3 U4077 ( .A(n2619), .Q(n1489) );
  NAND22 U4078 ( .A(n977), .B(n2251), .Q(n2619) );
  INV3 U4079 ( .A(\u_cdr/phd1/n11 ), .Q(n2251) );
  AOI221 U4080 ( .A(\u_cdr/phd1/w_en_f ), .B(\u_cdr/phd1/w_s3 ), .C(n302), .D(
        \u_cdr/phd1/w_s4 ), .Q(\u_cdr/phd1/n11 ) );
  INV3 U4081 ( .A(\u_cdr/phd1/f1/n2 ), .Q(n1502) );
  NAND22 U4082 ( .A(n976), .B(n1780), .Q(\u_cdr/phd1/f1/n2 ) );
  INV3 U4083 ( .A(\u_cdr/phd1/n14 ), .Q(n1780) );
  AOI221 U4084 ( .A(n2252), .B(\u_cdr/dir ), .C(\u_cdr/phd1/w_s1 ), .D(
        \u_cdr/phd1/n15 ), .Q(\u_cdr/phd1/n14 ) );
  INV3 U4085 ( .A(\u_inFIFO/os1/dff1/n2 ), .Q(n1507) );
  NAND22 U4086 ( .A(n976), .B(n1658), .Q(\u_inFIFO/os1/dff1/n2 ) );
  INV3 U4087 ( .A(\u_mux3/n3 ), .Q(n1658) );
  AOI221 U4088 ( .A(\sig_MUX_inMUX3[0] ), .B(n1687), .C(in_MUX_inSEL3), .D(
        sig_DEMUX_outDEMUX1[2]), .Q(\u_mux3/n3 ) );
  INV3 U4089 ( .A(\u_cordic/my_rotation/n84 ), .Q(n1528) );
  NAND22 U4090 ( .A(\u_cordic/my_rotation/next_delta [0]), .B(n974), .Q(
        \u_cordic/my_rotation/n84 ) );
  XNR21 U4091 ( .A(\u_cordic/my_rotation/present_angle[0][0] ), .B(n61), .Q(
        \u_cordic/my_rotation/next_delta [0]) );
  NAND22 U4092 ( .A(n976), .B(n312), .Q(\u_cdr/phd1/n16 ) );
  NOR31 U4093 ( .A(n314), .B(\u_decoder/fir_filter/state [1]), .C(n985), .Q(
        \u_decoder/fir_filter/N12 ) );
  AOI211 U4094 ( .A(n315), .B(n1089), .C(n987), .Q(n1490) );
  NOR21 U4095 ( .A(\u_decoder/iq_demod/state [0]), .B(\u_decoder/iq_demod/n69 ), .Q(\u_decoder/iq_demod/N13 ) );
  NOR21 U4096 ( .A(n980), .B(\u_coder/n148 ), .Q(\u_coder/N501 ) );
  NOR21 U4097 ( .A(n981), .B(\u_coder/n147 ), .Q(\u_coder/N499 ) );
  INV3 U4098 ( .A(\u_decoder/iq_demod/n68 ), .Q(n1315) );
  AOI221 U4099 ( .A(\u_decoder/iq_demod/I_if_buff[3] ), .B(
        \u_decoder/iq_demod/n61 ), .C(n1584), .D(sig_DEMUX_outDEMUX18[3]), .Q(
        \u_decoder/iq_demod/n68 ) );
  NOR21 U4100 ( .A(in_DEMUX_inSEL17), .B(n1674), .Q(sig_DEMUX_outDEMUX18[3])
         );
  INV3 U4101 ( .A(\u_decoder/iq_demod/n64 ), .Q(n1319) );
  AOI221 U4102 ( .A(\u_decoder/iq_demod/Q_if_buff[3] ), .B(
        \u_decoder/iq_demod/n61 ), .C(n1584), .D(sig_DEMUX_outDEMUX17[3]), .Q(
        \u_decoder/iq_demod/n64 ) );
  NOR21 U4103 ( .A(in_DEMUX_inSEL17), .B(n1666), .Q(sig_DEMUX_outDEMUX17[3])
         );
  INV3 U4104 ( .A(\u_decoder/iq_demod/n67 ), .Q(n1316) );
  AOI221 U4105 ( .A(sig_DEMUX_outDEMUX18[2]), .B(n1584), .C(
        \u_decoder/iq_demod/I_if_signed [2]), .D(\u_decoder/iq_demod/n61 ), 
        .Q(\u_decoder/iq_demod/n67 ) );
  NOR21 U4106 ( .A(in_DEMUX_inSEL17), .B(n1676), .Q(sig_DEMUX_outDEMUX18[2])
         );
  INV3 U4107 ( .A(\u_decoder/iq_demod/n66 ), .Q(n1317) );
  AOI221 U4108 ( .A(sig_DEMUX_outDEMUX18[1]), .B(n1584), .C(
        \u_decoder/iq_demod/I_if_signed [1]), .D(\u_decoder/iq_demod/n61 ), 
        .Q(\u_decoder/iq_demod/n66 ) );
  NOR21 U4109 ( .A(in_DEMUX_inSEL17), .B(n1678), .Q(sig_DEMUX_outDEMUX18[1])
         );
  INV3 U4110 ( .A(\u_decoder/iq_demod/n65 ), .Q(n1318) );
  AOI221 U4111 ( .A(sig_DEMUX_outDEMUX18[0]), .B(n1584), .C(
        \u_decoder/iq_demod/I_if_signed [0]), .D(\u_decoder/iq_demod/n61 ), 
        .Q(\u_decoder/iq_demod/n65 ) );
  NOR21 U4112 ( .A(in_DEMUX_inSEL17), .B(n1680), .Q(sig_DEMUX_outDEMUX18[0])
         );
  INV3 U4113 ( .A(\u_decoder/iq_demod/n63 ), .Q(n1320) );
  AOI221 U4114 ( .A(sig_DEMUX_outDEMUX17[2]), .B(n1584), .C(
        \u_decoder/iq_demod/Q_if_signed [2]), .D(\u_decoder/iq_demod/n61 ), 
        .Q(\u_decoder/iq_demod/n63 ) );
  NOR21 U4115 ( .A(in_DEMUX_inSEL17), .B(n1668), .Q(sig_DEMUX_outDEMUX17[2])
         );
  INV3 U4116 ( .A(\u_decoder/iq_demod/n62 ), .Q(n1321) );
  AOI221 U4117 ( .A(sig_DEMUX_outDEMUX17[1]), .B(n1584), .C(
        \u_decoder/iq_demod/Q_if_signed [1]), .D(\u_decoder/iq_demod/n61 ), 
        .Q(\u_decoder/iq_demod/n62 ) );
  NOR21 U4118 ( .A(in_DEMUX_inSEL17), .B(n1670), .Q(sig_DEMUX_outDEMUX17[1])
         );
  INV3 U4119 ( .A(\u_decoder/iq_demod/n60 ), .Q(n1322) );
  AOI221 U4120 ( .A(sig_DEMUX_outDEMUX17[0]), .B(n1584), .C(
        \u_decoder/iq_demod/Q_if_signed [0]), .D(\u_decoder/iq_demod/n61 ), 
        .Q(\u_decoder/iq_demod/n60 ) );
  NOR21 U4121 ( .A(in_DEMUX_inSEL17), .B(n1672), .Q(sig_DEMUX_outDEMUX17[0])
         );
  INV3 U4122 ( .A(n2644), .Q(n1495) );
  NAND22 U4123 ( .A(n977), .B(\u_inFIFO/os1/sigQout1 ), .Q(n2644) );
  INV3 U4124 ( .A(n2646), .Q(n1497) );
  NAND22 U4125 ( .A(n977), .B(\u_inFIFO/os2/sigQout1 ), .Q(n2646) );
  INV3 U4126 ( .A(n2648), .Q(n1499) );
  NAND22 U4127 ( .A(n977), .B(\u_outFIFO/os1/sigQout1 ), .Q(n2648) );
  INV3 U4128 ( .A(n2650), .Q(n1501) );
  NAND22 U4129 ( .A(n977), .B(\u_outFIFO/os2/sigQout1 ), .Q(n2650) );
  INV3 U4130 ( .A(\u_cordic/my_rotation/n65 ), .Q(n1509) );
  NAND22 U4131 ( .A(n976), .B(\u_cordic/cordic_to_rotation [3]), .Q(
        \u_cordic/my_rotation/n65 ) );
  INV3 U4132 ( .A(\u_cordic/my_rotation/n106 ), .Q(n1530) );
  NAND22 U4133 ( .A(\u_cordic/cordic_to_rotation [15]), .B(n974), .Q(
        \u_cordic/my_rotation/n106 ) );
  INV3 U4134 ( .A(\u_cordic/my_rotation/n107 ), .Q(n1531) );
  NAND22 U4135 ( .A(\u_cordic/cordic_to_rotation [14]), .B(n974), .Q(
        \u_cordic/my_rotation/n107 ) );
  INV3 U4136 ( .A(\u_cordic/my_rotation/n108 ), .Q(n1532) );
  NAND22 U4137 ( .A(\u_cordic/cordic_to_rotation [13]), .B(n973), .Q(
        \u_cordic/my_rotation/n108 ) );
  INV3 U4138 ( .A(\u_cordic/my_rotation/n109 ), .Q(n1533) );
  NAND22 U4139 ( .A(\u_cordic/cordic_to_rotation [12]), .B(n973), .Q(
        \u_cordic/my_rotation/n109 ) );
  INV3 U4140 ( .A(\u_cordic/my_rotation/n110 ), .Q(n1534) );
  NAND22 U4141 ( .A(\u_cordic/cordic_to_rotation [11]), .B(n973), .Q(
        \u_cordic/my_rotation/n110 ) );
  INV3 U4142 ( .A(\u_cordic/my_rotation/n111 ), .Q(n1535) );
  NAND22 U4143 ( .A(\u_cordic/cordic_to_rotation [10]), .B(n973), .Q(
        \u_cordic/my_rotation/n111 ) );
  INV3 U4144 ( .A(\u_cordic/my_rotation/n112 ), .Q(n1536) );
  NAND22 U4145 ( .A(\u_cordic/cordic_to_rotation [9]), .B(n973), .Q(
        \u_cordic/my_rotation/n112 ) );
  INV3 U4146 ( .A(\u_cordic/my_rotation/n113 ), .Q(n1537) );
  NAND22 U4147 ( .A(\u_cordic/cordic_to_rotation [8]), .B(n973), .Q(
        \u_cordic/my_rotation/n113 ) );
  INV3 U4148 ( .A(\u_cordic/my_rotation/n114 ), .Q(n1538) );
  NAND22 U4149 ( .A(\u_cordic/cordic_to_rotation [7]), .B(n973), .Q(
        \u_cordic/my_rotation/n114 ) );
  INV3 U4150 ( .A(\u_cordic/my_rotation/n115 ), .Q(n1539) );
  NAND22 U4151 ( .A(\u_cordic/cordic_to_rotation [6]), .B(n973), .Q(
        \u_cordic/my_rotation/n115 ) );
  INV3 U4152 ( .A(\u_cordic/my_rotation/n116 ), .Q(n1540) );
  NAND22 U4153 ( .A(\u_cordic/cordic_to_rotation [5]), .B(n974), .Q(
        \u_cordic/my_rotation/n116 ) );
  INV3 U4154 ( .A(\u_cordic/my_rotation/n117 ), .Q(n1541) );
  NAND22 U4155 ( .A(\u_cordic/cordic_to_rotation [4]), .B(n973), .Q(
        \u_cordic/my_rotation/n117 ) );
  INV3 U4156 ( .A(\u_cordic/my_rotation/n66 ), .Q(n1510) );
  NAND22 U4157 ( .A(\u_cordic/cordic_to_rotation [2]), .B(n975), .Q(
        \u_cordic/my_rotation/n66 ) );
  INV3 U4158 ( .A(\u_cordic/my_rotation/n67 ), .Q(n1511) );
  NAND22 U4159 ( .A(\u_cordic/cordic_to_rotation [1]), .B(n975), .Q(
        \u_cordic/my_rotation/n67 ) );
  INV3 U4160 ( .A(\u_cordic/my_rotation/n68 ), .Q(n1512) );
  NAND22 U4161 ( .A(\u_cordic/cordic_to_rotation [0]), .B(n975), .Q(
        \u_cordic/my_rotation/n68 ) );
  INV3 U4162 ( .A(\u_cordic/mycordic/n429 ), .Q(n1572) );
  NAND22 U4163 ( .A(\u_cordic/mycordic/present_C_table[1][2] ), .B(n970), .Q(
        \u_cordic/mycordic/n429 ) );
  INV3 U4164 ( .A(\u_cordic/mycordic/n426 ), .Q(n1569) );
  NAND22 U4165 ( .A(\u_cordic/mycordic/present_C_table[2][2] ), .B(n970), .Q(
        \u_cordic/mycordic/n426 ) );
  INV3 U4166 ( .A(\u_cordic/mycordic/n422 ), .Q(n1565) );
  NAND22 U4167 ( .A(\u_cordic/mycordic/present_C_table[3][2] ), .B(n971), .Q(
        \u_cordic/mycordic/n422 ) );
  INV3 U4168 ( .A(\u_cordic/mycordic/n419 ), .Q(n1562) );
  NAND22 U4169 ( .A(\u_cordic/mycordic/present_C_table[4][2] ), .B(n971), .Q(
        \u_cordic/mycordic/n419 ) );
  INV3 U4170 ( .A(\u_cordic/mycordic/n416 ), .Q(n1559) );
  NAND22 U4171 ( .A(\u_cordic/mycordic/present_C_table[5][2] ), .B(n971), .Q(
        \u_cordic/mycordic/n416 ) );
  INV3 U4172 ( .A(\u_cordic/mycordic/n412 ), .Q(n1555) );
  NAND22 U4173 ( .A(\u_cordic/mycordic/present_C_table[6][2] ), .B(n972), .Q(
        \u_cordic/mycordic/n412 ) );
  INV3 U4174 ( .A(\u_cordic/mycordic/n430 ), .Q(n1573) );
  NAND22 U4175 ( .A(\u_cordic/mycordic/present_C_table[1][1] ), .B(n970), .Q(
        \u_cordic/mycordic/n430 ) );
  INV3 U4176 ( .A(\u_cordic/mycordic/n427 ), .Q(n1570) );
  NAND22 U4177 ( .A(\u_cordic/mycordic/present_C_table[2][1] ), .B(n970), .Q(
        \u_cordic/mycordic/n427 ) );
  INV3 U4178 ( .A(\u_cordic/mycordic/n423 ), .Q(n1566) );
  NAND22 U4179 ( .A(\u_cordic/mycordic/present_C_table[3][1] ), .B(n971), .Q(
        \u_cordic/mycordic/n423 ) );
  INV3 U4180 ( .A(\u_cordic/mycordic/n420 ), .Q(n1563) );
  NAND22 U4181 ( .A(\u_cordic/mycordic/present_C_table[4][1] ), .B(n971), .Q(
        \u_cordic/mycordic/n420 ) );
  INV3 U4182 ( .A(\u_cordic/mycordic/n417 ), .Q(n1560) );
  NAND22 U4183 ( .A(\u_cordic/mycordic/present_C_table[5][1] ), .B(n971), .Q(
        \u_cordic/mycordic/n417 ) );
  INV3 U4184 ( .A(\u_cordic/mycordic/n414 ), .Q(n1557) );
  NAND22 U4185 ( .A(\u_cordic/mycordic/present_C_table[6][1] ), .B(n971), .Q(
        \u_cordic/mycordic/n414 ) );
  INV3 U4186 ( .A(\u_cordic/mycordic/n431 ), .Q(n1574) );
  NAND22 U4187 ( .A(\u_cordic/mycordic/present_C_table[1][0] ), .B(n970), .Q(
        \u_cordic/mycordic/n431 ) );
  INV3 U4188 ( .A(\u_cordic/mycordic/n428 ), .Q(n1571) );
  NAND22 U4189 ( .A(\u_cordic/mycordic/present_C_table[2][0] ), .B(n970), .Q(
        \u_cordic/mycordic/n428 ) );
  INV3 U4190 ( .A(\u_cordic/mycordic/n425 ), .Q(n1568) );
  NAND22 U4191 ( .A(\u_cordic/mycordic/present_C_table[3][0] ), .B(n970), .Q(
        \u_cordic/mycordic/n425 ) );
  INV3 U4192 ( .A(\u_cordic/mycordic/n421 ), .Q(n1564) );
  NAND22 U4193 ( .A(\u_cordic/mycordic/present_C_table[4][0] ), .B(n971), .Q(
        \u_cordic/mycordic/n421 ) );
  INV3 U4194 ( .A(\u_cordic/mycordic/n418 ), .Q(n1561) );
  NAND22 U4195 ( .A(\u_cordic/mycordic/present_C_table[5][0] ), .B(n971), .Q(
        \u_cordic/mycordic/n418 ) );
  INV3 U4196 ( .A(\u_cordic/mycordic/n415 ), .Q(n1558) );
  NAND22 U4197 ( .A(\u_cordic/mycordic/present_C_table[6][0] ), .B(n971), .Q(
        \u_cordic/mycordic/n415 ) );
  INV3 U4198 ( .A(in_DEMUX_inSEL17), .Q(n1696) );
  INV6 U4199 ( .A(\u_inFIFO/n116 ), .Q(n1614) );
  NAND22 U4200 ( .A(in_inFIFO_inData[3]), .B(n969), .Q(\u_inFIFO/n116 ) );
  INV6 U4201 ( .A(\u_inFIFO/n115 ), .Q(n1613) );
  NAND22 U4202 ( .A(in_inFIFO_inData[2]), .B(n969), .Q(\u_inFIFO/n115 ) );
  INV6 U4203 ( .A(\u_inFIFO/n114 ), .Q(n1612) );
  NAND22 U4204 ( .A(in_inFIFO_inData[1]), .B(n969), .Q(\u_inFIFO/n114 ) );
  INV6 U4205 ( .A(\u_inFIFO/n113 ), .Q(n1611) );
  NAND22 U4206 ( .A(in_inFIFO_inData[0]), .B(n969), .Q(\u_inFIFO/n113 ) );
  NOR31 U4207 ( .A(\u_demux1/n5 ), .B(in_DEMUX_inSEL1[2]), .C(
        in_DEMUX_inSEL1[1]), .Q(sig_DEMUX_outDEMUX1[0]) );
  INV3 U4208 ( .A(in_MUX_inSEL9[0]), .Q(n1691) );
  INV3 U4209 ( .A(in_MUX_inSEL9[1]), .Q(n1690) );
  NAND22 U4210 ( .A(in_DEMUX_inDEMUX1), .B(n1683), .Q(\u_demux1/n5 ) );
  INV3 U4211 ( .A(in_DEMUX_inSEL1[0]), .Q(n1683) );
  NAND22 U4212 ( .A(in_DEMUX_inDEMUX2), .B(n1686), .Q(n2693) );
  INV3 U4213 ( .A(in_DEMUX_inSEL2[0]), .Q(n1686) );
  AOI221 U4214 ( .A(\sig_MUX_inMUX14[0] ), .B(n1695), .C(\sig_MUX_inMUX13[0] ), 
        .D(in_MUX_inSEL15[0]), .Q(n2651) );
  AOI221 U4215 ( .A(\sig_MUX_inMUX5[0] ), .B(n1695), .C(in_MUX_inSEL15[0]), 
        .D(\sig_MUX_inMUX8[0] ), .Q(n2652) );
  NAND22 U4216 ( .A(sig_decod_outQ[0]), .B(n1691), .Q(n2663) );
  AOI221 U4217 ( .A(sig_coder_outSinQ[0]), .B(n1691), .C(in_MUX_inSEL9[0]), 
        .D(sig_coder_outSinQMasked[0]), .Q(n2664) );
  NAND22 U4218 ( .A(sig_decod_outQ[1]), .B(n1691), .Q(n2665) );
  AOI221 U4219 ( .A(sig_coder_outSinQ[1]), .B(n1691), .C(in_MUX_inSEL9[0]), 
        .D(sig_coder_outSinQMasked[1]), .Q(n2666) );
  NAND22 U4220 ( .A(sig_decod_outQ[2]), .B(n1691), .Q(n2667) );
  AOI221 U4221 ( .A(sig_coder_outSinQ[2]), .B(n1691), .C(in_MUX_inSEL9[0]), 
        .D(sig_coder_outSinQMasked[2]), .Q(n2668) );
  NAND22 U4222 ( .A(sig_decod_outQ[3]), .B(n1691), .Q(n2669) );
  AOI221 U4223 ( .A(sig_coder_outSinQ[3]), .B(n1691), .C(in_MUX_inSEL9[0]), 
        .D(sig_coder_outSinQMasked[3]), .Q(n2670) );
  AOI221 U4224 ( .A(sig_decod_outI[0]), .B(n1691), .C(sig_outFIFO_outData[0]), 
        .D(in_MUX_inSEL9[0]), .Q(n2655) );
  AOI221 U4225 ( .A(sig_coder_outSinI[0]), .B(n1691), .C(in_MUX_inSEL9[0]), 
        .D(sig_coder_outSinIMasked[0]), .Q(n2656) );
  AOI221 U4226 ( .A(sig_decod_outI[1]), .B(n1691), .C(sig_outFIFO_outData[1]), 
        .D(in_MUX_inSEL9[0]), .Q(n2657) );
  AOI221 U4227 ( .A(sig_coder_outSinI[1]), .B(n1691), .C(in_MUX_inSEL9[0]), 
        .D(sig_coder_outSinIMasked[1]), .Q(n2658) );
  AOI221 U4228 ( .A(sig_decod_outI[2]), .B(n1691), .C(sig_outFIFO_outData[2]), 
        .D(in_MUX_inSEL9[0]), .Q(n2659) );
  AOI221 U4229 ( .A(sig_coder_outSinI[2]), .B(n1691), .C(in_MUX_inSEL9[0]), 
        .D(sig_coder_outSinIMasked[2]), .Q(n2660) );
  AOI221 U4230 ( .A(sig_decod_outI[3]), .B(n1691), .C(sig_outFIFO_outData[3]), 
        .D(in_MUX_inSEL9[0]), .Q(n2661) );
  AOI221 U4231 ( .A(sig_coder_outSinI[3]), .B(n1691), .C(in_MUX_inSEL9[0]), 
        .D(sig_coder_outSinIMasked[3]), .Q(n2662) );
  INV3 U4232 ( .A(inReset), .Q(n980) );
  AOI221 U4233 ( .A(\sig_MUX_inMUX4[0] ), .B(n1695), .C(in_MUX_inSEL15[0]), 
        .D(\sig_MUX_inMUX3[0] ), .Q(n2654) );
  AOI221 U4234 ( .A(n1695), .B(\sig_MUX_inMUX11[0] ), .C(in_MUX_inSEL15[0]), 
        .D(\sig_MUX_inMUX12[0] ), .Q(n2653) );
  NOR31 U4235 ( .A(n2693), .B(in_DEMUX_inSEL2[1]), .C(n1684), .Q(
        sig_DEMUX_outDEMUX2[4]) );
  INV3 U4236 ( .A(in_DEMUX_inSEL2[2]), .Q(n1684) );
  NOR31 U4237 ( .A(\u_demux1/n5 ), .B(in_DEMUX_inSEL1[2]), .C(n1682), .Q(
        sig_DEMUX_outDEMUX1[2]) );
  NOR31 U4238 ( .A(n1685), .B(in_DEMUX_inSEL2[2]), .C(n2692), .Q(
        sig_DEMUX_outDEMUX2[3]) );
  INV3 U4239 ( .A(inReset), .Q(n984) );
  INV3 U4240 ( .A(inReset), .Q(n983) );
  INV3 U4241 ( .A(inReset), .Q(n981) );
  INV3 U4242 ( .A(inReset), .Q(n982) );
  NAND22 U4243 ( .A(in_DEMUX_inSEL1[0]), .B(in_DEMUX_inDEMUX1), .Q(
        \u_demux1/n4 ) );
  NAND22 U4244 ( .A(in_DEMUX_inSEL2[0]), .B(in_DEMUX_inDEMUX2), .Q(n2692) );
  INV3 U4245 ( .A(inReset), .Q(n985) );
  INV3 U4246 ( .A(inReset), .Q(n986) );
  INV3 U4247 ( .A(in_MUX_inSEL15[0]), .Q(n1695) );
  INV3 U4248 ( .A(inReset), .Q(n987) );
  NOR31 U4249 ( .A(\u_demux1/n5 ), .B(in_DEMUX_inSEL1[1]), .C(n1681), .Q(
        sig_DEMUX_outDEMUX1[4]) );
  INV3 U4250 ( .A(in_DEMUX_inSEL1[2]), .Q(n1681) );
  INV3 U4251 ( .A(in_MUX_inSEL6[1]), .Q(n1688) );
  INV3 U4252 ( .A(in_MUX_inSEL3), .Q(n1687) );
  INV3 U4253 ( .A(in_DEMUX_inDEMUX18[3]), .Q(n1674) );
  INV3 U4254 ( .A(in_DEMUX_inDEMUX18[2]), .Q(n1676) );
  INV3 U4255 ( .A(in_DEMUX_inDEMUX18[1]), .Q(n1678) );
  INV3 U4256 ( .A(in_DEMUX_inDEMUX18[0]), .Q(n1680) );
  INV3 U4257 ( .A(in_DEMUX_inDEMUX17[3]), .Q(n1666) );
  INV3 U4258 ( .A(in_DEMUX_inDEMUX17[2]), .Q(n1668) );
  INV3 U4259 ( .A(in_DEMUX_inDEMUX17[1]), .Q(n1670) );
  INV3 U4260 ( .A(in_DEMUX_inDEMUX17[0]), .Q(n1672) );
  INV3 U4261 ( .A(in_DEMUX_inSEL1[1]), .Q(n1682) );
  INV3 U4262 ( .A(in_DEMUX_inSEL2[1]), .Q(n1685) );
  INV3 U4263 ( .A(in_MUX_inSEL11), .Q(n1692) );
  INV3 U4264 ( .A(in_MUX_inSEL12), .Q(n1693) );
  INV3 U4265 ( .A(in_MUX_inSEL15[1]), .Q(n1694) );
  INV3 U4266 ( .A(n2645), .Q(n1496) );
  NAND22 U4267 ( .A(n977), .B(sig_DEMUX_outDEMUX2[0]), .Q(n2645) );
  NOR31 U4268 ( .A(n2693), .B(in_DEMUX_inSEL2[2]), .C(in_DEMUX_inSEL2[1]), .Q(
        sig_DEMUX_outDEMUX2[0]) );
  INV3 U4269 ( .A(n2647), .Q(n1498) );
  NAND22 U4270 ( .A(n977), .B(in_outFIFO_inReadEnable), .Q(n2647) );
  NAND22 U4271 ( .A(\u_cdr/div1/N34 ), .B(\u_cdr/w_nb_P [1]), .Q(n1047) );
  CLKIN3 U4272 ( .A(n1047), .Q(n988) );
  NAND22 U4273 ( .A(n1003), .B(n1008), .Q(\u_cdr/div1/n31 ) );
  NAND22 U4274 ( .A(\u_cdr/div1/n31 ), .B(\u_cdr/div1/n10 ), .Q(n991) );
  OAI212 U4275 ( .A(\u_cdr/cnt_d [1]), .B(\u_cdr/cnt_d [0]), .C(n990), .Q(
        n1025) );
  OAI222 U4276 ( .A(\u_cdr/div1/n26 ), .B(n991), .C(\u_cdr/div1/n10 ), .D(
        n1025), .Q(\u_cdr/div1/n37 ) );
  NAND22 U4277 ( .A(\u_cdr/div1/n9 ), .B(\u_cdr/div1/n10 ), .Q(n1021) );
  CLKIN3 U4278 ( .A(n1021), .Q(n1026) );
  NAND22 U4279 ( .A(\u_cdr/div1/n9 ), .B(\u_cdr/div1/n8 ), .Q(n1067) );
  CLKIN3 U4280 ( .A(n1067), .Q(n1069) );
  NAND22 U4281 ( .A(n1069), .B(\u_cdr/div1/n10 ), .Q(n996) );
  OAI212 U4282 ( .A(n1026), .B(\u_cdr/div1/n8 ), .C(n996), .Q(n1108) );
  CLKIN3 U4283 ( .A(n1108), .Q(n995) );
  NAND22 U4284 ( .A(n1025), .B(\u_cdr/phd1/n9 ), .Q(n1016) );
  NAND22 U4285 ( .A(\u_cdr/div1/n30 ), .B(n1025), .Q(n1020) );
  CLKIN3 U4286 ( .A(n1025), .Q(n1017) );
  NAND22 U4287 ( .A(\u_cdr/w_nb_P [1]), .B(\u_cdr/w_nb_P [2]), .Q(n1051) );
  CLKIN3 U4288 ( .A(n1051), .Q(n997) );
  OAI212 U4289 ( .A(\u_cdr/phd1/n9 ), .B(n997), .C(n1025), .Q(n992) );
  CLKIN3 U4290 ( .A(n996), .Q(n1027) );
  NAND22 U4291 ( .A(n1027), .B(n124), .Q(n1006) );
  OAI212 U4292 ( .A(n1027), .B(n124), .C(n1006), .Q(n1110) );
  CLKIN3 U4293 ( .A(n1110), .Q(n1002) );
  NAND22 U4294 ( .A(n997), .B(\u_cdr/w_nb_P [3]), .Q(n998) );
  CLKIN3 U4295 ( .A(n998), .Q(n1012) );
  OAI212 U4296 ( .A(\u_cdr/phd1/n9 ), .B(n1012), .C(n1025), .Q(n999) );
  CLKIN3 U4297 ( .A(n1003), .Q(n1004) );
  CLKIN3 U4298 ( .A(\u_cdr/div1/n26 ), .Q(n1009) );
  NAND22 U4299 ( .A(n1004), .B(n1009), .Q(n1005) );
  CLKIN3 U4300 ( .A(n1005), .Q(n1023) );
  CLKIN3 U4301 ( .A(n1006), .Q(n1007) );
  NAND22 U4302 ( .A(n1007), .B(\u_cdr/div1/n7 ), .Q(n1116) );
  OAI212 U4303 ( .A(n1007), .B(\u_cdr/div1/n7 ), .C(n1116), .Q(n1111) );
  CLKIN3 U4304 ( .A(n1008), .Q(n1010) );
  NAND22 U4305 ( .A(n1010), .B(n1009), .Q(n1011) );
  CLKIN3 U4306 ( .A(n1011), .Q(n1022) );
  NAND22 U4307 ( .A(n1012), .B(\u_cdr/w_nb_P [4]), .Q(n1013) );
  XNR21 U4308 ( .A(n1013), .B(\u_cdr/w_nb_P [5]), .Q(n1014) );
  OAI212 U4309 ( .A(\u_cdr/div1/n7 ), .B(n1025), .C(n1015), .Q(
        \u_cdr/div1/n38 ) );
  CLKIN3 U4310 ( .A(n1016), .Q(n1018) );
  NAND22 U4311 ( .A(n1020), .B(n1019), .Q(\u_cdr/div1/n39 ) );
  NAND22 U4312 ( .A(n1051), .B(n1021), .Q(n1109) );
  OAI212 U4313 ( .A(\u_cdr/div1/n9 ), .B(n1025), .C(n1024), .Q(
        \u_cdr/div1/n36 ) );
  NAND22 U4314 ( .A(n1026), .B(n29), .Q(n1029) );
  CLKIN3 U4315 ( .A(n1029), .Q(n1028) );
  NAND22 U4316 ( .A(n1027), .B(n29), .Q(n1030) );
  OAI212 U4317 ( .A(n1028), .B(\u_cdr/div1/n8 ), .C(n1030), .Q(n1081) );
  XNR21 U4318 ( .A(n1081), .B(\u_cdr/div1/cnt_div/cnt [3]), .Q(n2599) );
  OAI2112 U4319 ( .A(\u_cdr/div1/n9 ), .B(n29), .C(n1029), .D(n1051), .Q(n1102) );
  XNR21 U4320 ( .A(n1102), .B(\u_cdr/div1/cnt_div/cnt [2]), .Q(n2598) );
  CLKIN3 U4321 ( .A(n1030), .Q(n1031) );
  NAND22 U4322 ( .A(n1031), .B(n124), .Q(n1032) );
  OAI212 U4323 ( .A(n1031), .B(n124), .C(n1032), .Q(n1091) );
  XNR21 U4324 ( .A(n1091), .B(\u_cdr/div1/cnt_div/cnt [4]), .Q(n2597) );
  CLKIN3 U4325 ( .A(n1032), .Q(n1033) );
  NAND22 U4326 ( .A(n1033), .B(\u_cdr/div1/n7 ), .Q(n1132) );
  CLKIN3 U4327 ( .A(n1132), .Q(n1087) );
  XNR21 U4328 ( .A(n197), .B(\u_cdr/div1/N34 ), .Q(n1118) );
  CLKIN3 U4329 ( .A(n1118), .Q(n1036) );
  OAI212 U4330 ( .A(\u_cdr/div1/N34 ), .B(\u_cdr/w_nb_P [1]), .C(n1047), .Q(
        n1121) );
  CLKIN3 U4331 ( .A(n1121), .Q(n1045) );
  XNR21 U4332 ( .A(\u_cdr/div1/cnt_div/cnt [1]), .B(n1045), .Q(n1035) );
  OAI212 U4333 ( .A(n1033), .B(\u_cdr/div1/n7 ), .C(n1132), .Q(n1097) );
  CLKIN3 U4334 ( .A(n1097), .Q(n1122) );
  XNR21 U4335 ( .A(\u_cdr/div1/cnt_div/cnt [5]), .B(n1122), .Q(n1034) );
  XNR21 U4336 ( .A(n1081), .B(\u_cdr/dec1/cnt_dec/cnt [3]), .Q(n2603) );
  XNR21 U4337 ( .A(n1102), .B(\u_cdr/dec1/cnt_dec/cnt [2]), .Q(n2602) );
  XNR21 U4338 ( .A(n1091), .B(\u_cdr/dec1/cnt_dec/cnt [4]), .Q(n2601) );
  XNR21 U4339 ( .A(n29), .B(n196), .Q(n1039) );
  XNR21 U4340 ( .A(\u_cdr/dec1/cnt_dec/cnt [1]), .B(n1045), .Q(n1038) );
  XNR21 U4341 ( .A(\u_cdr/dec1/cnt_dec/cnt [5]), .B(n1122), .Q(n1037) );
  CLKIN3 U4342 ( .A(n1081), .Q(n1125) );
  CLKIN3 U4343 ( .A(n1102), .Q(n1124) );
  CLKIN3 U4344 ( .A(n1042), .Q(n1041) );
  CLKIN3 U4345 ( .A(n1091), .Q(n1123) );
  OAI212 U4346 ( .A(n1042), .B(n1091), .C(n1097), .Q(n1040) );
  NAND22 U4347 ( .A(n1044), .B(n1040), .Q(\u_cdr/phd1/cnt_phd/N14 ) );
  XNR21 U4348 ( .A(n1123), .B(n1041), .Q(\u_cdr/phd1/cnt_phd/N13 ) );
  NAND22 U4349 ( .A(n1102), .B(n1081), .Q(n1090) );
  NAND22 U4350 ( .A(n1132), .B(n1044), .Q(n2240) );
  NAND22 U4351 ( .A(\u_cdr/phd1/cnt_phd/cnt [0]), .B(n1121), .Q(n2608) );
  XNR21 U4352 ( .A(n1124), .B(n1045), .Q(n1142) );
  NAND22 U4353 ( .A(n1045), .B(n2620), .Q(n1043) );
  CLKIN3 U4354 ( .A(n1043), .Q(n1141) );
  NAND22 U4355 ( .A(n1132), .B(n1044), .Q(n2239) );
  CLKIN3 U4356 ( .A(n1044), .Q(\u_cdr/phd1/cnt_phd/N41 ) );
  XNR21 U4357 ( .A(n1081), .B(\u_cdr/phd1/cnt_phd/cnt [3]), .Q(n2616) );
  XNR21 U4358 ( .A(n1102), .B(\u_cdr/phd1/cnt_phd/cnt [2]), .Q(n2615) );
  XNR21 U4359 ( .A(n1091), .B(\u_cdr/phd1/cnt_phd/cnt [4]), .Q(n2614) );
  XNR21 U4360 ( .A(n2620), .B(\u_cdr/div1/N34 ), .Q(n1062) );
  CLKIN3 U4361 ( .A(n1062), .Q(n1076) );
  XNR21 U4362 ( .A(\u_cdr/phd1/cnt_phd/cnt [5]), .B(n1122), .Q(n1046) );
  XNR21 U4363 ( .A(\u_cdr/phd1/cnt_phd/cnt [1]), .B(n1045), .Q(n1061) );
  CLKIN3 U4364 ( .A(\u_cdr/dec1/n33 ), .Q(n1161) );
  CLKIN3 U4365 ( .A(\u_cdr/dec1/n32 ), .Q(n1162) );
  CLKIN3 U4366 ( .A(\u_cdr/dec1/n26 ), .Q(n1166) );
  CLKIN3 U4367 ( .A(\u_cdr/dec1/n29 ), .Q(n1165) );
  CLKIN3 U4368 ( .A(\u_cdr/dec1/n30 ), .Q(n1164) );
  CLKIN3 U4369 ( .A(\u_cdr/dec1/n31 ), .Q(n1163) );
  NAND22 U4370 ( .A(n1047), .B(\u_cdr/div1/n9 ), .Q(n1050) );
  CLKIN3 U4371 ( .A(n1050), .Q(n1048) );
  NAND22 U4372 ( .A(n1048), .B(\u_cdr/div1/n8 ), .Q(n1053) );
  OAI212 U4373 ( .A(n1048), .B(\u_cdr/div1/n8 ), .C(n1053), .Q(n1049) );
  XNR21 U4374 ( .A(n1049), .B(\u_cdr/phd1/cnt_phd/cnt [3]), .Q(n1060) );
  OAI212 U4375 ( .A(n29), .B(n1051), .C(n1050), .Q(n1052) );
  XNR21 U4376 ( .A(n1052), .B(\u_cdr/phd1/cnt_phd/cnt [2]), .Q(n1059) );
  CLKIN3 U4377 ( .A(n1053), .Q(n1054) );
  NAND22 U4378 ( .A(n1054), .B(n124), .Q(n1063) );
  OAI212 U4379 ( .A(n1054), .B(n124), .C(n1063), .Q(n1055) );
  XNR21 U4380 ( .A(n1055), .B(\u_cdr/phd1/cnt_phd/cnt [4]), .Q(n1058) );
  NAND22 U4381 ( .A(\u_cdr/w_nb_P [5]), .B(n1063), .Q(n1056) );
  XNR21 U4382 ( .A(n271), .B(n1056), .Q(n1057) );
  NAND41 U4383 ( .A(n1060), .B(n1059), .C(n1058), .D(n1057), .Q(n1066) );
  CLKIN3 U4384 ( .A(n1061), .Q(n1065) );
  OAI212 U4385 ( .A(\u_cdr/w_nb_P [5]), .B(n1063), .C(n1062), .Q(n1064) );
  OAI212 U4386 ( .A(\u_cdr/div1/n8 ), .B(\u_cdr/div1/n9 ), .C(n1067), .Q(n1068) );
  XNR21 U4387 ( .A(n1068), .B(\u_cdr/phd1/cnt_phd/cnt [3]), .Q(n1075) );
  XNR21 U4388 ( .A(\u_cdr/div1/n9 ), .B(\u_cdr/phd1/cnt_phd/cnt [2]), .Q(n1074) );
  NAND22 U4389 ( .A(n1069), .B(n124), .Q(n1077) );
  OAI212 U4390 ( .A(n1069), .B(n124), .C(n1077), .Q(n1070) );
  XNR21 U4391 ( .A(n1070), .B(\u_cdr/phd1/cnt_phd/cnt [4]), .Q(n1073) );
  NAND22 U4392 ( .A(\u_cdr/w_nb_P [5]), .B(n1077), .Q(n1071) );
  XNR21 U4393 ( .A(n271), .B(n1071), .Q(n1072) );
  NAND41 U4394 ( .A(n1075), .B(n1074), .C(n1073), .D(n1072), .Q(n1080) );
  XNR21 U4395 ( .A(\u_cdr/div1/n10 ), .B(\u_cdr/phd1/cnt_phd/cnt [1]), .Q(
        n1079) );
  OAI212 U4396 ( .A(\u_cdr/w_nb_P [5]), .B(n1077), .C(n1076), .Q(n1078) );
  XNR21 U4397 ( .A(n1091), .B(\u_cdr/dec1/cnt_dec/cnt [3]), .Q(n1085) );
  XNR21 U4398 ( .A(n1081), .B(\u_cdr/dec1/cnt_dec/cnt [2]), .Q(n1084) );
  XNR21 U4399 ( .A(n1097), .B(\u_cdr/dec1/cnt_dec/cnt [4]), .Q(n1083) );
  XNR21 U4400 ( .A(n1121), .B(\u_cdr/dec1/cnt_dec/cnt [0]), .Q(n1082) );
  NAND41 U4401 ( .A(n1085), .B(n1084), .C(n1083), .D(n1082), .Q(n1088) );
  XNR21 U4402 ( .A(n1102), .B(n278), .Q(n1086) );
  NAND22 U4403 ( .A(\u_cdr/dec1/w_s_r ), .B(n40), .Q(n1089) );
  CLKIN3 U4404 ( .A(n1090), .Q(n1092) );
  XOR31 U4405 ( .A(\u_cdr/dec1/cnt_r [3]), .B(n1123), .C(n1092), .Q(n1096) );
  NAND22 U4406 ( .A(n1092), .B(n1091), .Q(n1093) );
  CLKIN3 U4407 ( .A(n1093), .Q(n1098) );
  XOR31 U4408 ( .A(\u_cdr/dec1/cnt_r [4]), .B(n1122), .C(n1098), .Q(n1095) );
  NAND22 U4409 ( .A(\u_cdr/cnt_d [1]), .B(\u_cdr/cnt_d [0]), .Q(n1135) );
  NAND41 U4410 ( .A(n1096), .B(n1095), .C(n1132), .D(n1094), .Q(n1106) );
  NAND22 U4411 ( .A(n1098), .B(n1097), .Q(n1099) );
  XNR21 U4412 ( .A(n304), .B(n1099), .Q(n1101) );
  XOR31 U4413 ( .A(\u_cdr/dec1/cnt_r [2]), .B(n1125), .C(n1102), .Q(n1100) );
  NAND22 U4414 ( .A(n1101), .B(n1100), .Q(n1105) );
  XNR21 U4415 ( .A(n1102), .B(\u_cdr/dec1/cnt_r [1]), .Q(n1104) );
  XNR21 U4416 ( .A(n1121), .B(n250), .Q(n1103) );
  NAND22 U4417 ( .A(sig_DEMUX_outDEMUX1[4]), .B(in_MUX_inSEL12), .Q(n1107) );
  OAI212 U4418 ( .A(n40), .B(in_MUX_inSEL12), .C(n1107), .Q(n1659) );
  XNR21 U4419 ( .A(n1108), .B(\u_cdr/div1/cnt_div/cnt [3]), .Q(n1115) );
  XNR21 U4420 ( .A(n1109), .B(\u_cdr/div1/cnt_div/cnt [2]), .Q(n1114) );
  XNR21 U4421 ( .A(n1110), .B(\u_cdr/div1/cnt_div/cnt [4]), .Q(n1113) );
  XNR21 U4422 ( .A(n1111), .B(\u_cdr/div1/cnt_div/cnt [5]), .Q(n1112) );
  NAND41 U4423 ( .A(n1115), .B(n1114), .C(n1113), .D(n1112), .Q(n1120) );
  CLKIN3 U4424 ( .A(n1116), .Q(n1119) );
  XNR21 U4425 ( .A(\u_cdr/div1/cnt_div/cnt [1]), .B(\u_cdr/w_nb_P [1]), .Q(
        n1117) );
  XNR21 U4426 ( .A(n1121), .B(\u_cdr/dec1/cnt_r [1]), .Q(n1133) );
  XNR21 U4427 ( .A(n250), .B(\u_cdr/div1/N34 ), .Q(n1131) );
  XNR21 U4428 ( .A(\u_cdr/dec1/cnt_r [5]), .B(n1122), .Q(n1129) );
  XNR21 U4429 ( .A(\u_cdr/dec1/cnt_r [4]), .B(n1123), .Q(n1128) );
  XNR21 U4430 ( .A(\u_cdr/dec1/cnt_r [2]), .B(n1124), .Q(n1127) );
  XNR21 U4431 ( .A(\u_cdr/dec1/cnt_r [3]), .B(n1125), .Q(n1126) );
  NAND41 U4432 ( .A(n1133), .B(n1132), .C(n1131), .D(n1130), .Q(n1136) );
  CLKIN3 U4433 ( .A(n1134), .Q(n1140) );
  CLKIN3 U4434 ( .A(n1135), .Q(n1137) );
  CLKIN3 U4435 ( .A(n1138), .Q(n1139) );
  OAI212 U4436 ( .A(\u_inFIFO/outReadCount[1] ), .B(n2257), .C(\u_inFIFO/n85 ), 
        .Q(n2256) );
  OAI212 U4437 ( .A(\u_inFIFO/outReadCount[4] ), .B(\u_inFIFO/n82 ), .C(n2261), 
        .Q(n2262) );
  OAI222 U4438 ( .A(\u_inFIFO/outReadCount[1] ), .B(n2263), .C(n2263), .D(
        \u_inFIFO/n85 ), .Q(n2264) );
  OAI212 U4439 ( .A(\u_outFIFO/outReadCount[1] ), .B(n2304), .C(
        \u_outFIFO/n183 ), .Q(n2303) );
  OAI212 U4440 ( .A(\u_outFIFO/outReadCount[4] ), .B(\u_outFIFO/n180 ), .C(
        n2308), .Q(n2309) );
  OAI222 U4441 ( .A(\u_outFIFO/outReadCount[1] ), .B(n2310), .C(n2310), .D(
        \u_outFIFO/n183 ), .Q(n2311) );
  XNR31 U4442 ( .A(\u_decoder/iq_demod/dp_cluster_1/mult_149/A2[5] ), .B(n1959), .C(n2316), .Q(\u_decoder/iq_demod/dp_cluster_1/mult_I_sin_out [7]) );
  OAI212 U4443 ( .A(\u_decoder/iq_demod/dp_cluster_1/mult_149/A1[4] ), .B(
        n2317), .C(\u_decoder/iq_demod/dp_cluster_1/mult_149/A2[4] ), .Q(n2318) );
  XOR31 U4444 ( .A(\u_decoder/iq_demod/dp_cluster_1/mult_149/A2[4] ), .B(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/A1[4] ), .C(n2317), .Q(
        \u_decoder/iq_demod/dp_cluster_1/mult_I_sin_out [6]) );
  XNR31 U4445 ( .A(\u_decoder/iq_demod/dp_cluster_1/mult_150/A2[5] ), .B(n1952), .C(n2323), .Q(\u_decoder/iq_demod/dp_cluster_1/mult_Q_cos_out [7]) );
  OAI212 U4446 ( .A(\u_decoder/iq_demod/dp_cluster_1/mult_150/A1[4] ), .B(
        n2324), .C(\u_decoder/iq_demod/dp_cluster_1/mult_150/A2[4] ), .Q(n2325) );
  XOR31 U4447 ( .A(\u_decoder/iq_demod/dp_cluster_1/mult_150/A2[4] ), .B(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/A1[4] ), .C(n2324), .Q(
        \u_decoder/iq_demod/dp_cluster_1/mult_Q_cos_out [6]) );
  XNR31 U4448 ( .A(\u_decoder/iq_demod/dp_cluster_0/mult_148/A2[5] ), .B(n1960), .C(n2330), .Q(\u_decoder/iq_demod/dp_cluster_0/mult_I_cos_out [7]) );
  OAI212 U4449 ( .A(\u_decoder/iq_demod/dp_cluster_0/mult_148/A1[4] ), .B(
        n2331), .C(\u_decoder/iq_demod/dp_cluster_0/mult_148/A2[4] ), .Q(n2332) );
  XOR31 U4450 ( .A(\u_decoder/iq_demod/dp_cluster_0/mult_148/A2[4] ), .B(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/A1[4] ), .C(n2331), .Q(
        \u_decoder/iq_demod/dp_cluster_0/mult_I_cos_out [6]) );
  OAI212 U4451 ( .A(\u_decoder/iq_demod/dp_cluster_0/mult_151/A1[4] ), .B(
        n2338), .C(\u_decoder/iq_demod/dp_cluster_0/mult_151/A2[4] ), .Q(n2339) );
  OAI212 U4452 ( .A(n2347), .B(n2348), .C(n2349), .Q(n2346) );
  OAI212 U4453 ( .A(\u_decoder/fir_filter/dp_cluster_0/r177/A2[6] ), .B(n2350), 
        .C(n2351), .Q(\u_decoder/fir_filter/Q_data_mult_0 [8]) );
  OAI212 U4454 ( .A(\u_decoder/fir_filter/dp_cluster_0/r177/PROD1[4] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r177/A1[3] ), .C(n2354), .Q(n2355)
         );
  OAI212 U4455 ( .A(n1939), .B(n2344), .C(
        \u_decoder/fir_filter/dp_cluster_0/r177/A2[9] ), .Q(n2357) );
  OAI212 U4456 ( .A(n2345), .B(n1931), .C(n2358), .Q(n2344) );
  OAI212 U4457 ( .A(\u_decoder/fir_filter/dp_cluster_0/r177/A1[8] ), .B(n1924), 
        .C(\u_decoder/fir_filter/dp_cluster_0/r177/A2[8] ), .Q(n2358) );
  OAI222 U4458 ( .A(\u_decoder/fir_filter/dp_cluster_0/r177/A1[6] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r177/A2[6] ), .C(
        \u_decoder/fir_filter/dp_cluster_0/r177/A1[7] ), .D(
        \u_decoder/fir_filter/dp_cluster_0/r177/A2[7] ), .Q(n2362) );
  OAI212 U4459 ( .A(\u_decoder/fir_filter/dp_cluster_0/r178/PROD1[5] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r178/A1[4] ), .C(n2368), .Q(n2370)
         );
  OAI212 U4460 ( .A(n1939), .B(n2372), .C(
        \u_decoder/fir_filter/dp_cluster_0/r178/A2[10] ), .Q(n2373) );
  OAI212 U4461 ( .A(n1873), .B(n1872), .C(n2374), .Q(n2372) );
  OAI212 U4462 ( .A(\u_decoder/fir_filter/dp_cluster_0/r178/A1[9] ), .B(n2363), 
        .C(\u_decoder/fir_filter/dp_cluster_0/r178/A2[9] ), .Q(n2374) );
  OAI212 U4463 ( .A(n2364), .B(n1874), .C(n2375), .Q(n2363) );
  OAI212 U4464 ( .A(\u_decoder/fir_filter/dp_cluster_0/r178/A1[8] ), .B(n1875), 
        .C(\u_decoder/fir_filter/dp_cluster_0/r178/A2[8] ), .Q(n2375) );
  OAI212 U4465 ( .A(\u_decoder/fir_filter/dp_cluster_0/r178/A1[7] ), .B(n2365), 
        .C(\u_decoder/fir_filter/dp_cluster_0/r178/A2[7] ), .Q(n2376) );
  OAI212 U4466 ( .A(n1880), .B(n1879), .C(n2383), .Q(n2382) );
  OAI212 U4467 ( .A(\u_decoder/fir_filter/dp_cluster_0/r179/CARRYB[7][3] ), 
        .B(n2378), .C(\u_decoder/fir_filter/dp_cluster_0/r179/A2[9] ), .Q(
        n2383) );
  OAI212 U4468 ( .A(n2379), .B(n1881), .C(n2384), .Q(n2378) );
  OAI212 U4469 ( .A(\u_decoder/fir_filter/dp_cluster_0/r179/A1[8] ), .B(n1882), 
        .C(\u_decoder/fir_filter/dp_cluster_0/r179/A2[8] ), .Q(n2384) );
  OAI212 U4470 ( .A(\u_decoder/fir_filter/dp_cluster_0/r179/A1[7] ), .B(n1885), 
        .C(\u_decoder/fir_filter/dp_cluster_0/r179/A2[7] ), .Q(n2385) );
  OAI212 U4471 ( .A(n2390), .B(n2391), .C(n2392), .Q(
        \u_decoder/fir_filter/Q_data_mult_3 [10]) );
  OAI222 U4472 ( .A(\u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[7][5] ), 
        .B(\u_decoder/fir_filter/dp_cluster_0/r180/A2[11] ), .C(
        \u_decoder/fir_filter/dp_cluster_0/r180/A1[8] ), .D(
        \u_decoder/fir_filter/dp_cluster_0/r180/A2[8] ), .Q(n2401) );
  OAI212 U4473 ( .A(\u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[7][5] ), 
        .B(n2397), .C(\u_decoder/fir_filter/dp_cluster_0/r180/A2[11] ), .Q(
        n2402) );
  OAI212 U4474 ( .A(n2400), .B(n1913), .C(n2403), .Q(n2397) );
  OAI212 U4475 ( .A(n2391), .B(n2399), .C(n2389), .Q(n2404) );
  OAI212 U4476 ( .A(n2400), .B(n2406), .C(n2403), .Q(n2405) );
  OAI212 U4477 ( .A(n2390), .B(n2408), .C(n2391), .Q(n2387) );
  IMAJ31 U4478 ( .A(\u_decoder/fir_filter/dp_cluster_0/r180/A2[7] ), .B(n2395), 
        .C(\u_decoder/fir_filter/dp_cluster_0/r180/A1[7] ), .Q(n2390) );
  OAI212 U4479 ( .A(n2412), .B(n2413), .C(n2414), .Q(
        \u_decoder/fir_filter/Q_data_mult_4 [10]) );
  XOR31 U4480 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_308/A1[7] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/A2[7] ), .C(n2417), .Q(
        \u_decoder/fir_filter/Q_data_mult_4 [9]) );
  OAI222 U4481 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[7][5] ), 
        .B(\u_decoder/fir_filter/dp_cluster_0/mult_308/A2[11] ), .C(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/A1[8] ), .D(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/A2[8] ), .Q(n2423) );
  OAI212 U4482 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[7][5] ), 
        .B(n2419), .C(\u_decoder/fir_filter/dp_cluster_0/mult_308/A2[11] ), 
        .Q(n2424) );
  OAI212 U4483 ( .A(n2422), .B(n1897), .C(n2425), .Q(n2419) );
  OAI212 U4484 ( .A(n2413), .B(n2421), .C(n2411), .Q(n2426) );
  XOR31 U4485 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_308/A2[11] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[7][5] ), .C(n2427), 
        .Q(\u_decoder/fir_filter/Q_data_mult_4 [13]) );
  OAI212 U4486 ( .A(n2422), .B(n2428), .C(n2425), .Q(n2427) );
  OAI212 U4487 ( .A(n2412), .B(n2430), .C(n2413), .Q(n2409) );
  IMAJ31 U4488 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_308/A2[7] ), .B(
        n2417), .C(\u_decoder/fir_filter/dp_cluster_0/mult_308/A1[7] ), .Q(
        n2412) );
  OAI212 U4489 ( .A(n2434), .B(n2435), .C(n2436), .Q(n2433) );
  OAI212 U4490 ( .A(\u_decoder/fir_filter/dp_cluster_0/r164/A2[6] ), .B(n2437), 
        .C(n2438), .Q(\u_decoder/fir_filter/I_data_mult_0 [8]) );
  OAI212 U4491 ( .A(\u_decoder/fir_filter/dp_cluster_0/r164/PROD1[4] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r164/A1[3] ), .C(n2441), .Q(n2442)
         );
  OAI212 U4492 ( .A(n1868), .B(n2431), .C(
        \u_decoder/fir_filter/dp_cluster_0/r164/A2[9] ), .Q(n2444) );
  OAI212 U4493 ( .A(n2432), .B(n1860), .C(n2445), .Q(n2431) );
  OAI212 U4494 ( .A(\u_decoder/fir_filter/dp_cluster_0/r164/A1[8] ), .B(n1853), 
        .C(\u_decoder/fir_filter/dp_cluster_0/r164/A2[8] ), .Q(n2445) );
  OAI222 U4495 ( .A(\u_decoder/fir_filter/dp_cluster_0/r164/A1[6] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r164/A2[6] ), .C(
        \u_decoder/fir_filter/dp_cluster_0/r164/A1[7] ), .D(
        \u_decoder/fir_filter/dp_cluster_0/r164/A2[7] ), .Q(n2449) );
  OAI212 U4496 ( .A(\u_decoder/fir_filter/dp_cluster_0/r165/PROD1[5] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r165/A1[4] ), .C(n2455), .Q(n2457)
         );
  OAI212 U4497 ( .A(n1868), .B(n2459), .C(
        \u_decoder/fir_filter/dp_cluster_0/r165/A2[10] ), .Q(n2460) );
  OAI212 U4498 ( .A(n1802), .B(n1801), .C(n2461), .Q(n2459) );
  OAI212 U4499 ( .A(\u_decoder/fir_filter/dp_cluster_0/r165/A1[9] ), .B(n2450), 
        .C(\u_decoder/fir_filter/dp_cluster_0/r165/A2[9] ), .Q(n2461) );
  OAI212 U4500 ( .A(n2451), .B(n1803), .C(n2462), .Q(n2450) );
  OAI212 U4501 ( .A(\u_decoder/fir_filter/dp_cluster_0/r165/A1[8] ), .B(n1804), 
        .C(\u_decoder/fir_filter/dp_cluster_0/r165/A2[8] ), .Q(n2462) );
  OAI212 U4502 ( .A(\u_decoder/fir_filter/dp_cluster_0/r165/A1[7] ), .B(n2452), 
        .C(\u_decoder/fir_filter/dp_cluster_0/r165/A2[7] ), .Q(n2463) );
  OAI212 U4503 ( .A(n1809), .B(n1808), .C(n2470), .Q(n2469) );
  OAI212 U4504 ( .A(\u_decoder/fir_filter/dp_cluster_0/r166/CARRYB[7][3] ), 
        .B(n2465), .C(\u_decoder/fir_filter/dp_cluster_0/r166/A2[9] ), .Q(
        n2470) );
  OAI212 U4505 ( .A(n2466), .B(n1810), .C(n2471), .Q(n2465) );
  OAI212 U4506 ( .A(\u_decoder/fir_filter/dp_cluster_0/r166/A1[8] ), .B(n1811), 
        .C(\u_decoder/fir_filter/dp_cluster_0/r166/A2[8] ), .Q(n2471) );
  OAI212 U4507 ( .A(\u_decoder/fir_filter/dp_cluster_0/r166/A1[7] ), .B(n1814), 
        .C(\u_decoder/fir_filter/dp_cluster_0/r166/A2[7] ), .Q(n2472) );
  OAI212 U4508 ( .A(n2477), .B(n2478), .C(n2479), .Q(
        \u_decoder/fir_filter/I_data_mult_3 [10]) );
  OAI222 U4509 ( .A(\u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[7][5] ), 
        .B(\u_decoder/fir_filter/dp_cluster_0/r167/A2[11] ), .C(
        \u_decoder/fir_filter/dp_cluster_0/r167/A1[8] ), .D(
        \u_decoder/fir_filter/dp_cluster_0/r167/A2[8] ), .Q(n2488) );
  OAI212 U4510 ( .A(\u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[7][5] ), 
        .B(n2484), .C(\u_decoder/fir_filter/dp_cluster_0/r167/A2[11] ), .Q(
        n2489) );
  OAI212 U4511 ( .A(n2487), .B(n1842), .C(n2490), .Q(n2484) );
  OAI212 U4512 ( .A(n2478), .B(n2486), .C(n2476), .Q(n2491) );
  OAI212 U4513 ( .A(n2487), .B(n2493), .C(n2490), .Q(n2492) );
  OAI212 U4514 ( .A(n2477), .B(n2495), .C(n2478), .Q(n2474) );
  IMAJ31 U4515 ( .A(\u_decoder/fir_filter/dp_cluster_0/r167/A2[7] ), .B(n2482), 
        .C(\u_decoder/fir_filter/dp_cluster_0/r167/A1[7] ), .Q(n2477) );
  OAI212 U4516 ( .A(n2499), .B(n2500), .C(n2501), .Q(
        \u_decoder/fir_filter/I_data_mult_4 [10]) );
  XOR31 U4517 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_276/A1[7] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/A2[7] ), .C(n2504), .Q(
        \u_decoder/fir_filter/I_data_mult_4 [9]) );
  OAI222 U4518 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[7][5] ), 
        .B(\u_decoder/fir_filter/dp_cluster_0/mult_276/A2[11] ), .C(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/A1[8] ), .D(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/A2[8] ), .Q(n2510) );
  OAI212 U4519 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[7][5] ), 
        .B(n2506), .C(\u_decoder/fir_filter/dp_cluster_0/mult_276/A2[11] ), 
        .Q(n2511) );
  OAI212 U4520 ( .A(n2509), .B(n1826), .C(n2512), .Q(n2506) );
  OAI212 U4521 ( .A(n2500), .B(n2508), .C(n2498), .Q(n2513) );
  XOR31 U4522 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_276/A2[11] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[7][5] ), .C(n2514), 
        .Q(\u_decoder/fir_filter/I_data_mult_4 [13]) );
  OAI212 U4523 ( .A(n2509), .B(n2515), .C(n2512), .Q(n2514) );
  OAI212 U4524 ( .A(n2499), .B(n2517), .C(n2500), .Q(n2496) );
  IMAJ31 U4525 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_276/A2[7] ), .B(
        n2504), .C(\u_decoder/fir_filter/dp_cluster_0/mult_276/A1[7] ), .Q(
        n2499) );
  OAI212 U4526 ( .A(n73), .B(n7), .C(n2518), .Q(n2519) );
  OAI212 U4527 ( .A(\u_decoder/fir_filter/Q_data_mult_0_buff [2]), .B(n2519), 
        .C(\u_decoder/fir_filter/Q_data_add_1_buff [2]), .Q(n2520) );
  OAI212 U4528 ( .A(n1987), .B(n71), .C(n2520), .Q(n2521) );
  OAI212 U4529 ( .A(\u_decoder/fir_filter/Q_data_mult_0_buff [3]), .B(n2521), 
        .C(\u_decoder/fir_filter/Q_data_add_1_buff [3]), .Q(n2522) );
  OAI212 U4530 ( .A(n1985), .B(n112), .C(n2522), .Q(n2523) );
  OAI212 U4531 ( .A(\u_decoder/fir_filter/Q_data_mult_0_buff [4]), .B(n2523), 
        .C(\u_decoder/fir_filter/Q_data_add_1_buff [4]), .Q(n2524) );
  OAI212 U4532 ( .A(n1983), .B(n128), .C(n2524), .Q(n2525) );
  OAI212 U4533 ( .A(\u_decoder/fir_filter/Q_data_mult_0_buff [5]), .B(n2525), 
        .C(\u_decoder/fir_filter/Q_data_add_1_buff [5]), .Q(n2526) );
  OAI212 U4534 ( .A(n1981), .B(n129), .C(n2526), .Q(n2527) );
  OAI212 U4535 ( .A(\u_decoder/fir_filter/Q_data_mult_0_buff [6]), .B(n2527), 
        .C(\u_decoder/fir_filter/Q_data_add_1_buff [6]), .Q(n2528) );
  OAI212 U4536 ( .A(n1979), .B(n142), .C(n2528), .Q(n2530) );
  OAI212 U4537 ( .A(\u_decoder/fir_filter/Q_data_mult_0_buff [7]), .B(n2530), 
        .C(\u_decoder/fir_filter/Q_data_add_1_buff [7]), .Q(n2529) );
  OAI212 U4538 ( .A(\u_decoder/fir_filter/Q_data_mult_0_buff [8]), .B(n1975), 
        .C(\u_decoder/fir_filter/Q_data_add_1_buff [8]), .Q(n2531) );
  OAI212 U4539 ( .A(n2532), .B(n198), .C(n2531), .Q(n2534) );
  OAI212 U4540 ( .A(\u_decoder/fir_filter/Q_data_mult_0_buff [9]), .B(n2534), 
        .C(\u_decoder/fir_filter/Q_data_add_1_buff [9]), .Q(n2533) );
  OAI212 U4541 ( .A(\u_decoder/fir_filter/Q_data_mult_0_buff [10]), .B(n1971), 
        .C(\u_decoder/fir_filter/Q_data_add_1_buff [10]), .Q(n2535) );
  OAI212 U4542 ( .A(n2536), .B(n258), .C(n2535), .Q(
        \u_decoder/fir_filter/add_326/carry [11]) );
  OAI212 U4543 ( .A(n74), .B(n8), .C(n2537), .Q(n2538) );
  OAI212 U4544 ( .A(\u_decoder/fir_filter/I_data_mult_0_buff [2]), .B(n2538), 
        .C(\u_decoder/fir_filter/I_data_add_1_buff [2]), .Q(n2539) );
  OAI212 U4545 ( .A(n2107), .B(n72), .C(n2539), .Q(n2540) );
  OAI212 U4546 ( .A(\u_decoder/fir_filter/I_data_mult_0_buff [3]), .B(n2540), 
        .C(\u_decoder/fir_filter/I_data_add_1_buff [3]), .Q(n2541) );
  OAI212 U4547 ( .A(n2105), .B(n113), .C(n2541), .Q(n2542) );
  OAI212 U4548 ( .A(\u_decoder/fir_filter/I_data_mult_0_buff [4]), .B(n2542), 
        .C(\u_decoder/fir_filter/I_data_add_1_buff [4]), .Q(n2543) );
  OAI212 U4549 ( .A(n2103), .B(n130), .C(n2543), .Q(n2544) );
  OAI212 U4550 ( .A(\u_decoder/fir_filter/I_data_mult_0_buff [5]), .B(n2544), 
        .C(\u_decoder/fir_filter/I_data_add_1_buff [5]), .Q(n2545) );
  OAI212 U4551 ( .A(n2101), .B(n131), .C(n2545), .Q(n2546) );
  OAI212 U4552 ( .A(\u_decoder/fir_filter/I_data_mult_0_buff [6]), .B(n2546), 
        .C(\u_decoder/fir_filter/I_data_add_1_buff [6]), .Q(n2547) );
  OAI212 U4553 ( .A(n2099), .B(n143), .C(n2547), .Q(n2549) );
  OAI212 U4554 ( .A(\u_decoder/fir_filter/I_data_mult_0_buff [7]), .B(n2549), 
        .C(\u_decoder/fir_filter/I_data_add_1_buff [7]), .Q(n2548) );
  OAI212 U4555 ( .A(\u_decoder/fir_filter/I_data_mult_0_buff [8]), .B(n2095), 
        .C(\u_decoder/fir_filter/I_data_add_1_buff [8]), .Q(n2550) );
  OAI212 U4556 ( .A(n2551), .B(n199), .C(n2550), .Q(n2553) );
  OAI212 U4557 ( .A(\u_decoder/fir_filter/I_data_mult_0_buff [9]), .B(n2553), 
        .C(\u_decoder/fir_filter/I_data_add_1_buff [9]), .Q(n2552) );
  OAI212 U4558 ( .A(\u_decoder/fir_filter/I_data_mult_0_buff [10]), .B(n2091), 
        .C(\u_decoder/fir_filter/I_data_add_1_buff [10]), .Q(n2554) );
  OAI212 U4559 ( .A(n2555), .B(n259), .C(n2554), .Q(
        \u_decoder/fir_filter/add_294/carry [11]) );
  OAI212 U4560 ( .A(n168), .B(n32), .C(n2556), .Q(n2557) );
  OAI212 U4561 ( .A(\u_cordic/mycordic/present_Q_table[5][2] ), .B(n2557), .C(
        \u_cordic/mycordic/present_I_table[5][6] ), .Q(n2558) );
  OAI212 U4562 ( .A(n2212), .B(n156), .C(n2558), .Q(n2560) );
  OAI212 U4563 ( .A(\u_cordic/mycordic/present_Q_table[5][3] ), .B(n2560), .C(
        \u_cordic/mycordic/present_I_table[5][7] ), .Q(n2559) );
  OAI212 U4564 ( .A(\u_cordic/mycordic/present_Q_table[5][4] ), .B(n2208), .C(
        \u_cordic/mycordic/present_I_table[5][7] ), .Q(n2561) );
  OAI212 U4565 ( .A(n2562), .B(n217), .C(n2561), .Q(n2564) );
  OAI212 U4566 ( .A(\u_cordic/mycordic/present_Q_table[5][5] ), .B(n2564), .C(
        \u_cordic/mycordic/present_I_table[5][7] ), .Q(n2563) );
  OAI212 U4567 ( .A(\u_cordic/mycordic/present_Q_table[5][6] ), .B(n2204), .C(
        \u_cordic/mycordic/present_I_table[5][7] ), .Q(n2565) );
  OAI212 U4568 ( .A(n2566), .B(n269), .C(n2565), .Q(
        \u_cordic/mycordic/add_228/carry[7] ) );
  OAI222 U4569 ( .A(n2570), .B(n156), .C(
        \u_cordic/mycordic/present_I_table[5][6] ), .D(n2211), .Q(n2572) );
  OAI212 U4570 ( .A(\u_cordic/mycordic/present_Q_table[5][3] ), .B(n2572), .C(
        n182), .Q(n2571) );
  OAI212 U4571 ( .A(n2574), .B(n217), .C(n2207), .Q(n2576) );
  OAI212 U4572 ( .A(\u_cordic/mycordic/present_Q_table[5][5] ), .B(n2576), .C(
        n182), .Q(n2575) );
  OAI212 U4573 ( .A(n2578), .B(n269), .C(n2203), .Q(
        \u_cordic/mycordic/sub_223/carry[7] ) );
  OAI222 U4574 ( .A(n2580), .B(n201), .C(
        \u_cordic/mycordic/present_Q_table[4][4] ), .D(n2579), .Q(n2582) );
  OAI222 U4575 ( .A(n2584), .B(n155), .C(
        \u_cordic/mycordic/present_Q_table[4][6] ), .D(n2583), .Q(
        \u_cordic/mycordic/sub_216/carry [4]) );
  OAI212 U4576 ( .A(\u_cordic/mycordic/present_I_table[4][2] ), .B(n2219), .C(
        \u_cordic/mycordic/present_Q_table[4][5] ), .Q(n2586) );
  OAI212 U4577 ( .A(n2587), .B(n232), .C(n2586), .Q(n2589) );
  OAI212 U4578 ( .A(\u_cordic/mycordic/present_I_table[4][3] ), .B(n2589), .C(
        \u_cordic/mycordic/present_Q_table[4][6] ), .Q(n2588) );
  OAI222 U4579 ( .A(n1141), .B(n276), .C(n1142), .D(n1141), .Q(n2610) );
  OAI212 U4580 ( .A(\u_coder/n259 ), .B(\u_coder/n69 ), .C(\u_coder/stateQ[0] ), .Q(\u_coder/N1149 ) );
  OAI212 U4581 ( .A(\u_coder/n261 ), .B(\u_coder/n69 ), .C(\u_coder/stateI[0] ), .Q(\u_coder/N1143 ) );
endmodule

