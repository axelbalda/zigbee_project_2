
module TOP ( inClock, inReset, in_inFIFO_inData, in_outFIFO_inReadEnable, 
        in_DEMUX_inDEMUX1, in_DEMUX_inDEMUX2, in_DEMUX_inDEMUX17, 
        in_DEMUX_inDEMUX18, in_DEMUX_inSEL1, in_DEMUX_inSEL2, in_MUX_inSEL3, 
        in_MUX_inSEL6, in_MUX_inSEL9, in_MUX_inSEL11, in_MUX_inSEL12, 
        in_MUX_inSEL15, in_DEMUX_inSEL17, out_MUX_outMUX9, out_MUX_outMUX10, 
        out_MUX_outMUX15, out_MUX_outMUX16 );
  input [3:0] in_inFIFO_inData;
  input [3:0] in_DEMUX_inDEMUX17;
  input [3:0] in_DEMUX_inDEMUX18;
  input [2:0] in_DEMUX_inSEL1;
  input [2:0] in_DEMUX_inSEL2;
  input [1:0] in_MUX_inSEL6;
  input [1:0] in_MUX_inSEL9;
  input [1:0] in_MUX_inSEL15;
  output [3:0] out_MUX_outMUX9;
  output [3:0] out_MUX_outMUX10;
  input inClock, inReset, in_outFIFO_inReadEnable, in_DEMUX_inDEMUX1,
         in_DEMUX_inDEMUX2, in_MUX_inSEL3, in_MUX_inSEL11, in_MUX_inSEL12,
         in_DEMUX_inSEL17;
  output out_MUX_outMUX15, out_MUX_outMUX16;
  wire   \sig_MUX_inMUX3[0] , \sig_MUX_inMUX4[0] , \sig_MUX_inMUX5[0] ,
         \sig_MUX_inMUX8[0] , sig_MUX_outMUX8, \sig_MUX_inMUX11[0] ,
         \sig_MUX_inMUX14[0] , \sig_MUX_inMUX12[0] , \sig_MUX_inMUX13[0] ,
         \u_inFIFO/n751 , \u_inFIFO/n750 , \u_inFIFO/n749 , \u_inFIFO/n748 ,
         \u_inFIFO/n747 , \u_inFIFO/n746 , \u_inFIFO/n745 , \u_inFIFO/n744 ,
         \u_inFIFO/n743 , \u_inFIFO/n742 , \u_inFIFO/n741 , \u_inFIFO/n740 ,
         \u_inFIFO/n739 , \u_inFIFO/n738 , \u_inFIFO/n737 , \u_inFIFO/n736 ,
         \u_inFIFO/n735 , \u_inFIFO/n734 , \u_inFIFO/n733 , \u_inFIFO/n732 ,
         \u_inFIFO/n731 , \u_inFIFO/n730 , \u_inFIFO/n729 , \u_inFIFO/n728 ,
         \u_inFIFO/n727 , \u_inFIFO/n726 , \u_inFIFO/n725 , \u_inFIFO/n724 ,
         \u_inFIFO/n723 , \u_inFIFO/n722 , \u_inFIFO/n721 , \u_inFIFO/n720 ,
         \u_inFIFO/n719 , \u_inFIFO/n718 , \u_inFIFO/n717 , \u_inFIFO/n716 ,
         \u_inFIFO/n715 , \u_inFIFO/n714 , \u_inFIFO/n713 , \u_inFIFO/n712 ,
         \u_inFIFO/n711 , \u_inFIFO/n710 , \u_inFIFO/n709 , \u_inFIFO/n708 ,
         \u_inFIFO/n707 , \u_inFIFO/n706 , \u_inFIFO/n705 , \u_inFIFO/n704 ,
         \u_inFIFO/n703 , \u_inFIFO/n702 , \u_inFIFO/n701 , \u_inFIFO/n700 ,
         \u_inFIFO/n699 , \u_inFIFO/n698 , \u_inFIFO/n697 , \u_inFIFO/n696 ,
         \u_inFIFO/n695 , \u_inFIFO/n694 , \u_inFIFO/n693 , \u_inFIFO/n692 ,
         \u_inFIFO/n691 , \u_inFIFO/n690 , \u_inFIFO/n689 , \u_inFIFO/n688 ,
         \u_inFIFO/n687 , \u_inFIFO/n686 , \u_inFIFO/n685 , \u_inFIFO/n684 ,
         \u_inFIFO/n683 , \u_inFIFO/n682 , \u_inFIFO/n681 , \u_inFIFO/n680 ,
         \u_inFIFO/n679 , \u_inFIFO/n678 , \u_inFIFO/n677 , \u_inFIFO/n676 ,
         \u_inFIFO/n675 , \u_inFIFO/n674 , \u_inFIFO/n673 , \u_inFIFO/n672 ,
         \u_inFIFO/n671 , \u_inFIFO/n670 , \u_inFIFO/n669 , \u_inFIFO/n668 ,
         \u_inFIFO/n667 , \u_inFIFO/n666 , \u_inFIFO/n665 , \u_inFIFO/n664 ,
         \u_inFIFO/n663 , \u_inFIFO/n662 , \u_inFIFO/n661 , \u_inFIFO/n660 ,
         \u_inFIFO/n659 , \u_inFIFO/n658 , \u_inFIFO/n657 , \u_inFIFO/n656 ,
         \u_inFIFO/n655 , \u_inFIFO/n654 , \u_inFIFO/n653 , \u_inFIFO/n652 ,
         \u_inFIFO/n651 , \u_inFIFO/n650 , \u_inFIFO/n649 , \u_inFIFO/n648 ,
         \u_inFIFO/n647 , \u_inFIFO/n646 , \u_inFIFO/n645 , \u_inFIFO/n644 ,
         \u_inFIFO/n643 , \u_inFIFO/n642 , \u_inFIFO/n641 , \u_inFIFO/n640 ,
         \u_inFIFO/n639 , \u_inFIFO/n638 , \u_inFIFO/n637 , \u_inFIFO/n636 ,
         \u_inFIFO/n635 , \u_inFIFO/n634 , \u_inFIFO/n633 , \u_inFIFO/n632 ,
         \u_inFIFO/n631 , \u_inFIFO/n630 , \u_inFIFO/n629 , \u_inFIFO/n628 ,
         \u_inFIFO/n627 , \u_inFIFO/n626 , \u_inFIFO/n625 , \u_inFIFO/n624 ,
         \u_inFIFO/n623 , \u_inFIFO/n622 , \u_inFIFO/n621 , \u_inFIFO/n620 ,
         \u_inFIFO/n619 , \u_inFIFO/n618 , \u_inFIFO/n617 , \u_inFIFO/n616 ,
         \u_inFIFO/n615 , \u_inFIFO/n614 , \u_inFIFO/n613 , \u_inFIFO/n612 ,
         \u_inFIFO/n611 , \u_inFIFO/n610 , \u_inFIFO/n609 , \u_inFIFO/n608 ,
         \u_inFIFO/n607 , \u_inFIFO/n606 , \u_inFIFO/n605 , \u_inFIFO/n604 ,
         \u_inFIFO/n603 , \u_inFIFO/n602 , \u_inFIFO/n601 , \u_inFIFO/n600 ,
         \u_inFIFO/n599 , \u_inFIFO/n598 , \u_inFIFO/n597 , \u_inFIFO/n596 ,
         \u_inFIFO/n595 , \u_inFIFO/n594 , \u_inFIFO/n593 , \u_inFIFO/n592 ,
         \u_inFIFO/n591 , \u_inFIFO/n590 , \u_inFIFO/n589 , \u_inFIFO/n588 ,
         \u_inFIFO/n587 , \u_inFIFO/n586 , \u_inFIFO/n585 , \u_inFIFO/n584 ,
         \u_inFIFO/n582 , \u_inFIFO/n581 , \u_inFIFO/n580 , \u_inFIFO/n579 ,
         \u_inFIFO/n578 , \u_inFIFO/n577 , \u_inFIFO/n576 , \u_inFIFO/n575 ,
         \u_inFIFO/n574 , \u_inFIFO/n573 , \u_inFIFO/n572 , \u_inFIFO/n570 ,
         \u_inFIFO/n569 , \u_inFIFO/n568 , \u_inFIFO/n567 , \u_inFIFO/n566 ,
         \u_inFIFO/n565 , \u_inFIFO/n564 , \u_inFIFO/n563 , \u_inFIFO/n562 ,
         \u_inFIFO/n561 , \u_inFIFO/n560 , \u_inFIFO/n559 , \u_inFIFO/n558 ,
         \u_inFIFO/n557 , \u_inFIFO/n556 , \u_inFIFO/n555 , \u_inFIFO/n554 ,
         \u_inFIFO/n553 , \u_inFIFO/n552 , \u_inFIFO/n551 , \u_inFIFO/n550 ,
         \u_inFIFO/n549 , \u_inFIFO/n548 , \u_inFIFO/n547 , \u_inFIFO/n546 ,
         \u_inFIFO/n545 , \u_inFIFO/n544 , \u_inFIFO/n543 , \u_inFIFO/n542 ,
         \u_inFIFO/n541 , \u_inFIFO/n540 , \u_inFIFO/n539 , \u_inFIFO/n538 ,
         \u_inFIFO/n537 , \u_inFIFO/n536 , \u_inFIFO/n535 , \u_inFIFO/n534 ,
         \u_inFIFO/n533 , \u_inFIFO/n532 , \u_inFIFO/n531 , \u_inFIFO/n530 ,
         \u_inFIFO/n529 , \u_inFIFO/n528 , \u_inFIFO/n527 , \u_inFIFO/n526 ,
         \u_inFIFO/n525 , \u_inFIFO/n524 , \u_inFIFO/n523 , \u_inFIFO/n522 ,
         \u_inFIFO/n521 , \u_inFIFO/n520 , \u_inFIFO/n519 , \u_inFIFO/n518 ,
         \u_inFIFO/n517 , \u_inFIFO/n516 , \u_inFIFO/n515 , \u_inFIFO/n514 ,
         \u_inFIFO/n513 , \u_inFIFO/n512 , \u_inFIFO/n511 , \u_inFIFO/n510 ,
         \u_inFIFO/n509 , \u_inFIFO/n508 , \u_inFIFO/n507 , \u_inFIFO/n506 ,
         \u_inFIFO/n505 , \u_inFIFO/n504 , \u_inFIFO/n503 , \u_inFIFO/n502 ,
         \u_inFIFO/n501 , \u_inFIFO/n500 , \u_inFIFO/n499 , \u_inFIFO/n498 ,
         \u_inFIFO/n497 , \u_inFIFO/n496 , \u_inFIFO/n495 , \u_inFIFO/n494 ,
         \u_inFIFO/n493 , \u_inFIFO/n492 , \u_inFIFO/n491 , \u_inFIFO/n490 ,
         \u_inFIFO/n489 , \u_inFIFO/n488 , \u_inFIFO/n487 , \u_inFIFO/n486 ,
         \u_inFIFO/n485 , \u_inFIFO/n484 , \u_inFIFO/n483 , \u_inFIFO/n482 ,
         \u_inFIFO/n481 , \u_inFIFO/n480 , \u_inFIFO/n479 , \u_inFIFO/n478 ,
         \u_inFIFO/n477 , \u_inFIFO/n476 , \u_inFIFO/n475 , \u_inFIFO/n474 ,
         \u_inFIFO/n473 , \u_inFIFO/n472 , \u_inFIFO/n471 , \u_inFIFO/n470 ,
         \u_inFIFO/n469 , \u_inFIFO/n468 , \u_inFIFO/n467 , \u_inFIFO/n466 ,
         \u_inFIFO/n465 , \u_inFIFO/n464 , \u_inFIFO/n463 , \u_inFIFO/n462 ,
         \u_inFIFO/n461 , \u_inFIFO/n460 , \u_inFIFO/n459 , \u_inFIFO/n458 ,
         \u_inFIFO/n457 , \u_inFIFO/n456 , \u_inFIFO/n455 , \u_inFIFO/n454 ,
         \u_inFIFO/n453 , \u_inFIFO/n452 , \u_inFIFO/n451 , \u_inFIFO/n450 ,
         \u_inFIFO/n449 , \u_inFIFO/n448 , \u_inFIFO/n447 , \u_inFIFO/n446 ,
         \u_inFIFO/n445 , \u_inFIFO/n444 , \u_inFIFO/n443 , \u_inFIFO/n442 ,
         \u_inFIFO/n441 , \u_inFIFO/n440 , \u_inFIFO/n439 , \u_inFIFO/n438 ,
         \u_inFIFO/n437 , \u_inFIFO/n436 , \u_inFIFO/n435 , \u_inFIFO/n434 ,
         \u_inFIFO/n433 , \u_inFIFO/n432 , \u_inFIFO/n431 , \u_inFIFO/n430 ,
         \u_inFIFO/n429 , \u_inFIFO/n428 , \u_inFIFO/n427 , \u_inFIFO/n426 ,
         \u_inFIFO/n425 , \u_inFIFO/n424 , \u_inFIFO/n423 , \u_inFIFO/n422 ,
         \u_inFIFO/n421 , \u_inFIFO/n420 , \u_inFIFO/n419 , \u_inFIFO/n418 ,
         \u_inFIFO/n417 , \u_inFIFO/n416 , \u_inFIFO/n415 , \u_inFIFO/n414 ,
         \u_inFIFO/n413 , \u_inFIFO/n412 , \u_inFIFO/n411 , \u_inFIFO/n410 ,
         \u_inFIFO/n409 , \u_inFIFO/n408 , \u_inFIFO/n407 , \u_inFIFO/n406 ,
         \u_inFIFO/n405 , \u_inFIFO/n404 , \u_inFIFO/n403 , \u_inFIFO/n402 ,
         \u_inFIFO/n401 , \u_inFIFO/n400 , \u_inFIFO/n399 , \u_inFIFO/n398 ,
         \u_inFIFO/n397 , \u_inFIFO/n396 , \u_inFIFO/n395 , \u_inFIFO/n394 ,
         \u_inFIFO/n393 , \u_inFIFO/n392 , \u_inFIFO/n391 , \u_inFIFO/n390 ,
         \u_inFIFO/n389 , \u_inFIFO/n388 , \u_inFIFO/n387 , \u_inFIFO/n386 ,
         \u_inFIFO/n385 , \u_inFIFO/n384 , \u_inFIFO/n383 , \u_inFIFO/n382 ,
         \u_inFIFO/n381 , \u_inFIFO/n380 , \u_inFIFO/n379 , \u_inFIFO/n378 ,
         \u_inFIFO/n377 , \u_inFIFO/n376 , \u_inFIFO/n375 , \u_inFIFO/n374 ,
         \u_inFIFO/n373 , \u_inFIFO/n372 , \u_inFIFO/n371 , \u_inFIFO/n370 ,
         \u_inFIFO/n369 , \u_inFIFO/n368 , \u_inFIFO/n367 , \u_inFIFO/n366 ,
         \u_inFIFO/n365 , \u_inFIFO/n364 , \u_inFIFO/n363 , \u_inFIFO/n362 ,
         \u_inFIFO/n361 , \u_inFIFO/n360 , \u_inFIFO/n359 , \u_inFIFO/n358 ,
         \u_inFIFO/n357 , \u_inFIFO/n356 , \u_inFIFO/n355 , \u_inFIFO/n354 ,
         \u_inFIFO/n353 , \u_inFIFO/n352 , \u_inFIFO/n351 , \u_inFIFO/n350 ,
         \u_inFIFO/n349 , \u_inFIFO/n348 , \u_inFIFO/n347 , \u_inFIFO/n346 ,
         \u_inFIFO/n345 , \u_inFIFO/n344 , \u_inFIFO/n343 , \u_inFIFO/n342 ,
         \u_inFIFO/n341 , \u_inFIFO/n340 , \u_inFIFO/n339 , \u_inFIFO/n338 ,
         \u_inFIFO/n337 , \u_inFIFO/n336 , \u_inFIFO/n335 , \u_inFIFO/n334 ,
         \u_inFIFO/n333 , \u_inFIFO/n332 , \u_inFIFO/n331 , \u_inFIFO/n330 ,
         \u_inFIFO/n329 , \u_inFIFO/n328 , \u_inFIFO/n327 , \u_inFIFO/n326 ,
         \u_inFIFO/n325 , \u_inFIFO/n324 , \u_inFIFO/n323 , \u_inFIFO/n322 ,
         \u_inFIFO/n321 , \u_inFIFO/n320 , \u_inFIFO/n319 , \u_inFIFO/n318 ,
         \u_inFIFO/n317 , \u_inFIFO/n316 , \u_inFIFO/n315 , \u_inFIFO/n314 ,
         \u_inFIFO/n313 , \u_inFIFO/n312 , \u_inFIFO/n311 , \u_inFIFO/n310 ,
         \u_inFIFO/n309 , \u_inFIFO/n308 , \u_inFIFO/n307 , \u_inFIFO/n306 ,
         \u_inFIFO/n305 , \u_inFIFO/n304 , \u_inFIFO/n303 , \u_inFIFO/n302 ,
         \u_inFIFO/n301 , \u_inFIFO/n300 , \u_inFIFO/n299 , \u_inFIFO/n298 ,
         \u_inFIFO/n297 , \u_inFIFO/n296 , \u_inFIFO/n295 , \u_inFIFO/n294 ,
         \u_inFIFO/n293 , \u_inFIFO/n292 , \u_inFIFO/n291 , \u_inFIFO/n290 ,
         \u_inFIFO/n289 , \u_inFIFO/n288 , \u_inFIFO/n287 , \u_inFIFO/n286 ,
         \u_inFIFO/n285 , \u_inFIFO/n284 , \u_inFIFO/n283 , \u_inFIFO/n282 ,
         \u_inFIFO/n281 , \u_inFIFO/n280 , \u_inFIFO/n279 , \u_inFIFO/n278 ,
         \u_inFIFO/n277 , \u_inFIFO/n276 , \u_inFIFO/n275 , \u_inFIFO/n274 ,
         \u_inFIFO/n273 , \u_inFIFO/n272 , \u_inFIFO/n271 , \u_inFIFO/n270 ,
         \u_inFIFO/n269 , \u_inFIFO/n268 , \u_inFIFO/n267 , \u_inFIFO/n266 ,
         \u_inFIFO/n265 , \u_inFIFO/n264 , \u_inFIFO/n263 , \u_inFIFO/n262 ,
         \u_inFIFO/n261 , \u_inFIFO/n260 , \u_inFIFO/n259 , \u_inFIFO/n258 ,
         \u_inFIFO/n257 , \u_inFIFO/n256 , \u_inFIFO/n255 , \u_inFIFO/n254 ,
         \u_inFIFO/n253 , \u_inFIFO/n252 , \u_inFIFO/n251 , \u_inFIFO/n250 ,
         \u_inFIFO/n249 , \u_inFIFO/n248 , \u_inFIFO/n247 , \u_inFIFO/n246 ,
         \u_inFIFO/n245 , \u_inFIFO/n244 , \u_inFIFO/n243 , \u_inFIFO/n242 ,
         \u_inFIFO/n241 , \u_inFIFO/n240 , \u_inFIFO/n239 , \u_inFIFO/n238 ,
         \u_inFIFO/n237 , \u_inFIFO/n236 , \u_inFIFO/n235 , \u_inFIFO/n234 ,
         \u_inFIFO/n233 , \u_inFIFO/n232 , \u_inFIFO/n231 , \u_inFIFO/n230 ,
         \u_inFIFO/n229 , \u_inFIFO/n228 , \u_inFIFO/n227 , \u_inFIFO/n226 ,
         \u_inFIFO/n225 , \u_inFIFO/n224 , \u_inFIFO/n223 , \u_inFIFO/n222 ,
         \u_inFIFO/n221 , \u_inFIFO/n220 , \u_inFIFO/n219 , \u_inFIFO/n218 ,
         \u_inFIFO/n217 , \u_inFIFO/n216 , \u_inFIFO/n215 , \u_inFIFO/n212 ,
         \u_inFIFO/n207 , \u_inFIFO/n206 , \u_inFIFO/n205 , \u_inFIFO/n204 ,
         \u_inFIFO/n203 , \u_inFIFO/n202 , \u_inFIFO/n201 , \u_inFIFO/n200 ,
         \u_inFIFO/n198 , \u_inFIFO/n197 , \u_inFIFO/n188 , \u_inFIFO/n187 ,
         \u_inFIFO/n186 , \u_inFIFO/n185 , \u_inFIFO/n184 , \u_inFIFO/n183 ,
         \u_inFIFO/n182 , \u_inFIFO/n179 , \u_inFIFO/n177 , \u_inFIFO/n176 ,
         \u_inFIFO/n173 , \u_inFIFO/n154 , \u_inFIFO/N375 , \u_inFIFO/N217 ,
         \u_inFIFO/N216 , \u_inFIFO/N215 , \u_inFIFO/N214 , \u_inFIFO/N213 ,
         \u_inFIFO/N212 , \u_inFIFO/N203 , \u_inFIFO/N202 , \u_inFIFO/N201 ,
         \u_inFIFO/N200 , \u_inFIFO/FIFO[127][3] , \u_inFIFO/FIFO[127][2] ,
         \u_inFIFO/FIFO[127][1] , \u_inFIFO/FIFO[127][0] ,
         \u_inFIFO/FIFO[126][3] , \u_inFIFO/FIFO[126][2] ,
         \u_inFIFO/FIFO[126][1] , \u_inFIFO/FIFO[126][0] ,
         \u_inFIFO/FIFO[125][3] , \u_inFIFO/FIFO[125][2] ,
         \u_inFIFO/FIFO[125][1] , \u_inFIFO/FIFO[125][0] ,
         \u_inFIFO/FIFO[124][3] , \u_inFIFO/FIFO[124][2] ,
         \u_inFIFO/FIFO[124][1] , \u_inFIFO/FIFO[124][0] ,
         \u_inFIFO/FIFO[123][3] , \u_inFIFO/FIFO[123][2] ,
         \u_inFIFO/FIFO[123][1] , \u_inFIFO/FIFO[123][0] ,
         \u_inFIFO/FIFO[122][3] , \u_inFIFO/FIFO[122][2] ,
         \u_inFIFO/FIFO[122][1] , \u_inFIFO/FIFO[122][0] ,
         \u_inFIFO/FIFO[121][3] , \u_inFIFO/FIFO[121][2] ,
         \u_inFIFO/FIFO[121][1] , \u_inFIFO/FIFO[121][0] ,
         \u_inFIFO/FIFO[120][3] , \u_inFIFO/FIFO[120][2] ,
         \u_inFIFO/FIFO[120][1] , \u_inFIFO/FIFO[120][0] ,
         \u_inFIFO/FIFO[119][3] , \u_inFIFO/FIFO[119][2] ,
         \u_inFIFO/FIFO[119][1] , \u_inFIFO/FIFO[119][0] ,
         \u_inFIFO/FIFO[118][3] , \u_inFIFO/FIFO[118][2] ,
         \u_inFIFO/FIFO[118][1] , \u_inFIFO/FIFO[118][0] ,
         \u_inFIFO/FIFO[117][3] , \u_inFIFO/FIFO[117][2] ,
         \u_inFIFO/FIFO[117][1] , \u_inFIFO/FIFO[117][0] ,
         \u_inFIFO/FIFO[116][3] , \u_inFIFO/FIFO[116][2] ,
         \u_inFIFO/FIFO[116][1] , \u_inFIFO/FIFO[116][0] ,
         \u_inFIFO/FIFO[115][3] , \u_inFIFO/FIFO[115][2] ,
         \u_inFIFO/FIFO[115][1] , \u_inFIFO/FIFO[115][0] ,
         \u_inFIFO/FIFO[114][3] , \u_inFIFO/FIFO[114][2] ,
         \u_inFIFO/FIFO[114][1] , \u_inFIFO/FIFO[114][0] ,
         \u_inFIFO/FIFO[113][3] , \u_inFIFO/FIFO[113][2] ,
         \u_inFIFO/FIFO[113][1] , \u_inFIFO/FIFO[113][0] ,
         \u_inFIFO/FIFO[112][3] , \u_inFIFO/FIFO[112][2] ,
         \u_inFIFO/FIFO[112][1] , \u_inFIFO/FIFO[112][0] ,
         \u_inFIFO/FIFO[111][3] , \u_inFIFO/FIFO[111][2] ,
         \u_inFIFO/FIFO[111][1] , \u_inFIFO/FIFO[111][0] ,
         \u_inFIFO/FIFO[110][3] , \u_inFIFO/FIFO[110][2] ,
         \u_inFIFO/FIFO[110][1] , \u_inFIFO/FIFO[110][0] ,
         \u_inFIFO/FIFO[109][3] , \u_inFIFO/FIFO[109][2] ,
         \u_inFIFO/FIFO[109][1] , \u_inFIFO/FIFO[109][0] ,
         \u_inFIFO/FIFO[108][3] , \u_inFIFO/FIFO[108][2] ,
         \u_inFIFO/FIFO[108][1] , \u_inFIFO/FIFO[108][0] ,
         \u_inFIFO/FIFO[107][3] , \u_inFIFO/FIFO[107][2] ,
         \u_inFIFO/FIFO[107][1] , \u_inFIFO/FIFO[107][0] ,
         \u_inFIFO/FIFO[106][3] , \u_inFIFO/FIFO[106][2] ,
         \u_inFIFO/FIFO[106][1] , \u_inFIFO/FIFO[106][0] ,
         \u_inFIFO/FIFO[105][3] , \u_inFIFO/FIFO[105][2] ,
         \u_inFIFO/FIFO[105][1] , \u_inFIFO/FIFO[105][0] ,
         \u_inFIFO/FIFO[104][3] , \u_inFIFO/FIFO[104][2] ,
         \u_inFIFO/FIFO[104][1] , \u_inFIFO/FIFO[104][0] ,
         \u_inFIFO/FIFO[103][3] , \u_inFIFO/FIFO[103][2] ,
         \u_inFIFO/FIFO[103][1] , \u_inFIFO/FIFO[103][0] ,
         \u_inFIFO/FIFO[102][3] , \u_inFIFO/FIFO[102][2] ,
         \u_inFIFO/FIFO[102][1] , \u_inFIFO/FIFO[102][0] ,
         \u_inFIFO/FIFO[101][3] , \u_inFIFO/FIFO[101][2] ,
         \u_inFIFO/FIFO[101][1] , \u_inFIFO/FIFO[101][0] ,
         \u_inFIFO/FIFO[100][3] , \u_inFIFO/FIFO[100][2] ,
         \u_inFIFO/FIFO[100][1] , \u_inFIFO/FIFO[100][0] ,
         \u_inFIFO/FIFO[99][3] , \u_inFIFO/FIFO[99][2] ,
         \u_inFIFO/FIFO[99][1] , \u_inFIFO/FIFO[99][0] ,
         \u_inFIFO/FIFO[98][3] , \u_inFIFO/FIFO[98][2] ,
         \u_inFIFO/FIFO[98][1] , \u_inFIFO/FIFO[98][0] ,
         \u_inFIFO/FIFO[97][3] , \u_inFIFO/FIFO[97][2] ,
         \u_inFIFO/FIFO[97][1] , \u_inFIFO/FIFO[97][0] ,
         \u_inFIFO/FIFO[96][3] , \u_inFIFO/FIFO[96][2] ,
         \u_inFIFO/FIFO[96][1] , \u_inFIFO/FIFO[96][0] ,
         \u_inFIFO/FIFO[95][3] , \u_inFIFO/FIFO[95][2] ,
         \u_inFIFO/FIFO[95][1] , \u_inFIFO/FIFO[95][0] ,
         \u_inFIFO/FIFO[94][3] , \u_inFIFO/FIFO[94][2] ,
         \u_inFIFO/FIFO[94][1] , \u_inFIFO/FIFO[94][0] ,
         \u_inFIFO/FIFO[93][3] , \u_inFIFO/FIFO[93][2] ,
         \u_inFIFO/FIFO[93][1] , \u_inFIFO/FIFO[93][0] ,
         \u_inFIFO/FIFO[92][3] , \u_inFIFO/FIFO[92][2] ,
         \u_inFIFO/FIFO[92][1] , \u_inFIFO/FIFO[92][0] ,
         \u_inFIFO/FIFO[91][3] , \u_inFIFO/FIFO[91][2] ,
         \u_inFIFO/FIFO[91][1] , \u_inFIFO/FIFO[91][0] ,
         \u_inFIFO/FIFO[90][3] , \u_inFIFO/FIFO[90][2] ,
         \u_inFIFO/FIFO[90][1] , \u_inFIFO/FIFO[90][0] ,
         \u_inFIFO/FIFO[89][3] , \u_inFIFO/FIFO[89][2] ,
         \u_inFIFO/FIFO[89][1] , \u_inFIFO/FIFO[89][0] ,
         \u_inFIFO/FIFO[88][3] , \u_inFIFO/FIFO[88][2] ,
         \u_inFIFO/FIFO[88][1] , \u_inFIFO/FIFO[88][0] ,
         \u_inFIFO/FIFO[87][3] , \u_inFIFO/FIFO[87][2] ,
         \u_inFIFO/FIFO[87][1] , \u_inFIFO/FIFO[87][0] ,
         \u_inFIFO/FIFO[86][3] , \u_inFIFO/FIFO[86][2] ,
         \u_inFIFO/FIFO[86][1] , \u_inFIFO/FIFO[86][0] ,
         \u_inFIFO/FIFO[85][3] , \u_inFIFO/FIFO[85][2] ,
         \u_inFIFO/FIFO[85][1] , \u_inFIFO/FIFO[85][0] ,
         \u_inFIFO/FIFO[84][3] , \u_inFIFO/FIFO[84][2] ,
         \u_inFIFO/FIFO[84][1] , \u_inFIFO/FIFO[84][0] ,
         \u_inFIFO/FIFO[83][3] , \u_inFIFO/FIFO[83][2] ,
         \u_inFIFO/FIFO[83][1] , \u_inFIFO/FIFO[83][0] ,
         \u_inFIFO/FIFO[82][3] , \u_inFIFO/FIFO[82][2] ,
         \u_inFIFO/FIFO[82][1] , \u_inFIFO/FIFO[82][0] ,
         \u_inFIFO/FIFO[81][3] , \u_inFIFO/FIFO[81][2] ,
         \u_inFIFO/FIFO[81][1] , \u_inFIFO/FIFO[81][0] ,
         \u_inFIFO/FIFO[80][3] , \u_inFIFO/FIFO[80][2] ,
         \u_inFIFO/FIFO[80][1] , \u_inFIFO/FIFO[80][0] ,
         \u_inFIFO/FIFO[79][3] , \u_inFIFO/FIFO[79][2] ,
         \u_inFIFO/FIFO[79][1] , \u_inFIFO/FIFO[79][0] ,
         \u_inFIFO/FIFO[78][3] , \u_inFIFO/FIFO[78][2] ,
         \u_inFIFO/FIFO[78][1] , \u_inFIFO/FIFO[78][0] ,
         \u_inFIFO/FIFO[77][3] , \u_inFIFO/FIFO[77][2] ,
         \u_inFIFO/FIFO[77][1] , \u_inFIFO/FIFO[77][0] ,
         \u_inFIFO/FIFO[76][3] , \u_inFIFO/FIFO[76][2] ,
         \u_inFIFO/FIFO[76][1] , \u_inFIFO/FIFO[76][0] ,
         \u_inFIFO/FIFO[75][3] , \u_inFIFO/FIFO[75][2] ,
         \u_inFIFO/FIFO[75][1] , \u_inFIFO/FIFO[75][0] ,
         \u_inFIFO/FIFO[74][3] , \u_inFIFO/FIFO[74][2] ,
         \u_inFIFO/FIFO[74][1] , \u_inFIFO/FIFO[74][0] ,
         \u_inFIFO/FIFO[73][3] , \u_inFIFO/FIFO[73][2] ,
         \u_inFIFO/FIFO[73][1] , \u_inFIFO/FIFO[73][0] ,
         \u_inFIFO/FIFO[72][3] , \u_inFIFO/FIFO[72][2] ,
         \u_inFIFO/FIFO[72][1] , \u_inFIFO/FIFO[72][0] ,
         \u_inFIFO/FIFO[71][3] , \u_inFIFO/FIFO[71][2] ,
         \u_inFIFO/FIFO[71][1] , \u_inFIFO/FIFO[71][0] ,
         \u_inFIFO/FIFO[70][3] , \u_inFIFO/FIFO[70][2] ,
         \u_inFIFO/FIFO[70][1] , \u_inFIFO/FIFO[70][0] ,
         \u_inFIFO/FIFO[69][3] , \u_inFIFO/FIFO[69][2] ,
         \u_inFIFO/FIFO[69][1] , \u_inFIFO/FIFO[69][0] ,
         \u_inFIFO/FIFO[68][3] , \u_inFIFO/FIFO[68][2] ,
         \u_inFIFO/FIFO[68][1] , \u_inFIFO/FIFO[68][0] ,
         \u_inFIFO/FIFO[67][3] , \u_inFIFO/FIFO[67][2] ,
         \u_inFIFO/FIFO[67][1] , \u_inFIFO/FIFO[67][0] ,
         \u_inFIFO/FIFO[66][3] , \u_inFIFO/FIFO[66][2] ,
         \u_inFIFO/FIFO[66][1] , \u_inFIFO/FIFO[66][0] ,
         \u_inFIFO/FIFO[65][3] , \u_inFIFO/FIFO[65][2] ,
         \u_inFIFO/FIFO[65][1] , \u_inFIFO/FIFO[65][0] ,
         \u_inFIFO/FIFO[64][3] , \u_inFIFO/FIFO[64][2] ,
         \u_inFIFO/FIFO[64][1] , \u_inFIFO/FIFO[64][0] ,
         \u_inFIFO/FIFO[63][3] , \u_inFIFO/FIFO[63][2] ,
         \u_inFIFO/FIFO[63][1] , \u_inFIFO/FIFO[63][0] ,
         \u_inFIFO/FIFO[62][3] , \u_inFIFO/FIFO[62][2] ,
         \u_inFIFO/FIFO[62][1] , \u_inFIFO/FIFO[62][0] ,
         \u_inFIFO/FIFO[61][3] , \u_inFIFO/FIFO[61][2] ,
         \u_inFIFO/FIFO[61][1] , \u_inFIFO/FIFO[61][0] ,
         \u_inFIFO/FIFO[60][3] , \u_inFIFO/FIFO[60][2] ,
         \u_inFIFO/FIFO[60][1] , \u_inFIFO/FIFO[60][0] ,
         \u_inFIFO/FIFO[59][3] , \u_inFIFO/FIFO[59][2] ,
         \u_inFIFO/FIFO[59][1] , \u_inFIFO/FIFO[59][0] ,
         \u_inFIFO/FIFO[58][3] , \u_inFIFO/FIFO[58][2] ,
         \u_inFIFO/FIFO[58][1] , \u_inFIFO/FIFO[58][0] ,
         \u_inFIFO/FIFO[57][3] , \u_inFIFO/FIFO[57][2] ,
         \u_inFIFO/FIFO[57][1] , \u_inFIFO/FIFO[57][0] ,
         \u_inFIFO/FIFO[56][3] , \u_inFIFO/FIFO[56][2] ,
         \u_inFIFO/FIFO[56][1] , \u_inFIFO/FIFO[56][0] ,
         \u_inFIFO/FIFO[55][3] , \u_inFIFO/FIFO[55][2] ,
         \u_inFIFO/FIFO[55][1] , \u_inFIFO/FIFO[55][0] ,
         \u_inFIFO/FIFO[54][3] , \u_inFIFO/FIFO[54][2] ,
         \u_inFIFO/FIFO[54][1] , \u_inFIFO/FIFO[54][0] ,
         \u_inFIFO/FIFO[53][3] , \u_inFIFO/FIFO[53][2] ,
         \u_inFIFO/FIFO[53][1] , \u_inFIFO/FIFO[53][0] ,
         \u_inFIFO/FIFO[52][3] , \u_inFIFO/FIFO[52][2] ,
         \u_inFIFO/FIFO[52][1] , \u_inFIFO/FIFO[52][0] ,
         \u_inFIFO/FIFO[51][3] , \u_inFIFO/FIFO[51][2] ,
         \u_inFIFO/FIFO[51][1] , \u_inFIFO/FIFO[51][0] ,
         \u_inFIFO/FIFO[50][3] , \u_inFIFO/FIFO[50][2] ,
         \u_inFIFO/FIFO[50][1] , \u_inFIFO/FIFO[50][0] ,
         \u_inFIFO/FIFO[49][3] , \u_inFIFO/FIFO[49][2] ,
         \u_inFIFO/FIFO[49][1] , \u_inFIFO/FIFO[49][0] ,
         \u_inFIFO/FIFO[48][3] , \u_inFIFO/FIFO[48][2] ,
         \u_inFIFO/FIFO[48][1] , \u_inFIFO/FIFO[48][0] ,
         \u_inFIFO/FIFO[47][3] , \u_inFIFO/FIFO[47][2] ,
         \u_inFIFO/FIFO[47][1] , \u_inFIFO/FIFO[47][0] ,
         \u_inFIFO/FIFO[46][3] , \u_inFIFO/FIFO[46][2] ,
         \u_inFIFO/FIFO[46][1] , \u_inFIFO/FIFO[46][0] ,
         \u_inFIFO/FIFO[45][3] , \u_inFIFO/FIFO[45][2] ,
         \u_inFIFO/FIFO[45][1] , \u_inFIFO/FIFO[45][0] ,
         \u_inFIFO/FIFO[44][3] , \u_inFIFO/FIFO[44][2] ,
         \u_inFIFO/FIFO[44][1] , \u_inFIFO/FIFO[44][0] ,
         \u_inFIFO/FIFO[43][3] , \u_inFIFO/FIFO[43][2] ,
         \u_inFIFO/FIFO[43][1] , \u_inFIFO/FIFO[43][0] ,
         \u_inFIFO/FIFO[42][3] , \u_inFIFO/FIFO[42][2] ,
         \u_inFIFO/FIFO[42][1] , \u_inFIFO/FIFO[42][0] ,
         \u_inFIFO/FIFO[41][3] , \u_inFIFO/FIFO[41][2] ,
         \u_inFIFO/FIFO[41][1] , \u_inFIFO/FIFO[41][0] ,
         \u_inFIFO/FIFO[40][3] , \u_inFIFO/FIFO[40][2] ,
         \u_inFIFO/FIFO[40][1] , \u_inFIFO/FIFO[40][0] ,
         \u_inFIFO/FIFO[39][3] , \u_inFIFO/FIFO[39][2] ,
         \u_inFIFO/FIFO[39][1] , \u_inFIFO/FIFO[39][0] ,
         \u_inFIFO/FIFO[38][3] , \u_inFIFO/FIFO[38][2] ,
         \u_inFIFO/FIFO[38][1] , \u_inFIFO/FIFO[38][0] ,
         \u_inFIFO/FIFO[37][3] , \u_inFIFO/FIFO[37][2] ,
         \u_inFIFO/FIFO[37][1] , \u_inFIFO/FIFO[37][0] ,
         \u_inFIFO/FIFO[36][3] , \u_inFIFO/FIFO[36][2] ,
         \u_inFIFO/FIFO[36][1] , \u_inFIFO/FIFO[36][0] ,
         \u_inFIFO/FIFO[35][3] , \u_inFIFO/FIFO[35][2] ,
         \u_inFIFO/FIFO[35][1] , \u_inFIFO/FIFO[35][0] ,
         \u_inFIFO/FIFO[34][3] , \u_inFIFO/FIFO[34][2] ,
         \u_inFIFO/FIFO[34][1] , \u_inFIFO/FIFO[34][0] ,
         \u_inFIFO/FIFO[33][3] , \u_inFIFO/FIFO[33][2] ,
         \u_inFIFO/FIFO[33][1] , \u_inFIFO/FIFO[33][0] ,
         \u_inFIFO/FIFO[32][3] , \u_inFIFO/FIFO[32][2] ,
         \u_inFIFO/FIFO[32][1] , \u_inFIFO/FIFO[32][0] ,
         \u_inFIFO/FIFO[31][3] , \u_inFIFO/FIFO[31][2] ,
         \u_inFIFO/FIFO[31][1] , \u_inFIFO/FIFO[31][0] ,
         \u_inFIFO/FIFO[30][3] , \u_inFIFO/FIFO[30][2] ,
         \u_inFIFO/FIFO[30][1] , \u_inFIFO/FIFO[30][0] ,
         \u_inFIFO/FIFO[29][3] , \u_inFIFO/FIFO[29][2] ,
         \u_inFIFO/FIFO[29][1] , \u_inFIFO/FIFO[29][0] ,
         \u_inFIFO/FIFO[28][3] , \u_inFIFO/FIFO[28][2] ,
         \u_inFIFO/FIFO[28][1] , \u_inFIFO/FIFO[28][0] ,
         \u_inFIFO/FIFO[27][3] , \u_inFIFO/FIFO[27][2] ,
         \u_inFIFO/FIFO[27][1] , \u_inFIFO/FIFO[27][0] ,
         \u_inFIFO/FIFO[26][3] , \u_inFIFO/FIFO[26][2] ,
         \u_inFIFO/FIFO[26][1] , \u_inFIFO/FIFO[26][0] ,
         \u_inFIFO/FIFO[25][3] , \u_inFIFO/FIFO[25][2] ,
         \u_inFIFO/FIFO[25][1] , \u_inFIFO/FIFO[25][0] ,
         \u_inFIFO/FIFO[24][3] , \u_inFIFO/FIFO[24][2] ,
         \u_inFIFO/FIFO[24][1] , \u_inFIFO/FIFO[24][0] ,
         \u_inFIFO/FIFO[23][3] , \u_inFIFO/FIFO[23][2] ,
         \u_inFIFO/FIFO[23][1] , \u_inFIFO/FIFO[23][0] ,
         \u_inFIFO/FIFO[22][3] , \u_inFIFO/FIFO[22][2] ,
         \u_inFIFO/FIFO[22][1] , \u_inFIFO/FIFO[22][0] ,
         \u_inFIFO/FIFO[21][3] , \u_inFIFO/FIFO[21][2] ,
         \u_inFIFO/FIFO[21][1] , \u_inFIFO/FIFO[21][0] ,
         \u_inFIFO/FIFO[20][3] , \u_inFIFO/FIFO[20][2] ,
         \u_inFIFO/FIFO[20][1] , \u_inFIFO/FIFO[20][0] ,
         \u_inFIFO/FIFO[19][3] , \u_inFIFO/FIFO[19][2] ,
         \u_inFIFO/FIFO[19][1] , \u_inFIFO/FIFO[19][0] ,
         \u_inFIFO/FIFO[18][3] , \u_inFIFO/FIFO[18][2] ,
         \u_inFIFO/FIFO[18][1] , \u_inFIFO/FIFO[18][0] ,
         \u_inFIFO/FIFO[17][3] , \u_inFIFO/FIFO[17][2] ,
         \u_inFIFO/FIFO[17][1] , \u_inFIFO/FIFO[17][0] ,
         \u_inFIFO/FIFO[16][3] , \u_inFIFO/FIFO[16][2] ,
         \u_inFIFO/FIFO[16][1] , \u_inFIFO/FIFO[16][0] ,
         \u_inFIFO/FIFO[15][3] , \u_inFIFO/FIFO[15][2] ,
         \u_inFIFO/FIFO[15][1] , \u_inFIFO/FIFO[15][0] ,
         \u_inFIFO/FIFO[14][3] , \u_inFIFO/FIFO[14][2] ,
         \u_inFIFO/FIFO[14][1] , \u_inFIFO/FIFO[14][0] ,
         \u_inFIFO/FIFO[13][3] , \u_inFIFO/FIFO[13][2] ,
         \u_inFIFO/FIFO[13][1] , \u_inFIFO/FIFO[13][0] ,
         \u_inFIFO/FIFO[12][3] , \u_inFIFO/FIFO[12][2] ,
         \u_inFIFO/FIFO[12][1] , \u_inFIFO/FIFO[12][0] ,
         \u_inFIFO/FIFO[11][3] , \u_inFIFO/FIFO[11][2] ,
         \u_inFIFO/FIFO[11][1] , \u_inFIFO/FIFO[11][0] ,
         \u_inFIFO/FIFO[10][3] , \u_inFIFO/FIFO[10][2] ,
         \u_inFIFO/FIFO[10][1] , \u_inFIFO/FIFO[10][0] , \u_inFIFO/FIFO[9][3] ,
         \u_inFIFO/FIFO[9][2] , \u_inFIFO/FIFO[9][1] , \u_inFIFO/FIFO[9][0] ,
         \u_inFIFO/FIFO[8][3] , \u_inFIFO/FIFO[8][2] , \u_inFIFO/FIFO[8][1] ,
         \u_inFIFO/FIFO[8][0] , \u_inFIFO/FIFO[7][3] , \u_inFIFO/FIFO[7][2] ,
         \u_inFIFO/FIFO[7][1] , \u_inFIFO/FIFO[7][0] , \u_inFIFO/FIFO[6][3] ,
         \u_inFIFO/FIFO[6][2] , \u_inFIFO/FIFO[6][1] , \u_inFIFO/FIFO[6][0] ,
         \u_inFIFO/FIFO[5][3] , \u_inFIFO/FIFO[5][2] , \u_inFIFO/FIFO[5][1] ,
         \u_inFIFO/FIFO[5][0] , \u_inFIFO/FIFO[4][3] , \u_inFIFO/FIFO[4][2] ,
         \u_inFIFO/FIFO[4][1] , \u_inFIFO/FIFO[4][0] , \u_inFIFO/FIFO[3][3] ,
         \u_inFIFO/FIFO[3][2] , \u_inFIFO/FIFO[3][1] , \u_inFIFO/FIFO[3][0] ,
         \u_inFIFO/FIFO[2][3] , \u_inFIFO/FIFO[2][2] , \u_inFIFO/FIFO[2][1] ,
         \u_inFIFO/FIFO[2][0] , \u_inFIFO/FIFO[1][3] , \u_inFIFO/FIFO[1][2] ,
         \u_inFIFO/FIFO[1][1] , \u_inFIFO/FIFO[1][0] , \u_inFIFO/FIFO[0][3] ,
         \u_inFIFO/FIFO[0][2] , \u_inFIFO/FIFO[0][1] , \u_inFIFO/FIFO[0][0] ,
         \u_inFIFO/N196 , \u_inFIFO/N149 , \u_inFIFO/N148 , \u_inFIFO/N147 ,
         \u_inFIFO/N146 , \u_inFIFO/N145 , \u_inFIFO/N144 , \u_inFIFO/N143 ,
         \u_inFIFO/N140 , \u_inFIFO/N139 , \u_inFIFO/N138 , \u_inFIFO/N137 ,
         \u_inFIFO/N136 , \u_inFIFO/N135 , \u_inFIFO/N134 , \u_inFIFO/N133 ,
         \u_inFIFO/N131 , \u_inFIFO/N130 , \u_inFIFO/N129 , \u_inFIFO/N128 ,
         \u_inFIFO/N127 , \u_inFIFO/N126 , \u_inFIFO/N124 , \u_inFIFO/N123 ,
         \u_inFIFO/N122 , \u_inFIFO/N121 , \u_inFIFO/N120 , \u_inFIFO/N119 ,
         \u_inFIFO/sigEnableCounter , \u_inFIFO/N50 , \u_inFIFO/N49 ,
         \u_inFIFO/N48 , \u_inFIFO/N47 , \u_inFIFO/sig_fsm_start_W ,
         \u_inFIFO/sig_fsm_start_R , \u_inFIFO/outReadCount[0] ,
         \u_inFIFO/outReadCount[1] , \u_inFIFO/outReadCount[2] ,
         \u_inFIFO/outReadCount[3] , \u_inFIFO/outReadCount[4] ,
         \u_inFIFO/outReadCount[5] , \u_inFIFO/outReadCount[6] ,
         \u_inFIFO/outWriteCount[0] , \u_inFIFO/outWriteCount[1] ,
         \u_inFIFO/outWriteCount[2] , \u_inFIFO/outWriteCount[3] ,
         \u_inFIFO/outWriteCount[4] , \u_inFIFO/outWriteCount[5] ,
         \u_inFIFO/outWriteCount[6] , \u_inFIFO/outWriteCount[7] ,
         \u_inFIFO/N45 , \u_inFIFO/N44 , \u_inFIFO/N43 , \u_inFIFO/N41 ,
         \u_inFIFO/N40 , \u_inFIFO/N38 , \u_coder/n356 , \u_coder/n355 ,
         \u_coder/n354 , \u_coder/n353 , \u_coder/n352 , \u_coder/n351 ,
         \u_coder/n350 , \u_coder/n349 , \u_coder/n348 , \u_coder/n347 ,
         \u_coder/n346 , \u_coder/n345 , \u_coder/n344 , \u_coder/n343 ,
         \u_coder/n342 , \u_coder/n341 , \u_coder/n340 , \u_coder/n339 ,
         \u_coder/n338 , \u_coder/n337 , \u_coder/n336 , \u_coder/n335 ,
         \u_coder/n334 , \u_coder/n333 , \u_coder/n332 , \u_coder/n331 ,
         \u_coder/n330 , \u_coder/n329 , \u_coder/n328 , \u_coder/n327 ,
         \u_coder/n326 , \u_coder/n325 , \u_coder/n324 , \u_coder/n323 ,
         \u_coder/n322 , \u_coder/n321 , \u_coder/n320 , \u_coder/n319 ,
         \u_coder/n318 , \u_coder/n317 , \u_coder/n316 , \u_coder/n315 ,
         \u_coder/n314 , \u_coder/n313 , \u_coder/n312 , \u_coder/n311 ,
         \u_coder/n310 , \u_coder/n309 , \u_coder/n308 , \u_coder/n307 ,
         \u_coder/n306 , \u_coder/n305 , \u_coder/n304 , \u_coder/n303 ,
         \u_coder/n302 , \u_coder/n301 , \u_coder/n300 , \u_coder/n299 ,
         \u_coder/n298 , \u_coder/n297 , \u_coder/n296 , \u_coder/n295 ,
         \u_coder/n294 , \u_coder/n293 , \u_coder/n292 , \u_coder/n291 ,
         \u_coder/n290 , \u_coder/n289 , \u_coder/n288 , \u_coder/n287 ,
         \u_coder/n286 , \u_coder/n284 , \u_coder/n283 , \u_coder/n282 ,
         \u_coder/n281 , \u_coder/n280 , \u_coder/n279 , \u_coder/n278 ,
         \u_coder/n277 , \u_coder/n276 , \u_coder/n275 , \u_coder/n274 ,
         \u_coder/n273 , \u_coder/n272 , \u_coder/n271 , \u_coder/n270 ,
         \u_coder/n269 , \u_coder/n268 , \u_coder/n267 , \u_coder/n266 ,
         \u_coder/n265 , \u_coder/n264 , \u_coder/n263 , \u_coder/n262 ,
         \u_coder/n261 , \u_coder/n260 , \u_coder/n259 , \u_coder/n258 ,
         \u_coder/n257 , \u_coder/n256 , \u_coder/n255 , \u_coder/n254 ,
         \u_coder/n253 , \u_coder/n252 , \u_coder/n251 , \u_coder/n250 ,
         \u_coder/n249 , \u_coder/n248 , \u_coder/n247 , \u_coder/n246 ,
         \u_coder/n245 , \u_coder/n244 , \u_coder/n243 , \u_coder/n242 ,
         \u_coder/n241 , \u_coder/n240 , \u_coder/n239 , \u_coder/n238 ,
         \u_coder/n237 , \u_coder/n236 , \u_coder/n235 , \u_coder/n234 ,
         \u_coder/n233 , \u_coder/n232 , \u_coder/n231 , \u_coder/n230 ,
         \u_coder/n229 , \u_coder/n228 , \u_coder/n227 , \u_coder/n226 ,
         \u_coder/n225 , \u_coder/n224 , \u_coder/n223 , \u_coder/n221 ,
         \u_coder/n220 , \u_coder/n219 , \u_coder/n218 , \u_coder/n217 ,
         \u_coder/n216 , \u_coder/n214 , \u_coder/n213 , \u_coder/n212 ,
         \u_coder/n211 , \u_coder/n210 , \u_coder/n209 , \u_coder/n208 ,
         \u_coder/n207 , \u_coder/n206 , \u_coder/n205 , \u_coder/n204 ,
         \u_coder/n203 , \u_coder/n202 , \u_coder/n201 , \u_coder/n200 ,
         \u_coder/n199 , \u_coder/n198 , \u_coder/n197 , \u_coder/n196 ,
         \u_coder/n195 , \u_coder/n194 , \u_coder/n193 , \u_coder/n192 ,
         \u_coder/n191 , \u_coder/n190 , \u_coder/n189 , \u_coder/n188 ,
         \u_coder/n187 , \u_coder/n186 , \u_coder/n185 , \u_coder/n184 ,
         \u_coder/n183 , \u_coder/n182 , \u_coder/n181 , \u_coder/n180 ,
         \u_coder/n179 , \u_coder/n178 , \u_coder/n177 , \u_coder/n176 ,
         \u_coder/n175 , \u_coder/n174 , \u_coder/n173 , \u_coder/n170 ,
         \u_coder/n169 , \u_coder/n168 , \u_coder/n167 , \u_coder/n166 ,
         \u_coder/n165 , \u_coder/n164 , \u_coder/n163 , \u_coder/n162 ,
         \u_coder/n161 , \u_coder/n160 , \u_coder/n159 , \u_coder/n158 ,
         \u_coder/n157 , \u_coder/n156 , \u_coder/n155 , \u_coder/n154 ,
         \u_coder/n153 , \u_coder/n152 , \u_coder/n151 , \u_coder/n150 ,
         \u_coder/n149 , \u_coder/n148 , \u_coder/n147 , \u_coder/n146 ,
         \u_coder/n145 , \u_coder/n144 , \u_coder/n143 , \u_coder/n142 ,
         \u_coder/n141 , \u_coder/n140 , \u_coder/n139 , \u_coder/n138 ,
         \u_coder/n137 , \u_coder/n136 , \u_coder/n135 , \u_coder/n131 ,
         \u_coder/n130 , \u_coder/n129 , \u_coder/n128 , \u_coder/n127 ,
         \u_coder/n126 , \u_coder/n125 , \u_coder/n123 , \u_coder/n120 ,
         \u_coder/n118 , \u_coder/n117 , \u_coder/n105 , \u_coder/n104 ,
         \u_coder/n103 , \u_coder/n101 , \u_coder/n94 , \u_coder/n91 ,
         \u_coder/n88 , \u_coder/n33 , \u_coder/N1149 , \u_coder/N1143 ,
         \u_coder/N1032 , \u_coder/N1031 , \u_coder/N1030 , \u_coder/N1029 ,
         \u_coder/N1028 , \u_coder/N1027 , \u_coder/N1026 , \u_coder/N1025 ,
         \u_coder/N1024 , \u_coder/N1023 , \u_coder/N1022 , \u_coder/N1021 ,
         \u_coder/N1020 , \u_coder/N1019 , \u_coder/N1018 , \u_coder/N1017 ,
         \u_coder/N1016 , \u_coder/N1015 , \u_coder/N1014 , \u_coder/N974 ,
         \u_coder/N726 , \u_coder/N725 , \u_coder/N724 , \u_coder/N723 ,
         \u_coder/N722 , \u_coder/N721 , \u_coder/N720 , \u_coder/N719 ,
         \u_coder/N718 , \u_coder/N717 , \u_coder/N716 , \u_coder/N715 ,
         \u_coder/N714 , \u_coder/N713 , \u_coder/N712 , \u_coder/N711 ,
         \u_coder/N710 , \u_coder/N709 , \u_coder/N708 , \u_coder/N668 ,
         \u_coder/N522 , \u_coder/N521 , \u_coder/N520 , \u_coder/N519 ,
         \u_coder/N518 , \u_coder/N517 , \u_coder/N516 , \u_coder/N515 ,
         \u_coder/N514 , \u_coder/N513 , \u_coder/N512 , \u_coder/N511 ,
         \u_coder/N510 , \u_coder/N509 , \u_coder/N508 , \u_coder/N507 ,
         \u_coder/N506 , \u_coder/N505 , \u_coder/N504 , \u_coder/N503 ,
         \u_coder/N501 , \u_coder/N499 , \u_coder/my_clk_10M ,
         \u_coder/old_i_data , \u_coder/is9 , \u_coder/isPositiveQ ,
         \u_coder/isPositiveI , \u_coder/sin_was_positiveQ , \u_coder/IorQ ,
         \u_coder/stateQ[0] , \u_coder/stateI[0] , \u_coder/N476 ,
         \u_coder/N475 , \u_coder/N474 , \u_coder/N473 , \u_coder/N472 ,
         \u_coder/N471 , \u_coder/N470 , \u_coder/N469 , \u_coder/N468 ,
         \u_coder/N467 , \u_coder/N466 , \u_coder/N465 , \u_coder/N464 ,
         \u_coder/N463 , \u_coder/N462 , \u_coder/N461 , \u_coder/N460 ,
         \u_coder/N459 , \u_coder/clk_10M , \u_decoder/sample_ready ,
         \u_cordic/n32 , \u_cordic/n31 , \u_cordic/n30 , \u_cordic/n29 ,
         \u_cordic/n28 , \u_cordic/n27 , \u_cordic/n26 , \u_cordic/n25 ,
         \u_cordic/n24 , \u_cordic/n23 , \u_cordic/n22 , \u_cordic/n21 ,
         \u_cordic/n20 , \u_cordic/n19 , \u_cordic/n18 , \u_cordic/n17 ,
         \u_cordic/n16 , \u_cordic/n15 , \u_cordic/n12 , \u_cordic/n11 ,
         \u_cordic/n10 , \u_cordic/n9 , \u_cordic/N16 , \u_cordic/N15 ,
         \u_cordic/N14 , \u_cordic/dir , \u_cdr/n59 , \u_cdr/n58 , \u_cdr/n57 ,
         \u_cdr/n56 , \u_cdr/n55 , \u_cdr/n54 , \u_cdr/n53 , \u_cdr/n52 ,
         \u_cdr/n51 , \u_cdr/n50 , \u_cdr/n49 , \u_cdr/n48 , \u_cdr/n47 ,
         \u_cdr/n46 , \u_cdr/n45 , \u_cdr/n44 , \u_cdr/n43 , \u_cdr/n42 ,
         \u_cdr/n41 , \u_cdr/n40 , \u_cdr/n39 , \u_cdr/n38 , \u_cdr/n37 ,
         \u_cdr/n36 , \u_cdr/n35 , \u_cdr/n34 , \u_cdr/n33 , \u_cdr/n32 ,
         \u_cdr/n31 , \u_cdr/n30 , \u_cdr/n29 , \u_cdr/n28 , \u_cdr/n27 ,
         \u_cdr/n26 , \u_cdr/n25 , \u_cdr/n24 , \u_cdr/n23 , \u_cdr/n20 ,
         \u_cdr/n19 , \u_cdr/n18 , \u_cdr/n17 , \u_cdr/n16 , \u_cdr/n15 ,
         \u_cdr/n14 , \u_cdr/n3 , \u_cdr/N100 , \u_cdr/w_sE , \u_cdr/w_sT ,
         \u_cdr/dir , \u_cdr/flag , \u_outFIFO/n1561 , \u_outFIFO/n1560 ,
         \u_outFIFO/n1559 , \u_outFIFO/n1558 , \u_outFIFO/n1557 ,
         \u_outFIFO/n1556 , \u_outFIFO/n1555 , \u_outFIFO/n1554 ,
         \u_outFIFO/n1553 , \u_outFIFO/n1552 , \u_outFIFO/n1551 ,
         \u_outFIFO/n1550 , \u_outFIFO/n1549 , \u_outFIFO/n1548 ,
         \u_outFIFO/n1547 , \u_outFIFO/n1546 , \u_outFIFO/n1545 ,
         \u_outFIFO/n1544 , \u_outFIFO/n1543 , \u_outFIFO/n1542 ,
         \u_outFIFO/n1541 , \u_outFIFO/n1540 , \u_outFIFO/n1539 ,
         \u_outFIFO/n1538 , \u_outFIFO/n1537 , \u_outFIFO/n1536 ,
         \u_outFIFO/n1535 , \u_outFIFO/n1534 , \u_outFIFO/n1533 ,
         \u_outFIFO/n1532 , \u_outFIFO/n1531 , \u_outFIFO/n1530 ,
         \u_outFIFO/n1529 , \u_outFIFO/n1528 , \u_outFIFO/n1527 ,
         \u_outFIFO/n1526 , \u_outFIFO/n1525 , \u_outFIFO/n1524 ,
         \u_outFIFO/n1523 , \u_outFIFO/n1522 , \u_outFIFO/n1521 ,
         \u_outFIFO/n1520 , \u_outFIFO/n1519 , \u_outFIFO/n1518 ,
         \u_outFIFO/n1517 , \u_outFIFO/n1516 , \u_outFIFO/n1515 ,
         \u_outFIFO/n1514 , \u_outFIFO/n1513 , \u_outFIFO/n1512 ,
         \u_outFIFO/n1511 , \u_outFIFO/n1510 , \u_outFIFO/n1509 ,
         \u_outFIFO/n1508 , \u_outFIFO/n1507 , \u_outFIFO/n1506 ,
         \u_outFIFO/n1505 , \u_outFIFO/n1504 , \u_outFIFO/n1503 ,
         \u_outFIFO/n1502 , \u_outFIFO/n1501 , \u_outFIFO/n1500 ,
         \u_outFIFO/n1499 , \u_outFIFO/n1498 , \u_outFIFO/n1497 ,
         \u_outFIFO/n1496 , \u_outFIFO/n1495 , \u_outFIFO/n1494 ,
         \u_outFIFO/n1493 , \u_outFIFO/n1492 , \u_outFIFO/n1491 ,
         \u_outFIFO/n1490 , \u_outFIFO/n1489 , \u_outFIFO/n1488 ,
         \u_outFIFO/n1487 , \u_outFIFO/n1486 , \u_outFIFO/n1485 ,
         \u_outFIFO/n1484 , \u_outFIFO/n1483 , \u_outFIFO/n1482 ,
         \u_outFIFO/n1481 , \u_outFIFO/n1480 , \u_outFIFO/n1479 ,
         \u_outFIFO/n1478 , \u_outFIFO/n1477 , \u_outFIFO/n1476 ,
         \u_outFIFO/n1475 , \u_outFIFO/n1474 , \u_outFIFO/n1473 ,
         \u_outFIFO/n1472 , \u_outFIFO/n1471 , \u_outFIFO/n1470 ,
         \u_outFIFO/n1469 , \u_outFIFO/n1468 , \u_outFIFO/n1467 ,
         \u_outFIFO/n1466 , \u_outFIFO/n1465 , \u_outFIFO/n1464 ,
         \u_outFIFO/n1463 , \u_outFIFO/n1462 , \u_outFIFO/n1461 ,
         \u_outFIFO/n1460 , \u_outFIFO/n1459 , \u_outFIFO/n1458 ,
         \u_outFIFO/n1457 , \u_outFIFO/n1456 , \u_outFIFO/n1455 ,
         \u_outFIFO/n1454 , \u_outFIFO/n1453 , \u_outFIFO/n1452 ,
         \u_outFIFO/n1451 , \u_outFIFO/n1450 , \u_outFIFO/n1449 ,
         \u_outFIFO/n1448 , \u_outFIFO/n1447 , \u_outFIFO/n1446 ,
         \u_outFIFO/n1445 , \u_outFIFO/n1444 , \u_outFIFO/n1443 ,
         \u_outFIFO/n1442 , \u_outFIFO/n1441 , \u_outFIFO/n1440 ,
         \u_outFIFO/n1439 , \u_outFIFO/n1438 , \u_outFIFO/n1437 ,
         \u_outFIFO/n1436 , \u_outFIFO/n1435 , \u_outFIFO/n1434 ,
         \u_outFIFO/n1433 , \u_outFIFO/n1432 , \u_outFIFO/n1431 ,
         \u_outFIFO/n1430 , \u_outFIFO/n1429 , \u_outFIFO/n1428 ,
         \u_outFIFO/n1427 , \u_outFIFO/n1426 , \u_outFIFO/n1425 ,
         \u_outFIFO/n1424 , \u_outFIFO/n1423 , \u_outFIFO/n1422 ,
         \u_outFIFO/n1421 , \u_outFIFO/n1420 , \u_outFIFO/n1419 ,
         \u_outFIFO/n1418 , \u_outFIFO/n1417 , \u_outFIFO/n1416 ,
         \u_outFIFO/n1415 , \u_outFIFO/n1414 , \u_outFIFO/n1413 ,
         \u_outFIFO/n1412 , \u_outFIFO/n1411 , \u_outFIFO/n1410 ,
         \u_outFIFO/n1409 , \u_outFIFO/n1408 , \u_outFIFO/n1407 ,
         \u_outFIFO/n1406 , \u_outFIFO/n1405 , \u_outFIFO/n1404 ,
         \u_outFIFO/n1403 , \u_outFIFO/n1402 , \u_outFIFO/n1401 ,
         \u_outFIFO/n1400 , \u_outFIFO/n1399 , \u_outFIFO/n1398 ,
         \u_outFIFO/n1397 , \u_outFIFO/n1396 , \u_outFIFO/n1395 ,
         \u_outFIFO/n1394 , \u_outFIFO/n1392 , \u_outFIFO/n1391 ,
         \u_outFIFO/n1390 , \u_outFIFO/n1389 , \u_outFIFO/n1388 ,
         \u_outFIFO/n1387 , \u_outFIFO/n1386 , \u_outFIFO/n1385 ,
         \u_outFIFO/n1384 , \u_outFIFO/n1383 , \u_outFIFO/n1382 ,
         \u_outFIFO/n1381 , \u_outFIFO/n1380 , \u_outFIFO/n1379 ,
         \u_outFIFO/n1378 , \u_outFIFO/n1377 , \u_outFIFO/n1376 ,
         \u_outFIFO/n1375 , \u_outFIFO/n1374 , \u_outFIFO/n1373 ,
         \u_outFIFO/n1372 , \u_outFIFO/n1371 , \u_outFIFO/n1370 ,
         \u_outFIFO/n1369 , \u_outFIFO/n1368 , \u_outFIFO/n1367 ,
         \u_outFIFO/n1366 , \u_outFIFO/n1365 , \u_outFIFO/n1364 ,
         \u_outFIFO/n1363 , \u_outFIFO/n1362 , \u_outFIFO/n1361 ,
         \u_outFIFO/n1360 , \u_outFIFO/n1359 , \u_outFIFO/n1358 ,
         \u_outFIFO/n1357 , \u_outFIFO/n1356 , \u_outFIFO/n1355 ,
         \u_outFIFO/n1354 , \u_outFIFO/n1353 , \u_outFIFO/n1352 ,
         \u_outFIFO/n1351 , \u_outFIFO/n1350 , \u_outFIFO/n1349 ,
         \u_outFIFO/n1348 , \u_outFIFO/n1347 , \u_outFIFO/n1346 ,
         \u_outFIFO/n1345 , \u_outFIFO/n1344 , \u_outFIFO/n1343 ,
         \u_outFIFO/n1342 , \u_outFIFO/n1341 , \u_outFIFO/n1340 ,
         \u_outFIFO/n1339 , \u_outFIFO/n1338 , \u_outFIFO/n1337 ,
         \u_outFIFO/n1336 , \u_outFIFO/n1335 , \u_outFIFO/n1334 ,
         \u_outFIFO/n1333 , \u_outFIFO/n1332 , \u_outFIFO/n1331 ,
         \u_outFIFO/n1330 , \u_outFIFO/n1329 , \u_outFIFO/n1328 ,
         \u_outFIFO/n1327 , \u_outFIFO/n1326 , \u_outFIFO/n1325 ,
         \u_outFIFO/n1324 , \u_outFIFO/n1323 , \u_outFIFO/n1322 ,
         \u_outFIFO/n1321 , \u_outFIFO/n1320 , \u_outFIFO/n1319 ,
         \u_outFIFO/n1318 , \u_outFIFO/n1317 , \u_outFIFO/n1316 ,
         \u_outFIFO/n1315 , \u_outFIFO/n1314 , \u_outFIFO/n1313 ,
         \u_outFIFO/n1312 , \u_outFIFO/n1311 , \u_outFIFO/n1310 ,
         \u_outFIFO/n1309 , \u_outFIFO/n1308 , \u_outFIFO/n1307 ,
         \u_outFIFO/n1306 , \u_outFIFO/n1305 , \u_outFIFO/n1304 ,
         \u_outFIFO/n1303 , \u_outFIFO/n1302 , \u_outFIFO/n1301 ,
         \u_outFIFO/n1300 , \u_outFIFO/n1299 , \u_outFIFO/n1298 ,
         \u_outFIFO/n1297 , \u_outFIFO/n1296 , \u_outFIFO/n1295 ,
         \u_outFIFO/n1294 , \u_outFIFO/n1293 , \u_outFIFO/n1292 ,
         \u_outFIFO/n1291 , \u_outFIFO/n1290 , \u_outFIFO/n1289 ,
         \u_outFIFO/n1288 , \u_outFIFO/n1287 , \u_outFIFO/n1286 ,
         \u_outFIFO/n1285 , \u_outFIFO/n1284 , \u_outFIFO/n1283 ,
         \u_outFIFO/n1282 , \u_outFIFO/n1281 , \u_outFIFO/n1280 ,
         \u_outFIFO/n1279 , \u_outFIFO/n1278 , \u_outFIFO/n1277 ,
         \u_outFIFO/n1276 , \u_outFIFO/n1275 , \u_outFIFO/n1274 ,
         \u_outFIFO/n1273 , \u_outFIFO/n1272 , \u_outFIFO/n1271 ,
         \u_outFIFO/n1270 , \u_outFIFO/n1269 , \u_outFIFO/n1268 ,
         \u_outFIFO/n1267 , \u_outFIFO/n1266 , \u_outFIFO/n1265 ,
         \u_outFIFO/n1264 , \u_outFIFO/n1263 , \u_outFIFO/n1262 ,
         \u_outFIFO/n1261 , \u_outFIFO/n1260 , \u_outFIFO/n1259 ,
         \u_outFIFO/n1258 , \u_outFIFO/n1257 , \u_outFIFO/n1256 ,
         \u_outFIFO/n1255 , \u_outFIFO/n1254 , \u_outFIFO/n1253 ,
         \u_outFIFO/n1252 , \u_outFIFO/n1251 , \u_outFIFO/n1250 ,
         \u_outFIFO/n1249 , \u_outFIFO/n1248 , \u_outFIFO/n1247 ,
         \u_outFIFO/n1246 , \u_outFIFO/n1245 , \u_outFIFO/n1244 ,
         \u_outFIFO/n1243 , \u_outFIFO/n1242 , \u_outFIFO/n1241 ,
         \u_outFIFO/n1240 , \u_outFIFO/n1239 , \u_outFIFO/n1238 ,
         \u_outFIFO/n1237 , \u_outFIFO/n1236 , \u_outFIFO/n1235 ,
         \u_outFIFO/n1234 , \u_outFIFO/n1233 , \u_outFIFO/n1232 ,
         \u_outFIFO/n1231 , \u_outFIFO/n1230 , \u_outFIFO/n1229 ,
         \u_outFIFO/n1228 , \u_outFIFO/n1227 , \u_outFIFO/n1226 ,
         \u_outFIFO/n1225 , \u_outFIFO/n1224 , \u_outFIFO/n1223 ,
         \u_outFIFO/n1222 , \u_outFIFO/n1221 , \u_outFIFO/n1220 ,
         \u_outFIFO/n1219 , \u_outFIFO/n1218 , \u_outFIFO/n1217 ,
         \u_outFIFO/n1216 , \u_outFIFO/n1215 , \u_outFIFO/n1214 ,
         \u_outFIFO/n1213 , \u_outFIFO/n1212 , \u_outFIFO/n1211 ,
         \u_outFIFO/n1210 , \u_outFIFO/n1209 , \u_outFIFO/n1208 ,
         \u_outFIFO/n1207 , \u_outFIFO/n1206 , \u_outFIFO/n1205 ,
         \u_outFIFO/n1204 , \u_outFIFO/n1203 , \u_outFIFO/n1202 ,
         \u_outFIFO/n1201 , \u_outFIFO/n1200 , \u_outFIFO/n1199 ,
         \u_outFIFO/n1198 , \u_outFIFO/n1197 , \u_outFIFO/n1196 ,
         \u_outFIFO/n1195 , \u_outFIFO/n1194 , \u_outFIFO/n1193 ,
         \u_outFIFO/n1192 , \u_outFIFO/n1191 , \u_outFIFO/n1190 ,
         \u_outFIFO/n1189 , \u_outFIFO/n1188 , \u_outFIFO/n1187 ,
         \u_outFIFO/n1186 , \u_outFIFO/n1185 , \u_outFIFO/n1184 ,
         \u_outFIFO/n1183 , \u_outFIFO/n1182 , \u_outFIFO/n1181 ,
         \u_outFIFO/n1180 , \u_outFIFO/n1179 , \u_outFIFO/n1178 ,
         \u_outFIFO/n1177 , \u_outFIFO/n1176 , \u_outFIFO/n1175 ,
         \u_outFIFO/n1174 , \u_outFIFO/n1173 , \u_outFIFO/n1172 ,
         \u_outFIFO/n1171 , \u_outFIFO/n1170 , \u_outFIFO/n1169 ,
         \u_outFIFO/n1168 , \u_outFIFO/n1167 , \u_outFIFO/n1166 ,
         \u_outFIFO/n1165 , \u_outFIFO/n1164 , \u_outFIFO/n1163 ,
         \u_outFIFO/n1162 , \u_outFIFO/n1161 , \u_outFIFO/n1159 ,
         \u_outFIFO/n1158 , \u_outFIFO/n1157 , \u_outFIFO/n1156 ,
         \u_outFIFO/n1155 , \u_outFIFO/n1154 , \u_outFIFO/n1153 ,
         \u_outFIFO/n1152 , \u_outFIFO/n1151 , \u_outFIFO/n1150 ,
         \u_outFIFO/n1149 , \u_outFIFO/n1148 , \u_outFIFO/n1147 ,
         \u_outFIFO/n1146 , \u_outFIFO/n1145 , \u_outFIFO/n1144 ,
         \u_outFIFO/n1143 , \u_outFIFO/n1142 , \u_outFIFO/n1141 ,
         \u_outFIFO/n1140 , \u_outFIFO/n1139 , \u_outFIFO/n1138 ,
         \u_outFIFO/n1137 , \u_outFIFO/n1136 , \u_outFIFO/n1135 ,
         \u_outFIFO/n1134 , \u_outFIFO/n1133 , \u_outFIFO/n1132 ,
         \u_outFIFO/n1131 , \u_outFIFO/n1130 , \u_outFIFO/n1129 ,
         \u_outFIFO/n1128 , \u_outFIFO/n1127 , \u_outFIFO/n1126 ,
         \u_outFIFO/n1125 , \u_outFIFO/n1124 , \u_outFIFO/n1123 ,
         \u_outFIFO/n1122 , \u_outFIFO/n1121 , \u_outFIFO/n1120 ,
         \u_outFIFO/n1119 , \u_outFIFO/n1118 , \u_outFIFO/n1117 ,
         \u_outFIFO/n1116 , \u_outFIFO/n1115 , \u_outFIFO/n1114 ,
         \u_outFIFO/n1113 , \u_outFIFO/n1112 , \u_outFIFO/n1111 ,
         \u_outFIFO/n1110 , \u_outFIFO/n1109 , \u_outFIFO/n1108 ,
         \u_outFIFO/n1107 , \u_outFIFO/n1106 , \u_outFIFO/n1105 ,
         \u_outFIFO/n1104 , \u_outFIFO/n1103 , \u_outFIFO/n1102 ,
         \u_outFIFO/n1101 , \u_outFIFO/n1100 , \u_outFIFO/n1099 ,
         \u_outFIFO/n1098 , \u_outFIFO/n1097 , \u_outFIFO/n1096 ,
         \u_outFIFO/n1095 , \u_outFIFO/n1094 , \u_outFIFO/n1093 ,
         \u_outFIFO/n1092 , \u_outFIFO/n1091 , \u_outFIFO/n1090 ,
         \u_outFIFO/n1089 , \u_outFIFO/n1088 , \u_outFIFO/n1087 ,
         \u_outFIFO/n1086 , \u_outFIFO/n1085 , \u_outFIFO/n1084 ,
         \u_outFIFO/n1083 , \u_outFIFO/n1082 , \u_outFIFO/n1081 ,
         \u_outFIFO/n1080 , \u_outFIFO/n1079 , \u_outFIFO/n1078 ,
         \u_outFIFO/n1077 , \u_outFIFO/n1076 , \u_outFIFO/n1075 ,
         \u_outFIFO/n1074 , \u_outFIFO/n1073 , \u_outFIFO/n1072 ,
         \u_outFIFO/n1071 , \u_outFIFO/n1070 , \u_outFIFO/n1069 ,
         \u_outFIFO/n1068 , \u_outFIFO/n1067 , \u_outFIFO/n1066 ,
         \u_outFIFO/n1065 , \u_outFIFO/n1064 , \u_outFIFO/n1063 ,
         \u_outFIFO/n1062 , \u_outFIFO/n1061 , \u_outFIFO/n1060 ,
         \u_outFIFO/n1059 , \u_outFIFO/n1058 , \u_outFIFO/n1057 ,
         \u_outFIFO/n1056 , \u_outFIFO/n1055 , \u_outFIFO/n1054 ,
         \u_outFIFO/n1053 , \u_outFIFO/n1052 , \u_outFIFO/n1051 ,
         \u_outFIFO/n1050 , \u_outFIFO/n1049 , \u_outFIFO/n1048 ,
         \u_outFIFO/n1047 , \u_outFIFO/n1046 , \u_outFIFO/n1045 ,
         \u_outFIFO/n1044 , \u_outFIFO/n1043 , \u_outFIFO/n1042 ,
         \u_outFIFO/n1041 , \u_outFIFO/n1040 , \u_outFIFO/n1039 ,
         \u_outFIFO/n1038 , \u_outFIFO/n1037 , \u_outFIFO/n1036 ,
         \u_outFIFO/n1035 , \u_outFIFO/n1034 , \u_outFIFO/n1033 ,
         \u_outFIFO/n1032 , \u_outFIFO/n1031 , \u_outFIFO/n1030 ,
         \u_outFIFO/n1029 , \u_outFIFO/n1028 , \u_outFIFO/n1027 ,
         \u_outFIFO/n1026 , \u_outFIFO/n1025 , \u_outFIFO/n1024 ,
         \u_outFIFO/n1023 , \u_outFIFO/n1022 , \u_outFIFO/n1021 ,
         \u_outFIFO/n1020 , \u_outFIFO/n1019 , \u_outFIFO/n1018 ,
         \u_outFIFO/n1017 , \u_outFIFO/n1016 , \u_outFIFO/n1015 ,
         \u_outFIFO/n1014 , \u_outFIFO/n1013 , \u_outFIFO/n1012 ,
         \u_outFIFO/n1011 , \u_outFIFO/n1010 , \u_outFIFO/n1009 ,
         \u_outFIFO/n1008 , \u_outFIFO/n1007 , \u_outFIFO/n1006 ,
         \u_outFIFO/n1005 , \u_outFIFO/n1004 , \u_outFIFO/n1003 ,
         \u_outFIFO/n1002 , \u_outFIFO/n1001 , \u_outFIFO/n1000 ,
         \u_outFIFO/n999 , \u_outFIFO/n998 , \u_outFIFO/n997 ,
         \u_outFIFO/n996 , \u_outFIFO/n995 , \u_outFIFO/n994 ,
         \u_outFIFO/n993 , \u_outFIFO/n992 , \u_outFIFO/n991 ,
         \u_outFIFO/n990 , \u_outFIFO/n989 , \u_outFIFO/n988 ,
         \u_outFIFO/n987 , \u_outFIFO/n986 , \u_outFIFO/n985 ,
         \u_outFIFO/n984 , \u_outFIFO/n983 , \u_outFIFO/n982 ,
         \u_outFIFO/n981 , \u_outFIFO/n980 , \u_outFIFO/n979 ,
         \u_outFIFO/n978 , \u_outFIFO/n977 , \u_outFIFO/n976 ,
         \u_outFIFO/n975 , \u_outFIFO/n974 , \u_outFIFO/n973 ,
         \u_outFIFO/n972 , \u_outFIFO/n971 , \u_outFIFO/n970 ,
         \u_outFIFO/n969 , \u_outFIFO/n968 , \u_outFIFO/n967 ,
         \u_outFIFO/n966 , \u_outFIFO/n965 , \u_outFIFO/n964 ,
         \u_outFIFO/n963 , \u_outFIFO/n962 , \u_outFIFO/n961 ,
         \u_outFIFO/n960 , \u_outFIFO/n959 , \u_outFIFO/n958 ,
         \u_outFIFO/n957 , \u_outFIFO/n956 , \u_outFIFO/n955 ,
         \u_outFIFO/n954 , \u_outFIFO/n953 , \u_outFIFO/n952 ,
         \u_outFIFO/n951 , \u_outFIFO/n950 , \u_outFIFO/n949 ,
         \u_outFIFO/n948 , \u_outFIFO/n947 , \u_outFIFO/n946 ,
         \u_outFIFO/n945 , \u_outFIFO/n944 , \u_outFIFO/n943 ,
         \u_outFIFO/n942 , \u_outFIFO/n941 , \u_outFIFO/n940 ,
         \u_outFIFO/n939 , \u_outFIFO/n938 , \u_outFIFO/n937 ,
         \u_outFIFO/n936 , \u_outFIFO/n935 , \u_outFIFO/n934 ,
         \u_outFIFO/n933 , \u_outFIFO/n932 , \u_outFIFO/n931 ,
         \u_outFIFO/n930 , \u_outFIFO/n929 , \u_outFIFO/n928 ,
         \u_outFIFO/n927 , \u_outFIFO/n926 , \u_outFIFO/n925 ,
         \u_outFIFO/n924 , \u_outFIFO/n923 , \u_outFIFO/n922 ,
         \u_outFIFO/n921 , \u_outFIFO/n920 , \u_outFIFO/n919 ,
         \u_outFIFO/n918 , \u_outFIFO/n917 , \u_outFIFO/n916 ,
         \u_outFIFO/n915 , \u_outFIFO/n914 , \u_outFIFO/n913 ,
         \u_outFIFO/n912 , \u_outFIFO/n911 , \u_outFIFO/n910 ,
         \u_outFIFO/n909 , \u_outFIFO/n908 , \u_outFIFO/n907 ,
         \u_outFIFO/n906 , \u_outFIFO/n905 , \u_outFIFO/n904 ,
         \u_outFIFO/n903 , \u_outFIFO/n902 , \u_outFIFO/n901 ,
         \u_outFIFO/n900 , \u_outFIFO/n899 , \u_outFIFO/n898 ,
         \u_outFIFO/n897 , \u_outFIFO/n896 , \u_outFIFO/n895 ,
         \u_outFIFO/n894 , \u_outFIFO/n893 , \u_outFIFO/n892 ,
         \u_outFIFO/n891 , \u_outFIFO/n890 , \u_outFIFO/n889 ,
         \u_outFIFO/n888 , \u_outFIFO/n887 , \u_outFIFO/n886 ,
         \u_outFIFO/n885 , \u_outFIFO/n884 , \u_outFIFO/n883 ,
         \u_outFIFO/n882 , \u_outFIFO/n881 , \u_outFIFO/n880 ,
         \u_outFIFO/n879 , \u_outFIFO/n878 , \u_outFIFO/n877 ,
         \u_outFIFO/n876 , \u_outFIFO/n875 , \u_outFIFO/n874 ,
         \u_outFIFO/n873 , \u_outFIFO/n872 , \u_outFIFO/n871 ,
         \u_outFIFO/n870 , \u_outFIFO/n869 , \u_outFIFO/n868 ,
         \u_outFIFO/n867 , \u_outFIFO/n866 , \u_outFIFO/n865 ,
         \u_outFIFO/n864 , \u_outFIFO/n863 , \u_outFIFO/n862 ,
         \u_outFIFO/n861 , \u_outFIFO/n860 , \u_outFIFO/n859 ,
         \u_outFIFO/n858 , \u_outFIFO/n857 , \u_outFIFO/n856 ,
         \u_outFIFO/n855 , \u_outFIFO/n854 , \u_outFIFO/n853 ,
         \u_outFIFO/n852 , \u_outFIFO/n851 , \u_outFIFO/n850 ,
         \u_outFIFO/n849 , \u_outFIFO/n848 , \u_outFIFO/n847 ,
         \u_outFIFO/n846 , \u_outFIFO/n845 , \u_outFIFO/n844 ,
         \u_outFIFO/n843 , \u_outFIFO/n842 , \u_outFIFO/n841 ,
         \u_outFIFO/n840 , \u_outFIFO/n839 , \u_outFIFO/n838 ,
         \u_outFIFO/n837 , \u_outFIFO/n836 , \u_outFIFO/n835 ,
         \u_outFIFO/n834 , \u_outFIFO/n833 , \u_outFIFO/n832 ,
         \u_outFIFO/n831 , \u_outFIFO/n830 , \u_outFIFO/n829 ,
         \u_outFIFO/n828 , \u_outFIFO/n827 , \u_outFIFO/n826 ,
         \u_outFIFO/n825 , \u_outFIFO/n824 , \u_outFIFO/n823 ,
         \u_outFIFO/n822 , \u_outFIFO/n821 , \u_outFIFO/n820 ,
         \u_outFIFO/n819 , \u_outFIFO/n818 , \u_outFIFO/n817 ,
         \u_outFIFO/n816 , \u_outFIFO/n815 , \u_outFIFO/n814 ,
         \u_outFIFO/n813 , \u_outFIFO/n812 , \u_outFIFO/n811 ,
         \u_outFIFO/n810 , \u_outFIFO/n809 , \u_outFIFO/n808 ,
         \u_outFIFO/n807 , \u_outFIFO/n806 , \u_outFIFO/n805 ,
         \u_outFIFO/n804 , \u_outFIFO/n803 , \u_outFIFO/n802 ,
         \u_outFIFO/n801 , \u_outFIFO/n800 , \u_outFIFO/n799 ,
         \u_outFIFO/n798 , \u_outFIFO/n797 , \u_outFIFO/n796 ,
         \u_outFIFO/n795 , \u_outFIFO/n794 , \u_outFIFO/n793 ,
         \u_outFIFO/n792 , \u_outFIFO/n791 , \u_outFIFO/n790 ,
         \u_outFIFO/n789 , \u_outFIFO/n788 , \u_outFIFO/n787 ,
         \u_outFIFO/n786 , \u_outFIFO/n785 , \u_outFIFO/n784 ,
         \u_outFIFO/n783 , \u_outFIFO/n782 , \u_outFIFO/n781 ,
         \u_outFIFO/n780 , \u_outFIFO/n779 , \u_outFIFO/n778 ,
         \u_outFIFO/n777 , \u_outFIFO/n776 , \u_outFIFO/n775 ,
         \u_outFIFO/n774 , \u_outFIFO/n773 , \u_outFIFO/n772 ,
         \u_outFIFO/n771 , \u_outFIFO/n770 , \u_outFIFO/n769 ,
         \u_outFIFO/n768 , \u_outFIFO/n767 , \u_outFIFO/n766 ,
         \u_outFIFO/n765 , \u_outFIFO/n764 , \u_outFIFO/n763 ,
         \u_outFIFO/n762 , \u_outFIFO/n761 , \u_outFIFO/n760 ,
         \u_outFIFO/n759 , \u_outFIFO/n758 , \u_outFIFO/n757 ,
         \u_outFIFO/n756 , \u_outFIFO/n755 , \u_outFIFO/n754 ,
         \u_outFIFO/n753 , \u_outFIFO/n752 , \u_outFIFO/n751 ,
         \u_outFIFO/n750 , \u_outFIFO/n749 , \u_outFIFO/n748 ,
         \u_outFIFO/n747 , \u_outFIFO/n746 , \u_outFIFO/n745 ,
         \u_outFIFO/n744 , \u_outFIFO/n743 , \u_outFIFO/n742 ,
         \u_outFIFO/n741 , \u_outFIFO/n740 , \u_outFIFO/n739 ,
         \u_outFIFO/n738 , \u_outFIFO/n737 , \u_outFIFO/n736 ,
         \u_outFIFO/n735 , \u_outFIFO/n734 , \u_outFIFO/n733 ,
         \u_outFIFO/n732 , \u_outFIFO/n731 , \u_outFIFO/n730 ,
         \u_outFIFO/n729 , \u_outFIFO/n728 , \u_outFIFO/n727 ,
         \u_outFIFO/n726 , \u_outFIFO/n725 , \u_outFIFO/n724 ,
         \u_outFIFO/n723 , \u_outFIFO/n722 , \u_outFIFO/n721 ,
         \u_outFIFO/n720 , \u_outFIFO/n719 , \u_outFIFO/n718 ,
         \u_outFIFO/n717 , \u_outFIFO/n716 , \u_outFIFO/n715 ,
         \u_outFIFO/n714 , \u_outFIFO/n713 , \u_outFIFO/n712 ,
         \u_outFIFO/n711 , \u_outFIFO/n710 , \u_outFIFO/n709 ,
         \u_outFIFO/n708 , \u_outFIFO/n707 , \u_outFIFO/n706 ,
         \u_outFIFO/n705 , \u_outFIFO/n704 , \u_outFIFO/n703 ,
         \u_outFIFO/n702 , \u_outFIFO/n701 , \u_outFIFO/n700 ,
         \u_outFIFO/n699 , \u_outFIFO/n698 , \u_outFIFO/n697 ,
         \u_outFIFO/n696 , \u_outFIFO/n695 , \u_outFIFO/n694 ,
         \u_outFIFO/n693 , \u_outFIFO/n692 , \u_outFIFO/n691 ,
         \u_outFIFO/n690 , \u_outFIFO/n689 , \u_outFIFO/n688 ,
         \u_outFIFO/n687 , \u_outFIFO/n686 , \u_outFIFO/n685 ,
         \u_outFIFO/n684 , \u_outFIFO/n683 , \u_outFIFO/n682 ,
         \u_outFIFO/n681 , \u_outFIFO/n680 , \u_outFIFO/n679 ,
         \u_outFIFO/n678 , \u_outFIFO/n677 , \u_outFIFO/n676 ,
         \u_outFIFO/n675 , \u_outFIFO/n674 , \u_outFIFO/n673 ,
         \u_outFIFO/n672 , \u_outFIFO/n671 , \u_outFIFO/n670 ,
         \u_outFIFO/n669 , \u_outFIFO/n668 , \u_outFIFO/n667 ,
         \u_outFIFO/n666 , \u_outFIFO/n665 , \u_outFIFO/n664 ,
         \u_outFIFO/n663 , \u_outFIFO/n662 , \u_outFIFO/n661 ,
         \u_outFIFO/n660 , \u_outFIFO/n659 , \u_outFIFO/n658 ,
         \u_outFIFO/n657 , \u_outFIFO/n656 , \u_outFIFO/n655 ,
         \u_outFIFO/n654 , \u_outFIFO/n653 , \u_outFIFO/n652 ,
         \u_outFIFO/n651 , \u_outFIFO/n650 , \u_outFIFO/n649 ,
         \u_outFIFO/n648 , \u_outFIFO/n647 , \u_outFIFO/n646 ,
         \u_outFIFO/n645 , \u_outFIFO/n644 , \u_outFIFO/n643 ,
         \u_outFIFO/n642 , \u_outFIFO/n641 , \u_outFIFO/n640 ,
         \u_outFIFO/n639 , \u_outFIFO/n638 , \u_outFIFO/n637 ,
         \u_outFIFO/n636 , \u_outFIFO/n635 , \u_outFIFO/n634 ,
         \u_outFIFO/n633 , \u_outFIFO/n632 , \u_outFIFO/n631 ,
         \u_outFIFO/n630 , \u_outFIFO/n629 , \u_outFIFO/n628 ,
         \u_outFIFO/n627 , \u_outFIFO/n626 , \u_outFIFO/n625 ,
         \u_outFIFO/n624 , \u_outFIFO/n623 , \u_outFIFO/n622 ,
         \u_outFIFO/n621 , \u_outFIFO/n620 , \u_outFIFO/n619 ,
         \u_outFIFO/n618 , \u_outFIFO/n617 , \u_outFIFO/n616 ,
         \u_outFIFO/n615 , \u_outFIFO/n614 , \u_outFIFO/n613 ,
         \u_outFIFO/n612 , \u_outFIFO/n611 , \u_outFIFO/n610 ,
         \u_outFIFO/n609 , \u_outFIFO/n608 , \u_outFIFO/n607 ,
         \u_outFIFO/n606 , \u_outFIFO/n605 , \u_outFIFO/n604 ,
         \u_outFIFO/n603 , \u_outFIFO/n602 , \u_outFIFO/n601 ,
         \u_outFIFO/n600 , \u_outFIFO/n599 , \u_outFIFO/n598 ,
         \u_outFIFO/n597 , \u_outFIFO/n596 , \u_outFIFO/n595 ,
         \u_outFIFO/n594 , \u_outFIFO/n593 , \u_outFIFO/n592 ,
         \u_outFIFO/n591 , \u_outFIFO/n590 , \u_outFIFO/n589 ,
         \u_outFIFO/n588 , \u_outFIFO/n587 , \u_outFIFO/n586 ,
         \u_outFIFO/n585 , \u_outFIFO/n584 , \u_outFIFO/n583 ,
         \u_outFIFO/n582 , \u_outFIFO/n581 , \u_outFIFO/n580 ,
         \u_outFIFO/n579 , \u_outFIFO/n578 , \u_outFIFO/n577 ,
         \u_outFIFO/n576 , \u_outFIFO/n575 , \u_outFIFO/n574 ,
         \u_outFIFO/n573 , \u_outFIFO/n572 , \u_outFIFO/n571 ,
         \u_outFIFO/n570 , \u_outFIFO/n569 , \u_outFIFO/n568 ,
         \u_outFIFO/n567 , \u_outFIFO/n566 , \u_outFIFO/n565 ,
         \u_outFIFO/n564 , \u_outFIFO/n563 , \u_outFIFO/n562 ,
         \u_outFIFO/n561 , \u_outFIFO/n560 , \u_outFIFO/n559 ,
         \u_outFIFO/n558 , \u_outFIFO/n557 , \u_outFIFO/n556 ,
         \u_outFIFO/n555 , \u_outFIFO/n554 , \u_outFIFO/n553 ,
         \u_outFIFO/n552 , \u_outFIFO/n551 , \u_outFIFO/n550 ,
         \u_outFIFO/n549 , \u_outFIFO/n548 , \u_outFIFO/n547 ,
         \u_outFIFO/n546 , \u_outFIFO/n545 , \u_outFIFO/n544 ,
         \u_outFIFO/n543 , \u_outFIFO/n542 , \u_outFIFO/n541 ,
         \u_outFIFO/n540 , \u_outFIFO/n539 , \u_outFIFO/n538 ,
         \u_outFIFO/n537 , \u_outFIFO/n536 , \u_outFIFO/n535 ,
         \u_outFIFO/n534 , \u_outFIFO/n533 , \u_outFIFO/n532 ,
         \u_outFIFO/n531 , \u_outFIFO/n530 , \u_outFIFO/n529 ,
         \u_outFIFO/n528 , \u_outFIFO/n527 , \u_outFIFO/n526 ,
         \u_outFIFO/n525 , \u_outFIFO/n524 , \u_outFIFO/n523 ,
         \u_outFIFO/n522 , \u_outFIFO/n521 , \u_outFIFO/n520 ,
         \u_outFIFO/n519 , \u_outFIFO/n518 , \u_outFIFO/n517 ,
         \u_outFIFO/n516 , \u_outFIFO/n515 , \u_outFIFO/n514 ,
         \u_outFIFO/n513 , \u_outFIFO/n512 , \u_outFIFO/n511 ,
         \u_outFIFO/n510 , \u_outFIFO/n509 , \u_outFIFO/n508 ,
         \u_outFIFO/n507 , \u_outFIFO/n506 , \u_outFIFO/n505 ,
         \u_outFIFO/n504 , \u_outFIFO/n503 , \u_outFIFO/n502 ,
         \u_outFIFO/n501 , \u_outFIFO/n500 , \u_outFIFO/n499 ,
         \u_outFIFO/n498 , \u_outFIFO/n497 , \u_outFIFO/n496 ,
         \u_outFIFO/n495 , \u_outFIFO/n494 , \u_outFIFO/n493 ,
         \u_outFIFO/n492 , \u_outFIFO/n491 , \u_outFIFO/n490 ,
         \u_outFIFO/n489 , \u_outFIFO/n488 , \u_outFIFO/n487 ,
         \u_outFIFO/n486 , \u_outFIFO/n485 , \u_outFIFO/n484 ,
         \u_outFIFO/n483 , \u_outFIFO/n482 , \u_outFIFO/n481 ,
         \u_outFIFO/n480 , \u_outFIFO/n479 , \u_outFIFO/n478 ,
         \u_outFIFO/n477 , \u_outFIFO/n476 , \u_outFIFO/n475 ,
         \u_outFIFO/n474 , \u_outFIFO/n473 , \u_outFIFO/n472 ,
         \u_outFIFO/n471 , \u_outFIFO/n470 , \u_outFIFO/n469 ,
         \u_outFIFO/n468 , \u_outFIFO/n467 , \u_outFIFO/n466 ,
         \u_outFIFO/n465 , \u_outFIFO/n464 , \u_outFIFO/n463 ,
         \u_outFIFO/n462 , \u_outFIFO/n461 , \u_outFIFO/n460 ,
         \u_outFIFO/n459 , \u_outFIFO/n458 , \u_outFIFO/n457 ,
         \u_outFIFO/n456 , \u_outFIFO/n455 , \u_outFIFO/n454 ,
         \u_outFIFO/n453 , \u_outFIFO/n452 , \u_outFIFO/n451 ,
         \u_outFIFO/n450 , \u_outFIFO/n449 , \u_outFIFO/n448 ,
         \u_outFIFO/n447 , \u_outFIFO/n446 , \u_outFIFO/n445 ,
         \u_outFIFO/n444 , \u_outFIFO/n443 , \u_outFIFO/n442 ,
         \u_outFIFO/n441 , \u_outFIFO/n440 , \u_outFIFO/n439 ,
         \u_outFIFO/n438 , \u_outFIFO/n437 , \u_outFIFO/n436 ,
         \u_outFIFO/n435 , \u_outFIFO/n434 , \u_outFIFO/n433 ,
         \u_outFIFO/n432 , \u_outFIFO/n431 , \u_outFIFO/n430 ,
         \u_outFIFO/n429 , \u_outFIFO/n428 , \u_outFIFO/n427 ,
         \u_outFIFO/n426 , \u_outFIFO/n425 , \u_outFIFO/n424 ,
         \u_outFIFO/n423 , \u_outFIFO/n422 , \u_outFIFO/n421 ,
         \u_outFIFO/n420 , \u_outFIFO/n419 , \u_outFIFO/n418 ,
         \u_outFIFO/n417 , \u_outFIFO/n416 , \u_outFIFO/n415 ,
         \u_outFIFO/n414 , \u_outFIFO/n413 , \u_outFIFO/n412 ,
         \u_outFIFO/n411 , \u_outFIFO/n410 , \u_outFIFO/n409 ,
         \u_outFIFO/n408 , \u_outFIFO/n407 , \u_outFIFO/n406 ,
         \u_outFIFO/n405 , \u_outFIFO/n404 , \u_outFIFO/n403 ,
         \u_outFIFO/n402 , \u_outFIFO/n401 , \u_outFIFO/n400 ,
         \u_outFIFO/n399 , \u_outFIFO/n398 , \u_outFIFO/n397 ,
         \u_outFIFO/n396 , \u_outFIFO/n395 , \u_outFIFO/n394 ,
         \u_outFIFO/n393 , \u_outFIFO/n392 , \u_outFIFO/n391 ,
         \u_outFIFO/n390 , \u_outFIFO/n389 , \u_outFIFO/n388 ,
         \u_outFIFO/n387 , \u_outFIFO/n386 , \u_outFIFO/n385 ,
         \u_outFIFO/n384 , \u_outFIFO/n383 , \u_outFIFO/n382 ,
         \u_outFIFO/n381 , \u_outFIFO/n380 , \u_outFIFO/n379 ,
         \u_outFIFO/n378 , \u_outFIFO/n377 , \u_outFIFO/n376 ,
         \u_outFIFO/n375 , \u_outFIFO/n374 , \u_outFIFO/n373 ,
         \u_outFIFO/n372 , \u_outFIFO/n371 , \u_outFIFO/n370 ,
         \u_outFIFO/n369 , \u_outFIFO/n368 , \u_outFIFO/n367 ,
         \u_outFIFO/n366 , \u_outFIFO/n365 , \u_outFIFO/n364 ,
         \u_outFIFO/n363 , \u_outFIFO/n362 , \u_outFIFO/n361 ,
         \u_outFIFO/n360 , \u_outFIFO/n359 , \u_outFIFO/n358 ,
         \u_outFIFO/n357 , \u_outFIFO/n356 , \u_outFIFO/n355 ,
         \u_outFIFO/n354 , \u_outFIFO/n353 , \u_outFIFO/n352 ,
         \u_outFIFO/n351 , \u_outFIFO/n350 , \u_outFIFO/n349 ,
         \u_outFIFO/n348 , \u_outFIFO/n347 , \u_outFIFO/n346 ,
         \u_outFIFO/n345 , \u_outFIFO/n344 , \u_outFIFO/n343 ,
         \u_outFIFO/n342 , \u_outFIFO/n341 , \u_outFIFO/n340 ,
         \u_outFIFO/n339 , \u_outFIFO/n338 , \u_outFIFO/n337 ,
         \u_outFIFO/n336 , \u_outFIFO/n335 , \u_outFIFO/n334 ,
         \u_outFIFO/n333 , \u_outFIFO/n332 , \u_outFIFO/n331 ,
         \u_outFIFO/n330 , \u_outFIFO/n329 , \u_outFIFO/n328 ,
         \u_outFIFO/n327 , \u_outFIFO/n326 , \u_outFIFO/n325 ,
         \u_outFIFO/n324 , \u_outFIFO/n323 , \u_outFIFO/n322 ,
         \u_outFIFO/n321 , \u_outFIFO/n320 , \u_outFIFO/n319 ,
         \u_outFIFO/n318 , \u_outFIFO/n317 , \u_outFIFO/n316 ,
         \u_outFIFO/n315 , \u_outFIFO/n314 , \u_outFIFO/n313 ,
         \u_outFIFO/n312 , \u_outFIFO/n311 , \u_outFIFO/n310 ,
         \u_outFIFO/n309 , \u_outFIFO/n308 , \u_outFIFO/n301 ,
         \u_outFIFO/n300 , \u_outFIFO/n299 , \u_outFIFO/n298 ,
         \u_outFIFO/n297 , \u_outFIFO/n296 , \u_outFIFO/n295 ,
         \u_outFIFO/n285 , \u_outFIFO/n284 , \u_outFIFO/n280 ,
         \u_outFIFO/n279 , \u_outFIFO/n278 , \u_outFIFO/n277 ,
         \u_outFIFO/n276 , \u_outFIFO/n275 , \u_outFIFO/n267 ,
         \u_outFIFO/n266 , \u_outFIFO/n265 , \u_outFIFO/n264 ,
         \u_outFIFO/n263 , \u_outFIFO/n262 , \u_outFIFO/n261 ,
         \u_outFIFO/n260 , \u_outFIFO/n258 , \u_outFIFO/n257 ,
         \u_outFIFO/n256 , \u_outFIFO/n254 , \u_outFIFO/n253 ,
         \u_outFIFO/N1270 , \u_outFIFO/N1269 , \u_outFIFO/N220 ,
         \u_outFIFO/N219 , \u_outFIFO/N218 , \u_outFIFO/N217 ,
         \u_outFIFO/N216 , \u_outFIFO/N205 , \u_outFIFO/N204 ,
         \u_outFIFO/N203 , \u_outFIFO/N202 , \u_outFIFO/FIFO[127][3] ,
         \u_outFIFO/FIFO[127][2] , \u_outFIFO/FIFO[127][1] ,
         \u_outFIFO/FIFO[127][0] , \u_outFIFO/FIFO[126][3] ,
         \u_outFIFO/FIFO[126][2] , \u_outFIFO/FIFO[126][1] ,
         \u_outFIFO/FIFO[126][0] , \u_outFIFO/FIFO[125][3] ,
         \u_outFIFO/FIFO[125][2] , \u_outFIFO/FIFO[125][1] ,
         \u_outFIFO/FIFO[125][0] , \u_outFIFO/FIFO[124][3] ,
         \u_outFIFO/FIFO[124][2] , \u_outFIFO/FIFO[124][1] ,
         \u_outFIFO/FIFO[124][0] , \u_outFIFO/FIFO[123][3] ,
         \u_outFIFO/FIFO[123][2] , \u_outFIFO/FIFO[123][1] ,
         \u_outFIFO/FIFO[123][0] , \u_outFIFO/FIFO[122][3] ,
         \u_outFIFO/FIFO[122][2] , \u_outFIFO/FIFO[122][1] ,
         \u_outFIFO/FIFO[122][0] , \u_outFIFO/FIFO[121][3] ,
         \u_outFIFO/FIFO[121][2] , \u_outFIFO/FIFO[121][1] ,
         \u_outFIFO/FIFO[121][0] , \u_outFIFO/FIFO[120][3] ,
         \u_outFIFO/FIFO[120][2] , \u_outFIFO/FIFO[120][1] ,
         \u_outFIFO/FIFO[120][0] , \u_outFIFO/FIFO[119][3] ,
         \u_outFIFO/FIFO[119][2] , \u_outFIFO/FIFO[119][1] ,
         \u_outFIFO/FIFO[119][0] , \u_outFIFO/FIFO[118][3] ,
         \u_outFIFO/FIFO[118][2] , \u_outFIFO/FIFO[118][1] ,
         \u_outFIFO/FIFO[118][0] , \u_outFIFO/FIFO[117][3] ,
         \u_outFIFO/FIFO[117][2] , \u_outFIFO/FIFO[117][1] ,
         \u_outFIFO/FIFO[117][0] , \u_outFIFO/FIFO[116][3] ,
         \u_outFIFO/FIFO[116][2] , \u_outFIFO/FIFO[116][1] ,
         \u_outFIFO/FIFO[116][0] , \u_outFIFO/FIFO[115][3] ,
         \u_outFIFO/FIFO[115][2] , \u_outFIFO/FIFO[115][1] ,
         \u_outFIFO/FIFO[115][0] , \u_outFIFO/FIFO[114][3] ,
         \u_outFIFO/FIFO[114][2] , \u_outFIFO/FIFO[114][1] ,
         \u_outFIFO/FIFO[114][0] , \u_outFIFO/FIFO[113][3] ,
         \u_outFIFO/FIFO[113][2] , \u_outFIFO/FIFO[113][1] ,
         \u_outFIFO/FIFO[113][0] , \u_outFIFO/FIFO[112][3] ,
         \u_outFIFO/FIFO[112][2] , \u_outFIFO/FIFO[112][1] ,
         \u_outFIFO/FIFO[112][0] , \u_outFIFO/FIFO[111][3] ,
         \u_outFIFO/FIFO[111][2] , \u_outFIFO/FIFO[111][1] ,
         \u_outFIFO/FIFO[111][0] , \u_outFIFO/FIFO[110][3] ,
         \u_outFIFO/FIFO[110][2] , \u_outFIFO/FIFO[110][1] ,
         \u_outFIFO/FIFO[110][0] , \u_outFIFO/FIFO[109][3] ,
         \u_outFIFO/FIFO[109][2] , \u_outFIFO/FIFO[109][1] ,
         \u_outFIFO/FIFO[109][0] , \u_outFIFO/FIFO[108][3] ,
         \u_outFIFO/FIFO[108][2] , \u_outFIFO/FIFO[108][1] ,
         \u_outFIFO/FIFO[108][0] , \u_outFIFO/FIFO[107][3] ,
         \u_outFIFO/FIFO[107][2] , \u_outFIFO/FIFO[107][1] ,
         \u_outFIFO/FIFO[107][0] , \u_outFIFO/FIFO[106][3] ,
         \u_outFIFO/FIFO[106][2] , \u_outFIFO/FIFO[106][1] ,
         \u_outFIFO/FIFO[106][0] , \u_outFIFO/FIFO[105][3] ,
         \u_outFIFO/FIFO[105][2] , \u_outFIFO/FIFO[105][1] ,
         \u_outFIFO/FIFO[105][0] , \u_outFIFO/FIFO[104][3] ,
         \u_outFIFO/FIFO[104][2] , \u_outFIFO/FIFO[104][1] ,
         \u_outFIFO/FIFO[104][0] , \u_outFIFO/FIFO[103][3] ,
         \u_outFIFO/FIFO[103][2] , \u_outFIFO/FIFO[103][1] ,
         \u_outFIFO/FIFO[103][0] , \u_outFIFO/FIFO[102][3] ,
         \u_outFIFO/FIFO[102][2] , \u_outFIFO/FIFO[102][1] ,
         \u_outFIFO/FIFO[102][0] , \u_outFIFO/FIFO[101][3] ,
         \u_outFIFO/FIFO[101][2] , \u_outFIFO/FIFO[101][1] ,
         \u_outFIFO/FIFO[101][0] , \u_outFIFO/FIFO[100][3] ,
         \u_outFIFO/FIFO[100][2] , \u_outFIFO/FIFO[100][1] ,
         \u_outFIFO/FIFO[100][0] , \u_outFIFO/FIFO[99][3] ,
         \u_outFIFO/FIFO[99][2] , \u_outFIFO/FIFO[99][1] ,
         \u_outFIFO/FIFO[99][0] , \u_outFIFO/FIFO[98][3] ,
         \u_outFIFO/FIFO[98][2] , \u_outFIFO/FIFO[98][1] ,
         \u_outFIFO/FIFO[98][0] , \u_outFIFO/FIFO[97][3] ,
         \u_outFIFO/FIFO[97][2] , \u_outFIFO/FIFO[97][1] ,
         \u_outFIFO/FIFO[97][0] , \u_outFIFO/FIFO[96][3] ,
         \u_outFIFO/FIFO[96][2] , \u_outFIFO/FIFO[96][1] ,
         \u_outFIFO/FIFO[96][0] , \u_outFIFO/FIFO[95][3] ,
         \u_outFIFO/FIFO[95][2] , \u_outFIFO/FIFO[95][1] ,
         \u_outFIFO/FIFO[95][0] , \u_outFIFO/FIFO[94][3] ,
         \u_outFIFO/FIFO[94][2] , \u_outFIFO/FIFO[94][1] ,
         \u_outFIFO/FIFO[94][0] , \u_outFIFO/FIFO[93][3] ,
         \u_outFIFO/FIFO[93][2] , \u_outFIFO/FIFO[93][1] ,
         \u_outFIFO/FIFO[93][0] , \u_outFIFO/FIFO[92][3] ,
         \u_outFIFO/FIFO[92][2] , \u_outFIFO/FIFO[92][1] ,
         \u_outFIFO/FIFO[92][0] , \u_outFIFO/FIFO[91][3] ,
         \u_outFIFO/FIFO[91][2] , \u_outFIFO/FIFO[91][1] ,
         \u_outFIFO/FIFO[91][0] , \u_outFIFO/FIFO[90][3] ,
         \u_outFIFO/FIFO[90][2] , \u_outFIFO/FIFO[90][1] ,
         \u_outFIFO/FIFO[90][0] , \u_outFIFO/FIFO[89][3] ,
         \u_outFIFO/FIFO[89][2] , \u_outFIFO/FIFO[89][1] ,
         \u_outFIFO/FIFO[89][0] , \u_outFIFO/FIFO[88][3] ,
         \u_outFIFO/FIFO[88][2] , \u_outFIFO/FIFO[88][1] ,
         \u_outFIFO/FIFO[88][0] , \u_outFIFO/FIFO[87][3] ,
         \u_outFIFO/FIFO[87][2] , \u_outFIFO/FIFO[87][1] ,
         \u_outFIFO/FIFO[87][0] , \u_outFIFO/FIFO[86][3] ,
         \u_outFIFO/FIFO[86][2] , \u_outFIFO/FIFO[86][1] ,
         \u_outFIFO/FIFO[86][0] , \u_outFIFO/FIFO[85][3] ,
         \u_outFIFO/FIFO[85][2] , \u_outFIFO/FIFO[85][1] ,
         \u_outFIFO/FIFO[85][0] , \u_outFIFO/FIFO[84][3] ,
         \u_outFIFO/FIFO[84][2] , \u_outFIFO/FIFO[84][1] ,
         \u_outFIFO/FIFO[84][0] , \u_outFIFO/FIFO[83][3] ,
         \u_outFIFO/FIFO[83][2] , \u_outFIFO/FIFO[83][1] ,
         \u_outFIFO/FIFO[83][0] , \u_outFIFO/FIFO[82][3] ,
         \u_outFIFO/FIFO[82][2] , \u_outFIFO/FIFO[82][1] ,
         \u_outFIFO/FIFO[82][0] , \u_outFIFO/FIFO[81][3] ,
         \u_outFIFO/FIFO[81][2] , \u_outFIFO/FIFO[81][1] ,
         \u_outFIFO/FIFO[81][0] , \u_outFIFO/FIFO[80][3] ,
         \u_outFIFO/FIFO[80][2] , \u_outFIFO/FIFO[80][1] ,
         \u_outFIFO/FIFO[80][0] , \u_outFIFO/FIFO[79][3] ,
         \u_outFIFO/FIFO[79][2] , \u_outFIFO/FIFO[79][1] ,
         \u_outFIFO/FIFO[79][0] , \u_outFIFO/FIFO[78][3] ,
         \u_outFIFO/FIFO[78][2] , \u_outFIFO/FIFO[78][1] ,
         \u_outFIFO/FIFO[78][0] , \u_outFIFO/FIFO[77][3] ,
         \u_outFIFO/FIFO[77][2] , \u_outFIFO/FIFO[77][1] ,
         \u_outFIFO/FIFO[77][0] , \u_outFIFO/FIFO[76][3] ,
         \u_outFIFO/FIFO[76][2] , \u_outFIFO/FIFO[76][1] ,
         \u_outFIFO/FIFO[76][0] , \u_outFIFO/FIFO[75][3] ,
         \u_outFIFO/FIFO[75][2] , \u_outFIFO/FIFO[75][1] ,
         \u_outFIFO/FIFO[75][0] , \u_outFIFO/FIFO[74][3] ,
         \u_outFIFO/FIFO[74][2] , \u_outFIFO/FIFO[74][1] ,
         \u_outFIFO/FIFO[74][0] , \u_outFIFO/FIFO[73][3] ,
         \u_outFIFO/FIFO[73][2] , \u_outFIFO/FIFO[73][1] ,
         \u_outFIFO/FIFO[73][0] , \u_outFIFO/FIFO[72][3] ,
         \u_outFIFO/FIFO[72][2] , \u_outFIFO/FIFO[72][1] ,
         \u_outFIFO/FIFO[72][0] , \u_outFIFO/FIFO[71][3] ,
         \u_outFIFO/FIFO[71][2] , \u_outFIFO/FIFO[71][1] ,
         \u_outFIFO/FIFO[71][0] , \u_outFIFO/FIFO[70][3] ,
         \u_outFIFO/FIFO[70][2] , \u_outFIFO/FIFO[70][1] ,
         \u_outFIFO/FIFO[70][0] , \u_outFIFO/FIFO[69][3] ,
         \u_outFIFO/FIFO[69][2] , \u_outFIFO/FIFO[69][1] ,
         \u_outFIFO/FIFO[69][0] , \u_outFIFO/FIFO[68][3] ,
         \u_outFIFO/FIFO[68][2] , \u_outFIFO/FIFO[68][1] ,
         \u_outFIFO/FIFO[68][0] , \u_outFIFO/FIFO[67][3] ,
         \u_outFIFO/FIFO[67][2] , \u_outFIFO/FIFO[67][1] ,
         \u_outFIFO/FIFO[67][0] , \u_outFIFO/FIFO[66][3] ,
         \u_outFIFO/FIFO[66][2] , \u_outFIFO/FIFO[66][1] ,
         \u_outFIFO/FIFO[66][0] , \u_outFIFO/FIFO[65][3] ,
         \u_outFIFO/FIFO[65][2] , \u_outFIFO/FIFO[65][1] ,
         \u_outFIFO/FIFO[65][0] , \u_outFIFO/FIFO[64][3] ,
         \u_outFIFO/FIFO[64][2] , \u_outFIFO/FIFO[64][1] ,
         \u_outFIFO/FIFO[64][0] , \u_outFIFO/FIFO[63][3] ,
         \u_outFIFO/FIFO[63][2] , \u_outFIFO/FIFO[63][1] ,
         \u_outFIFO/FIFO[63][0] , \u_outFIFO/FIFO[62][3] ,
         \u_outFIFO/FIFO[62][2] , \u_outFIFO/FIFO[62][1] ,
         \u_outFIFO/FIFO[62][0] , \u_outFIFO/FIFO[61][3] ,
         \u_outFIFO/FIFO[61][2] , \u_outFIFO/FIFO[61][1] ,
         \u_outFIFO/FIFO[61][0] , \u_outFIFO/FIFO[60][3] ,
         \u_outFIFO/FIFO[60][2] , \u_outFIFO/FIFO[60][1] ,
         \u_outFIFO/FIFO[60][0] , \u_outFIFO/FIFO[59][3] ,
         \u_outFIFO/FIFO[59][2] , \u_outFIFO/FIFO[59][1] ,
         \u_outFIFO/FIFO[59][0] , \u_outFIFO/FIFO[58][3] ,
         \u_outFIFO/FIFO[58][2] , \u_outFIFO/FIFO[58][1] ,
         \u_outFIFO/FIFO[58][0] , \u_outFIFO/FIFO[57][3] ,
         \u_outFIFO/FIFO[57][2] , \u_outFIFO/FIFO[57][1] ,
         \u_outFIFO/FIFO[57][0] , \u_outFIFO/FIFO[56][3] ,
         \u_outFIFO/FIFO[56][2] , \u_outFIFO/FIFO[56][1] ,
         \u_outFIFO/FIFO[56][0] , \u_outFIFO/FIFO[55][3] ,
         \u_outFIFO/FIFO[55][2] , \u_outFIFO/FIFO[55][1] ,
         \u_outFIFO/FIFO[55][0] , \u_outFIFO/FIFO[54][3] ,
         \u_outFIFO/FIFO[54][2] , \u_outFIFO/FIFO[54][1] ,
         \u_outFIFO/FIFO[54][0] , \u_outFIFO/FIFO[53][3] ,
         \u_outFIFO/FIFO[53][2] , \u_outFIFO/FIFO[53][1] ,
         \u_outFIFO/FIFO[53][0] , \u_outFIFO/FIFO[52][3] ,
         \u_outFIFO/FIFO[52][2] , \u_outFIFO/FIFO[52][1] ,
         \u_outFIFO/FIFO[52][0] , \u_outFIFO/FIFO[51][3] ,
         \u_outFIFO/FIFO[51][2] , \u_outFIFO/FIFO[51][1] ,
         \u_outFIFO/FIFO[51][0] , \u_outFIFO/FIFO[50][3] ,
         \u_outFIFO/FIFO[50][2] , \u_outFIFO/FIFO[50][1] ,
         \u_outFIFO/FIFO[50][0] , \u_outFIFO/FIFO[49][3] ,
         \u_outFIFO/FIFO[49][2] , \u_outFIFO/FIFO[49][1] ,
         \u_outFIFO/FIFO[49][0] , \u_outFIFO/FIFO[48][3] ,
         \u_outFIFO/FIFO[48][2] , \u_outFIFO/FIFO[48][1] ,
         \u_outFIFO/FIFO[48][0] , \u_outFIFO/FIFO[47][3] ,
         \u_outFIFO/FIFO[47][2] , \u_outFIFO/FIFO[47][1] ,
         \u_outFIFO/FIFO[47][0] , \u_outFIFO/FIFO[46][3] ,
         \u_outFIFO/FIFO[46][2] , \u_outFIFO/FIFO[46][1] ,
         \u_outFIFO/FIFO[46][0] , \u_outFIFO/FIFO[45][3] ,
         \u_outFIFO/FIFO[45][2] , \u_outFIFO/FIFO[45][1] ,
         \u_outFIFO/FIFO[45][0] , \u_outFIFO/FIFO[44][3] ,
         \u_outFIFO/FIFO[44][2] , \u_outFIFO/FIFO[44][1] ,
         \u_outFIFO/FIFO[44][0] , \u_outFIFO/FIFO[43][3] ,
         \u_outFIFO/FIFO[43][2] , \u_outFIFO/FIFO[43][1] ,
         \u_outFIFO/FIFO[43][0] , \u_outFIFO/FIFO[42][3] ,
         \u_outFIFO/FIFO[42][2] , \u_outFIFO/FIFO[42][1] ,
         \u_outFIFO/FIFO[42][0] , \u_outFIFO/FIFO[41][3] ,
         \u_outFIFO/FIFO[41][2] , \u_outFIFO/FIFO[41][1] ,
         \u_outFIFO/FIFO[41][0] , \u_outFIFO/FIFO[40][3] ,
         \u_outFIFO/FIFO[40][2] , \u_outFIFO/FIFO[40][1] ,
         \u_outFIFO/FIFO[40][0] , \u_outFIFO/FIFO[39][3] ,
         \u_outFIFO/FIFO[39][2] , \u_outFIFO/FIFO[39][1] ,
         \u_outFIFO/FIFO[39][0] , \u_outFIFO/FIFO[38][3] ,
         \u_outFIFO/FIFO[38][2] , \u_outFIFO/FIFO[38][1] ,
         \u_outFIFO/FIFO[38][0] , \u_outFIFO/FIFO[37][3] ,
         \u_outFIFO/FIFO[37][2] , \u_outFIFO/FIFO[37][1] ,
         \u_outFIFO/FIFO[37][0] , \u_outFIFO/FIFO[36][3] ,
         \u_outFIFO/FIFO[36][2] , \u_outFIFO/FIFO[36][1] ,
         \u_outFIFO/FIFO[36][0] , \u_outFIFO/FIFO[35][3] ,
         \u_outFIFO/FIFO[35][2] , \u_outFIFO/FIFO[35][1] ,
         \u_outFIFO/FIFO[35][0] , \u_outFIFO/FIFO[34][3] ,
         \u_outFIFO/FIFO[34][2] , \u_outFIFO/FIFO[34][1] ,
         \u_outFIFO/FIFO[34][0] , \u_outFIFO/FIFO[33][3] ,
         \u_outFIFO/FIFO[33][2] , \u_outFIFO/FIFO[33][1] ,
         \u_outFIFO/FIFO[33][0] , \u_outFIFO/FIFO[32][3] ,
         \u_outFIFO/FIFO[32][2] , \u_outFIFO/FIFO[32][1] ,
         \u_outFIFO/FIFO[32][0] , \u_outFIFO/FIFO[31][3] ,
         \u_outFIFO/FIFO[31][2] , \u_outFIFO/FIFO[31][1] ,
         \u_outFIFO/FIFO[31][0] , \u_outFIFO/FIFO[30][3] ,
         \u_outFIFO/FIFO[30][2] , \u_outFIFO/FIFO[30][1] ,
         \u_outFIFO/FIFO[30][0] , \u_outFIFO/FIFO[29][3] ,
         \u_outFIFO/FIFO[29][2] , \u_outFIFO/FIFO[29][1] ,
         \u_outFIFO/FIFO[29][0] , \u_outFIFO/FIFO[28][3] ,
         \u_outFIFO/FIFO[28][2] , \u_outFIFO/FIFO[28][1] ,
         \u_outFIFO/FIFO[28][0] , \u_outFIFO/FIFO[27][3] ,
         \u_outFIFO/FIFO[27][2] , \u_outFIFO/FIFO[27][1] ,
         \u_outFIFO/FIFO[27][0] , \u_outFIFO/FIFO[26][3] ,
         \u_outFIFO/FIFO[26][2] , \u_outFIFO/FIFO[26][1] ,
         \u_outFIFO/FIFO[26][0] , \u_outFIFO/FIFO[25][3] ,
         \u_outFIFO/FIFO[25][2] , \u_outFIFO/FIFO[25][1] ,
         \u_outFIFO/FIFO[25][0] , \u_outFIFO/FIFO[24][3] ,
         \u_outFIFO/FIFO[24][2] , \u_outFIFO/FIFO[24][1] ,
         \u_outFIFO/FIFO[24][0] , \u_outFIFO/FIFO[23][3] ,
         \u_outFIFO/FIFO[23][2] , \u_outFIFO/FIFO[23][1] ,
         \u_outFIFO/FIFO[23][0] , \u_outFIFO/FIFO[22][3] ,
         \u_outFIFO/FIFO[22][2] , \u_outFIFO/FIFO[22][1] ,
         \u_outFIFO/FIFO[22][0] , \u_outFIFO/FIFO[21][3] ,
         \u_outFIFO/FIFO[21][2] , \u_outFIFO/FIFO[21][1] ,
         \u_outFIFO/FIFO[21][0] , \u_outFIFO/FIFO[20][3] ,
         \u_outFIFO/FIFO[20][2] , \u_outFIFO/FIFO[20][1] ,
         \u_outFIFO/FIFO[20][0] , \u_outFIFO/FIFO[19][3] ,
         \u_outFIFO/FIFO[19][2] , \u_outFIFO/FIFO[19][1] ,
         \u_outFIFO/FIFO[19][0] , \u_outFIFO/FIFO[18][3] ,
         \u_outFIFO/FIFO[18][2] , \u_outFIFO/FIFO[18][1] ,
         \u_outFIFO/FIFO[18][0] , \u_outFIFO/FIFO[17][3] ,
         \u_outFIFO/FIFO[17][2] , \u_outFIFO/FIFO[17][1] ,
         \u_outFIFO/FIFO[17][0] , \u_outFIFO/FIFO[16][3] ,
         \u_outFIFO/FIFO[16][2] , \u_outFIFO/FIFO[16][1] ,
         \u_outFIFO/FIFO[16][0] , \u_outFIFO/FIFO[15][3] ,
         \u_outFIFO/FIFO[15][2] , \u_outFIFO/FIFO[15][1] ,
         \u_outFIFO/FIFO[15][0] , \u_outFIFO/FIFO[14][3] ,
         \u_outFIFO/FIFO[14][2] , \u_outFIFO/FIFO[14][1] ,
         \u_outFIFO/FIFO[14][0] , \u_outFIFO/FIFO[13][3] ,
         \u_outFIFO/FIFO[13][2] , \u_outFIFO/FIFO[13][1] ,
         \u_outFIFO/FIFO[13][0] , \u_outFIFO/FIFO[12][3] ,
         \u_outFIFO/FIFO[12][2] , \u_outFIFO/FIFO[12][1] ,
         \u_outFIFO/FIFO[12][0] , \u_outFIFO/FIFO[11][3] ,
         \u_outFIFO/FIFO[11][2] , \u_outFIFO/FIFO[11][1] ,
         \u_outFIFO/FIFO[11][0] , \u_outFIFO/FIFO[10][3] ,
         \u_outFIFO/FIFO[10][2] , \u_outFIFO/FIFO[10][1] ,
         \u_outFIFO/FIFO[10][0] , \u_outFIFO/FIFO[9][3] ,
         \u_outFIFO/FIFO[9][2] , \u_outFIFO/FIFO[9][1] ,
         \u_outFIFO/FIFO[9][0] , \u_outFIFO/FIFO[8][3] ,
         \u_outFIFO/FIFO[8][2] , \u_outFIFO/FIFO[8][1] ,
         \u_outFIFO/FIFO[8][0] , \u_outFIFO/FIFO[7][3] ,
         \u_outFIFO/FIFO[7][2] , \u_outFIFO/FIFO[7][1] ,
         \u_outFIFO/FIFO[7][0] , \u_outFIFO/FIFO[6][3] ,
         \u_outFIFO/FIFO[6][2] , \u_outFIFO/FIFO[6][1] ,
         \u_outFIFO/FIFO[6][0] , \u_outFIFO/FIFO[5][3] ,
         \u_outFIFO/FIFO[5][2] , \u_outFIFO/FIFO[5][1] ,
         \u_outFIFO/FIFO[5][0] , \u_outFIFO/FIFO[4][3] ,
         \u_outFIFO/FIFO[4][2] , \u_outFIFO/FIFO[4][1] ,
         \u_outFIFO/FIFO[4][0] , \u_outFIFO/FIFO[3][3] ,
         \u_outFIFO/FIFO[3][2] , \u_outFIFO/FIFO[3][1] ,
         \u_outFIFO/FIFO[3][0] , \u_outFIFO/FIFO[2][3] ,
         \u_outFIFO/FIFO[2][2] , \u_outFIFO/FIFO[2][1] ,
         \u_outFIFO/FIFO[2][0] , \u_outFIFO/FIFO[1][3] ,
         \u_outFIFO/FIFO[1][2] , \u_outFIFO/FIFO[1][1] ,
         \u_outFIFO/FIFO[1][0] , \u_outFIFO/FIFO[0][3] ,
         \u_outFIFO/FIFO[0][2] , \u_outFIFO/FIFO[0][1] ,
         \u_outFIFO/FIFO[0][0] , \u_outFIFO/N198 , \u_outFIFO/N150 ,
         \u_outFIFO/N149 , \u_outFIFO/N148 , \u_outFIFO/N147 ,
         \u_outFIFO/N146 , \u_outFIFO/N145 , \u_outFIFO/N144 ,
         \u_outFIFO/N143 , \u_outFIFO/N141 , \u_outFIFO/N140 ,
         \u_outFIFO/N139 , \u_outFIFO/N138 , \u_outFIFO/N137 ,
         \u_outFIFO/N136 , \u_outFIFO/N132 , \u_outFIFO/N131 ,
         \u_outFIFO/N130 , \u_outFIFO/N129 , \u_outFIFO/N128 ,
         \u_outFIFO/N126 , \u_outFIFO/N125 , \u_outFIFO/N124 ,
         \u_outFIFO/N123 , \u_outFIFO/N122 , \u_outFIFO/N121 ,
         \u_outFIFO/N120 , \u_outFIFO/sigEnableCounter , \u_outFIFO/N50 ,
         \u_outFIFO/N49 , \u_outFIFO/N48 , \u_outFIFO/N47 ,
         \u_outFIFO/sig_fsm_start_W , \u_outFIFO/sig_fsm_start_R ,
         \u_outFIFO/outReadCount[0] , \u_outFIFO/outReadCount[1] ,
         \u_outFIFO/outReadCount[2] , \u_outFIFO/outReadCount[3] ,
         \u_outFIFO/outReadCount[4] , \u_outFIFO/outReadCount[5] ,
         \u_outFIFO/outReadCount[6] , \u_outFIFO/outWriteCount[0] ,
         \u_outFIFO/outWriteCount[1] , \u_outFIFO/outWriteCount[2] ,
         \u_outFIFO/outWriteCount[3] , \u_outFIFO/outWriteCount[4] ,
         \u_outFIFO/outWriteCount[5] , \u_outFIFO/outWriteCount[6] ,
         \u_outFIFO/outWriteCount[7] , \u_outFIFO/N45 , \u_outFIFO/N44 ,
         \u_outFIFO/N43 , \u_outFIFO/N42 , \u_outFIFO/N40 , \u_outFIFO/N39 ,
         \u_demux1/n5 , \u_demux1/n4 , \u_mux3/n3 , \u_mux8/n4 , \u_mux8/n3 ,
         \u_inFIFO/os1/sigQout2 , \u_inFIFO/os1/sigQout1 ,
         \u_decoder/iq_demod/n71 , \u_decoder/iq_demod/n70 ,
         \u_decoder/iq_demod/n69 , \u_decoder/iq_demod/n68 ,
         \u_decoder/iq_demod/n67 , \u_decoder/iq_demod/n66 ,
         \u_decoder/iq_demod/n65 , \u_decoder/iq_demod/n64 ,
         \u_decoder/iq_demod/n63 , \u_decoder/iq_demod/n62 ,
         \u_decoder/iq_demod/n61 , \u_decoder/iq_demod/n60 ,
         \u_decoder/iq_demod/n59 , \u_decoder/iq_demod/n58 ,
         \u_decoder/iq_demod/n57 , \u_decoder/iq_demod/n56 ,
         \u_decoder/iq_demod/n55 , \u_decoder/iq_demod/n54 ,
         \u_decoder/iq_demod/n53 , \u_decoder/iq_demod/n52 ,
         \u_decoder/iq_demod/n51 , \u_decoder/iq_demod/n50 ,
         \u_decoder/iq_demod/n49 , \u_decoder/iq_demod/n48 ,
         \u_decoder/iq_demod/n47 , \u_decoder/iq_demod/n46 ,
         \u_decoder/iq_demod/n45 , \u_decoder/iq_demod/n44 ,
         \u_decoder/iq_demod/n43 , \u_decoder/iq_demod/n42 ,
         \u_decoder/iq_demod/n41 , \u_decoder/iq_demod/n30 ,
         \u_decoder/iq_demod/I_if_buff[3] , \u_decoder/iq_demod/Q_if_buff[3] ,
         \u_decoder/iq_demod/N13 , \u_decoder/fir_filter/n1451 ,
         \u_decoder/fir_filter/n1450 , \u_decoder/fir_filter/n1449 ,
         \u_decoder/fir_filter/n1448 , \u_decoder/fir_filter/n1447 ,
         \u_decoder/fir_filter/n1446 , \u_decoder/fir_filter/n1445 ,
         \u_decoder/fir_filter/n1444 , \u_decoder/fir_filter/n1443 ,
         \u_decoder/fir_filter/n1442 , \u_decoder/fir_filter/n1441 ,
         \u_decoder/fir_filter/n1440 , \u_decoder/fir_filter/n1439 ,
         \u_decoder/fir_filter/n1438 , \u_decoder/fir_filter/n1437 ,
         \u_decoder/fir_filter/n1436 , \u_decoder/fir_filter/n1434 ,
         \u_decoder/fir_filter/n1433 , \u_decoder/fir_filter/n1432 ,
         \u_decoder/fir_filter/n1431 , \u_decoder/fir_filter/n1430 ,
         \u_decoder/fir_filter/n1429 , \u_decoder/fir_filter/n1428 ,
         \u_decoder/fir_filter/n1427 , \u_decoder/fir_filter/n1426 ,
         \u_decoder/fir_filter/n1425 , \u_decoder/fir_filter/n1424 ,
         \u_decoder/fir_filter/n1423 , \u_decoder/fir_filter/n1422 ,
         \u_decoder/fir_filter/n1421 , \u_decoder/fir_filter/n1420 ,
         \u_decoder/fir_filter/n1418 , \u_decoder/fir_filter/n1417 ,
         \u_decoder/fir_filter/n1416 , \u_decoder/fir_filter/n1415 ,
         \u_decoder/fir_filter/n1414 , \u_decoder/fir_filter/n1413 ,
         \u_decoder/fir_filter/n1412 , \u_decoder/fir_filter/n1411 ,
         \u_decoder/fir_filter/n1410 , \u_decoder/fir_filter/n1409 ,
         \u_decoder/fir_filter/n1408 , \u_decoder/fir_filter/n1407 ,
         \u_decoder/fir_filter/n1406 , \u_decoder/fir_filter/n1405 ,
         \u_decoder/fir_filter/n1402 , \u_decoder/fir_filter/n1401 ,
         \u_decoder/fir_filter/n1400 , \u_decoder/fir_filter/n1399 ,
         \u_decoder/fir_filter/n1398 , \u_decoder/fir_filter/n1397 ,
         \u_decoder/fir_filter/n1396 , \u_decoder/fir_filter/n1395 ,
         \u_decoder/fir_filter/n1394 , \u_decoder/fir_filter/n1393 ,
         \u_decoder/fir_filter/n1392 , \u_decoder/fir_filter/n1391 ,
         \u_decoder/fir_filter/n1390 , \u_decoder/fir_filter/n1389 ,
         \u_decoder/fir_filter/n1388 , \u_decoder/fir_filter/n1386 ,
         \u_decoder/fir_filter/n1385 , \u_decoder/fir_filter/n1384 ,
         \u_decoder/fir_filter/n1383 , \u_decoder/fir_filter/n1382 ,
         \u_decoder/fir_filter/n1381 , \u_decoder/fir_filter/n1380 ,
         \u_decoder/fir_filter/n1379 , \u_decoder/fir_filter/n1378 ,
         \u_decoder/fir_filter/n1377 , \u_decoder/fir_filter/n1376 ,
         \u_decoder/fir_filter/n1375 , \u_decoder/fir_filter/n1374 ,
         \u_decoder/fir_filter/n1373 , \u_decoder/fir_filter/n1372 ,
         \u_decoder/fir_filter/n1370 , \u_decoder/fir_filter/n1369 ,
         \u_decoder/fir_filter/n1368 , \u_decoder/fir_filter/n1367 ,
         \u_decoder/fir_filter/n1366 , \u_decoder/fir_filter/n1365 ,
         \u_decoder/fir_filter/n1364 , \u_decoder/fir_filter/n1363 ,
         \u_decoder/fir_filter/n1362 , \u_decoder/fir_filter/n1361 ,
         \u_decoder/fir_filter/n1360 , \u_decoder/fir_filter/n1359 ,
         \u_decoder/fir_filter/n1358 , \u_decoder/fir_filter/n1357 ,
         \u_decoder/fir_filter/n1354 , \u_decoder/fir_filter/n1353 ,
         \u_decoder/fir_filter/n1352 , \u_decoder/fir_filter/n1351 ,
         \u_decoder/fir_filter/n1350 , \u_decoder/fir_filter/n1349 ,
         \u_decoder/fir_filter/n1348 , \u_decoder/fir_filter/n1347 ,
         \u_decoder/fir_filter/n1346 , \u_decoder/fir_filter/n1345 ,
         \u_decoder/fir_filter/n1344 , \u_decoder/fir_filter/n1343 ,
         \u_decoder/fir_filter/n1342 , \u_decoder/fir_filter/n1341 ,
         \u_decoder/fir_filter/n1340 , \u_decoder/fir_filter/n1338 ,
         \u_decoder/fir_filter/n1337 , \u_decoder/fir_filter/n1336 ,
         \u_decoder/fir_filter/n1335 , \u_decoder/fir_filter/n1334 ,
         \u_decoder/fir_filter/n1333 , \u_decoder/fir_filter/n1332 ,
         \u_decoder/fir_filter/n1331 , \u_decoder/fir_filter/n1330 ,
         \u_decoder/fir_filter/n1329 , \u_decoder/fir_filter/n1328 ,
         \u_decoder/fir_filter/n1327 , \u_decoder/fir_filter/n1326 ,
         \u_decoder/fir_filter/n1325 , \u_decoder/fir_filter/n1324 ,
         \u_decoder/fir_filter/n1317 , \u_decoder/fir_filter/n1316 ,
         \u_decoder/fir_filter/n1315 , \u_decoder/fir_filter/n1314 ,
         \u_decoder/fir_filter/n1313 , \u_decoder/fir_filter/n1312 ,
         \u_decoder/fir_filter/n1311 , \u_decoder/fir_filter/n1310 ,
         \u_decoder/fir_filter/n1309 , \u_decoder/fir_filter/n1308 ,
         \u_decoder/fir_filter/n1307 , \u_decoder/fir_filter/n1306 ,
         \u_decoder/fir_filter/n1305 , \u_decoder/fir_filter/n1304 ,
         \u_decoder/fir_filter/n1303 , \u_decoder/fir_filter/n1302 ,
         \u_decoder/fir_filter/n1301 , \u_decoder/fir_filter/n1300 ,
         \u_decoder/fir_filter/n1299 , \u_decoder/fir_filter/n1298 ,
         \u_decoder/fir_filter/n1297 , \u_decoder/fir_filter/n1296 ,
         \u_decoder/fir_filter/n1295 , \u_decoder/fir_filter/n1294 ,
         \u_decoder/fir_filter/n1293 , \u_decoder/fir_filter/n1292 ,
         \u_decoder/fir_filter/n1291 , \u_decoder/fir_filter/n1290 ,
         \u_decoder/fir_filter/n1289 , \u_decoder/fir_filter/n1288 ,
         \u_decoder/fir_filter/n1286 , \u_decoder/fir_filter/n1285 ,
         \u_decoder/fir_filter/n1284 , \u_decoder/fir_filter/n1283 ,
         \u_decoder/fir_filter/n1282 , \u_decoder/fir_filter/n1281 ,
         \u_decoder/fir_filter/n1280 , \u_decoder/fir_filter/n1279 ,
         \u_decoder/fir_filter/n1278 , \u_decoder/fir_filter/n1277 ,
         \u_decoder/fir_filter/n1276 , \u_decoder/fir_filter/n1275 ,
         \u_decoder/fir_filter/n1274 , \u_decoder/fir_filter/n1273 ,
         \u_decoder/fir_filter/n1272 , \u_decoder/fir_filter/n1270 ,
         \u_decoder/fir_filter/n1269 , \u_decoder/fir_filter/n1268 ,
         \u_decoder/fir_filter/n1267 , \u_decoder/fir_filter/n1266 ,
         \u_decoder/fir_filter/n1265 , \u_decoder/fir_filter/n1264 ,
         \u_decoder/fir_filter/n1263 , \u_decoder/fir_filter/n1262 ,
         \u_decoder/fir_filter/n1261 , \u_decoder/fir_filter/n1260 ,
         \u_decoder/fir_filter/n1259 , \u_decoder/fir_filter/n1258 ,
         \u_decoder/fir_filter/n1257 , \u_decoder/fir_filter/n1254 ,
         \u_decoder/fir_filter/n1253 , \u_decoder/fir_filter/n1252 ,
         \u_decoder/fir_filter/n1251 , \u_decoder/fir_filter/n1250 ,
         \u_decoder/fir_filter/n1249 , \u_decoder/fir_filter/n1248 ,
         \u_decoder/fir_filter/n1247 , \u_decoder/fir_filter/n1246 ,
         \u_decoder/fir_filter/n1245 , \u_decoder/fir_filter/n1244 ,
         \u_decoder/fir_filter/n1243 , \u_decoder/fir_filter/n1242 ,
         \u_decoder/fir_filter/n1241 , \u_decoder/fir_filter/n1240 ,
         \u_decoder/fir_filter/n1238 , \u_decoder/fir_filter/n1237 ,
         \u_decoder/fir_filter/n1236 , \u_decoder/fir_filter/n1235 ,
         \u_decoder/fir_filter/n1234 , \u_decoder/fir_filter/n1233 ,
         \u_decoder/fir_filter/n1232 , \u_decoder/fir_filter/n1231 ,
         \u_decoder/fir_filter/n1230 , \u_decoder/fir_filter/n1229 ,
         \u_decoder/fir_filter/n1228 , \u_decoder/fir_filter/n1227 ,
         \u_decoder/fir_filter/n1226 , \u_decoder/fir_filter/n1225 ,
         \u_decoder/fir_filter/n1224 , \u_decoder/fir_filter/n1222 ,
         \u_decoder/fir_filter/n1221 , \u_decoder/fir_filter/n1220 ,
         \u_decoder/fir_filter/n1219 , \u_decoder/fir_filter/n1218 ,
         \u_decoder/fir_filter/n1217 , \u_decoder/fir_filter/n1216 ,
         \u_decoder/fir_filter/n1215 , \u_decoder/fir_filter/n1214 ,
         \u_decoder/fir_filter/n1213 , \u_decoder/fir_filter/n1212 ,
         \u_decoder/fir_filter/n1211 , \u_decoder/fir_filter/n1210 ,
         \u_decoder/fir_filter/n1209 , \u_decoder/fir_filter/n1206 ,
         \u_decoder/fir_filter/n1205 , \u_decoder/fir_filter/n1204 ,
         \u_decoder/fir_filter/n1203 , \u_decoder/fir_filter/n1202 ,
         \u_decoder/fir_filter/n1201 , \u_decoder/fir_filter/n1200 ,
         \u_decoder/fir_filter/n1199 , \u_decoder/fir_filter/n1198 ,
         \u_decoder/fir_filter/n1197 , \u_decoder/fir_filter/n1196 ,
         \u_decoder/fir_filter/n1195 , \u_decoder/fir_filter/n1194 ,
         \u_decoder/fir_filter/n1193 , \u_decoder/fir_filter/n1192 ,
         \u_decoder/fir_filter/n1190 , \u_decoder/fir_filter/n1189 ,
         \u_decoder/fir_filter/n1188 , \u_decoder/fir_filter/n1187 ,
         \u_decoder/fir_filter/n1186 , \u_decoder/fir_filter/n1185 ,
         \u_decoder/fir_filter/n1184 , \u_decoder/fir_filter/n1183 ,
         \u_decoder/fir_filter/n1182 , \u_decoder/fir_filter/n1181 ,
         \u_decoder/fir_filter/n1180 , \u_decoder/fir_filter/n1179 ,
         \u_decoder/fir_filter/n1178 , \u_decoder/fir_filter/n1177 ,
         \u_decoder/fir_filter/n1176 , \u_decoder/fir_filter/n1169 ,
         \u_decoder/fir_filter/n1168 , \u_decoder/fir_filter/n1167 ,
         \u_decoder/fir_filter/n1166 , \u_decoder/fir_filter/n1165 ,
         \u_decoder/fir_filter/n1164 , \u_decoder/fir_filter/n1163 ,
         \u_decoder/fir_filter/n1162 , \u_decoder/fir_filter/n1161 ,
         \u_decoder/fir_filter/n1160 , \u_decoder/fir_filter/n1159 ,
         \u_decoder/fir_filter/n1158 , \u_decoder/fir_filter/n1157 ,
         \u_decoder/fir_filter/n1156 , \u_decoder/fir_filter/n1155 ,
         \u_decoder/fir_filter/n1154 , \u_decoder/fir_filter/n1153 ,
         \u_decoder/fir_filter/n1152 , \u_decoder/fir_filter/n1151 ,
         \u_decoder/fir_filter/n1150 , \u_decoder/fir_filter/n1149 ,
         \u_decoder/fir_filter/n1148 , \u_decoder/fir_filter/n1147 ,
         \u_decoder/fir_filter/n1146 , \u_decoder/fir_filter/n1145 ,
         \u_decoder/fir_filter/n1144 , \u_decoder/fir_filter/n1143 ,
         \u_decoder/fir_filter/n1142 , \u_decoder/fir_filter/n1141 ,
         \u_decoder/fir_filter/n1140 , \u_decoder/fir_filter/n1139 ,
         \u_decoder/fir_filter/n1138 , \u_decoder/fir_filter/n1137 ,
         \u_decoder/fir_filter/n1136 , \u_decoder/fir_filter/n1135 ,
         \u_decoder/fir_filter/n1134 , \u_decoder/fir_filter/n1132 ,
         \u_decoder/fir_filter/n1131 , \u_decoder/fir_filter/n1130 ,
         \u_decoder/fir_filter/n1129 , \u_decoder/fir_filter/n1128 ,
         \u_decoder/fir_filter/n1127 , \u_decoder/fir_filter/n1126 ,
         \u_decoder/fir_filter/n1125 , \u_decoder/fir_filter/n1124 ,
         \u_decoder/fir_filter/n1123 , \u_decoder/fir_filter/n1122 ,
         \u_decoder/fir_filter/n1121 , \u_decoder/fir_filter/n1120 ,
         \u_decoder/fir_filter/n1119 , \u_decoder/fir_filter/n1118 ,
         \u_decoder/fir_filter/n1116 , \u_decoder/fir_filter/n1115 ,
         \u_decoder/fir_filter/n1114 , \u_decoder/fir_filter/n1113 ,
         \u_decoder/fir_filter/n1112 , \u_decoder/fir_filter/n1111 ,
         \u_decoder/fir_filter/n1110 , \u_decoder/fir_filter/n1109 ,
         \u_decoder/fir_filter/n1108 , \u_decoder/fir_filter/n1107 ,
         \u_decoder/fir_filter/n1106 , \u_decoder/fir_filter/n1105 ,
         \u_decoder/fir_filter/n1104 , \u_decoder/fir_filter/n1103 ,
         \u_decoder/fir_filter/n1102 , \u_decoder/fir_filter/n1100 ,
         \u_decoder/fir_filter/n1099 , \u_decoder/fir_filter/n1098 ,
         \u_decoder/fir_filter/n1097 , \u_decoder/fir_filter/n1096 ,
         \u_decoder/fir_filter/n1095 , \u_decoder/fir_filter/n1094 ,
         \u_decoder/fir_filter/n1093 , \u_decoder/fir_filter/n1092 ,
         \u_decoder/fir_filter/n1091 , \u_decoder/fir_filter/n1090 ,
         \u_decoder/fir_filter/n1089 , \u_decoder/fir_filter/n1088 ,
         \u_decoder/fir_filter/n1087 , \u_decoder/fir_filter/n1086 ,
         \u_decoder/fir_filter/n1084 , \u_decoder/fir_filter/n1083 ,
         \u_decoder/fir_filter/n1082 , \u_decoder/fir_filter/n1081 ,
         \u_decoder/fir_filter/n1080 , \u_decoder/fir_filter/n1079 ,
         \u_decoder/fir_filter/n1078 , \u_decoder/fir_filter/n1077 ,
         \u_decoder/fir_filter/n1076 , \u_decoder/fir_filter/n1075 ,
         \u_decoder/fir_filter/n1074 , \u_decoder/fir_filter/n1073 ,
         \u_decoder/fir_filter/n1072 , \u_decoder/fir_filter/n1071 ,
         \u_decoder/fir_filter/n1070 , \u_decoder/fir_filter/n1068 ,
         \u_decoder/fir_filter/n1067 , \u_decoder/fir_filter/n1066 ,
         \u_decoder/fir_filter/n1065 , \u_decoder/fir_filter/n1064 ,
         \u_decoder/fir_filter/n1063 , \u_decoder/fir_filter/n1062 ,
         \u_decoder/fir_filter/n1061 , \u_decoder/fir_filter/n1060 ,
         \u_decoder/fir_filter/n1059 , \u_decoder/fir_filter/n1058 ,
         \u_decoder/fir_filter/n1057 , \u_decoder/fir_filter/n1056 ,
         \u_decoder/fir_filter/n1055 , \u_decoder/fir_filter/n1054 ,
         \u_decoder/fir_filter/n1052 , \u_decoder/fir_filter/n1051 ,
         \u_decoder/fir_filter/n1050 , \u_decoder/fir_filter/n1049 ,
         \u_decoder/fir_filter/n1048 , \u_decoder/fir_filter/n1047 ,
         \u_decoder/fir_filter/n1046 , \u_decoder/fir_filter/n1045 ,
         \u_decoder/fir_filter/n1044 , \u_decoder/fir_filter/n1043 ,
         \u_decoder/fir_filter/n1042 , \u_decoder/fir_filter/n1041 ,
         \u_decoder/fir_filter/n1040 , \u_decoder/fir_filter/n1039 ,
         \u_decoder/fir_filter/n1038 , \u_decoder/fir_filter/n1037 ,
         \u_decoder/fir_filter/n1035 , \u_decoder/fir_filter/n1034 ,
         \u_decoder/fir_filter/n1033 , \u_decoder/fir_filter/n1032 ,
         \u_decoder/fir_filter/n1031 , \u_decoder/fir_filter/n1030 ,
         \u_decoder/fir_filter/n1029 , \u_decoder/fir_filter/n1028 ,
         \u_decoder/fir_filter/n1027 , \u_decoder/fir_filter/n1026 ,
         \u_decoder/fir_filter/n1025 , \u_decoder/fir_filter/n1024 ,
         \u_decoder/fir_filter/n1023 , \u_decoder/fir_filter/n1022 ,
         \u_decoder/fir_filter/n1021 , \u_decoder/fir_filter/n1020 ,
         \u_decoder/fir_filter/n1019 , \u_decoder/fir_filter/n1011 ,
         \u_decoder/fir_filter/n1010 , \u_decoder/fir_filter/n1009 ,
         \u_decoder/fir_filter/n1008 , \u_decoder/fir_filter/n1007 ,
         \u_decoder/fir_filter/n1006 , \u_decoder/fir_filter/n1005 ,
         \u_decoder/fir_filter/n1004 , \u_decoder/fir_filter/n1003 ,
         \u_decoder/fir_filter/n1002 , \u_decoder/fir_filter/n1001 ,
         \u_decoder/fir_filter/n1000 , \u_decoder/fir_filter/n999 ,
         \u_decoder/fir_filter/n998 , \u_decoder/fir_filter/n997 ,
         \u_decoder/fir_filter/n996 , \u_decoder/fir_filter/n995 ,
         \u_decoder/fir_filter/n994 , \u_decoder/fir_filter/n993 ,
         \u_decoder/fir_filter/n992 , \u_decoder/fir_filter/n991 ,
         \u_decoder/fir_filter/n990 , \u_decoder/fir_filter/n989 ,
         \u_decoder/fir_filter/n988 , \u_decoder/fir_filter/n987 ,
         \u_decoder/fir_filter/n986 , \u_decoder/fir_filter/n985 ,
         \u_decoder/fir_filter/n984 , \u_decoder/fir_filter/n983 ,
         \u_decoder/fir_filter/n982 , \u_decoder/fir_filter/n975 ,
         \u_decoder/fir_filter/n974 , \u_decoder/fir_filter/n973 ,
         \u_decoder/fir_filter/n972 , \u_decoder/fir_filter/n971 ,
         \u_decoder/fir_filter/n970 , \u_decoder/fir_filter/n969 ,
         \u_decoder/fir_filter/n968 , \u_decoder/fir_filter/n967 ,
         \u_decoder/fir_filter/n966 , \u_decoder/fir_filter/n965 ,
         \u_decoder/fir_filter/n964 , \u_decoder/fir_filter/n963 ,
         \u_decoder/fir_filter/n962 , \u_decoder/fir_filter/n961 ,
         \u_decoder/fir_filter/n954 , \u_decoder/fir_filter/n953 ,
         \u_decoder/fir_filter/n952 , \u_decoder/fir_filter/n951 ,
         \u_decoder/fir_filter/n950 , \u_decoder/fir_filter/n949 ,
         \u_decoder/fir_filter/n948 , \u_decoder/fir_filter/n947 ,
         \u_decoder/fir_filter/n946 , \u_decoder/fir_filter/n945 ,
         \u_decoder/fir_filter/n944 , \u_decoder/fir_filter/n943 ,
         \u_decoder/fir_filter/n942 , \u_decoder/fir_filter/n941 ,
         \u_decoder/fir_filter/n940 , \u_decoder/fir_filter/n933 ,
         \u_decoder/fir_filter/n932 , \u_decoder/fir_filter/n931 ,
         \u_decoder/fir_filter/n930 , \u_decoder/fir_filter/n929 ,
         \u_decoder/fir_filter/n928 , \u_decoder/fir_filter/n927 ,
         \u_decoder/fir_filter/n926 , \u_decoder/fir_filter/n925 ,
         \u_decoder/fir_filter/n924 , \u_decoder/fir_filter/n923 ,
         \u_decoder/fir_filter/n922 , \u_decoder/fir_filter/n921 ,
         \u_decoder/fir_filter/n920 , \u_decoder/fir_filter/n919 ,
         \u_decoder/fir_filter/n912 , \u_decoder/fir_filter/n911 ,
         \u_decoder/fir_filter/n910 , \u_decoder/fir_filter/n909 ,
         \u_decoder/fir_filter/n908 , \u_decoder/fir_filter/n907 ,
         \u_decoder/fir_filter/n906 , \u_decoder/fir_filter/n905 ,
         \u_decoder/fir_filter/n904 , \u_decoder/fir_filter/n903 ,
         \u_decoder/fir_filter/n902 , \u_decoder/fir_filter/n901 ,
         \u_decoder/fir_filter/n900 , \u_decoder/fir_filter/n899 ,
         \u_decoder/fir_filter/n898 , \u_decoder/fir_filter/n891 ,
         \u_decoder/fir_filter/n890 , \u_decoder/fir_filter/n889 ,
         \u_decoder/fir_filter/n888 , \u_decoder/fir_filter/n887 ,
         \u_decoder/fir_filter/n886 , \u_decoder/fir_filter/n885 ,
         \u_decoder/fir_filter/n884 , \u_decoder/fir_filter/n883 ,
         \u_decoder/fir_filter/n882 , \u_decoder/fir_filter/n881 ,
         \u_decoder/fir_filter/n880 , \u_decoder/fir_filter/n879 ,
         \u_decoder/fir_filter/n878 , \u_decoder/fir_filter/n877 ,
         \u_decoder/fir_filter/n870 , \u_decoder/fir_filter/n869 ,
         \u_decoder/fir_filter/n868 , \u_decoder/fir_filter/n867 ,
         \u_decoder/fir_filter/n866 , \u_decoder/fir_filter/n865 ,
         \u_decoder/fir_filter/n864 , \u_decoder/fir_filter/n863 ,
         \u_decoder/fir_filter/n862 , \u_decoder/fir_filter/n861 ,
         \u_decoder/fir_filter/n860 , \u_decoder/fir_filter/n859 ,
         \u_decoder/fir_filter/n858 , \u_decoder/fir_filter/n857 ,
         \u_decoder/fir_filter/n856 , \u_decoder/fir_filter/n855 ,
         \u_decoder/fir_filter/n854 , \u_decoder/fir_filter/n853 ,
         \u_decoder/fir_filter/n852 , \u_decoder/fir_filter/n851 ,
         \u_decoder/fir_filter/n850 , \u_decoder/fir_filter/n849 ,
         \u_decoder/fir_filter/n848 , \u_decoder/fir_filter/n847 ,
         \u_decoder/fir_filter/n846 , \u_decoder/fir_filter/n845 ,
         \u_decoder/fir_filter/n844 , \u_decoder/fir_filter/n843 ,
         \u_decoder/fir_filter/n842 , \u_decoder/fir_filter/n841 ,
         \u_decoder/fir_filter/n840 , \u_decoder/fir_filter/n839 ,
         \u_decoder/fir_filter/n838 , \u_decoder/fir_filter/n837 ,
         \u_decoder/fir_filter/n835 , \u_decoder/fir_filter/n834 ,
         \u_decoder/fir_filter/n833 , \u_decoder/fir_filter/n832 ,
         \u_decoder/fir_filter/n831 , \u_decoder/fir_filter/n830 ,
         \u_decoder/fir_filter/n829 , \u_decoder/fir_filter/n828 ,
         \u_decoder/fir_filter/n827 , \u_decoder/fir_filter/n826 ,
         \u_decoder/fir_filter/n825 , \u_decoder/fir_filter/n824 ,
         \u_decoder/fir_filter/n823 , \u_decoder/fir_filter/n822 ,
         \u_decoder/fir_filter/n821 , \u_decoder/fir_filter/n819 ,
         \u_decoder/fir_filter/n818 , \u_decoder/fir_filter/n817 ,
         \u_decoder/fir_filter/n816 , \u_decoder/fir_filter/n815 ,
         \u_decoder/fir_filter/n814 , \u_decoder/fir_filter/n813 ,
         \u_decoder/fir_filter/n812 , \u_decoder/fir_filter/n811 ,
         \u_decoder/fir_filter/n810 , \u_decoder/fir_filter/n809 ,
         \u_decoder/fir_filter/n808 , \u_decoder/fir_filter/n807 ,
         \u_decoder/fir_filter/n806 , \u_decoder/fir_filter/n805 ,
         \u_decoder/fir_filter/n803 , \u_decoder/fir_filter/n802 ,
         \u_decoder/fir_filter/n801 , \u_decoder/fir_filter/n800 ,
         \u_decoder/fir_filter/n799 , \u_decoder/fir_filter/n798 ,
         \u_decoder/fir_filter/n797 , \u_decoder/fir_filter/n796 ,
         \u_decoder/fir_filter/n795 , \u_decoder/fir_filter/n794 ,
         \u_decoder/fir_filter/n793 , \u_decoder/fir_filter/n792 ,
         \u_decoder/fir_filter/n791 , \u_decoder/fir_filter/n790 ,
         \u_decoder/fir_filter/n789 , \u_decoder/fir_filter/n787 ,
         \u_decoder/fir_filter/n786 , \u_decoder/fir_filter/n785 ,
         \u_decoder/fir_filter/n784 , \u_decoder/fir_filter/n783 ,
         \u_decoder/fir_filter/n782 , \u_decoder/fir_filter/n781 ,
         \u_decoder/fir_filter/n780 , \u_decoder/fir_filter/n779 ,
         \u_decoder/fir_filter/n778 , \u_decoder/fir_filter/n777 ,
         \u_decoder/fir_filter/n776 , \u_decoder/fir_filter/n775 ,
         \u_decoder/fir_filter/n774 , \u_decoder/fir_filter/n773 ,
         \u_decoder/fir_filter/n771 , \u_decoder/fir_filter/n770 ,
         \u_decoder/fir_filter/n769 , \u_decoder/fir_filter/n768 ,
         \u_decoder/fir_filter/n767 , \u_decoder/fir_filter/n766 ,
         \u_decoder/fir_filter/n765 , \u_decoder/fir_filter/n764 ,
         \u_decoder/fir_filter/n763 , \u_decoder/fir_filter/n762 ,
         \u_decoder/fir_filter/n761 , \u_decoder/fir_filter/n760 ,
         \u_decoder/fir_filter/n759 , \u_decoder/fir_filter/n758 ,
         \u_decoder/fir_filter/n757 , \u_decoder/fir_filter/n755 ,
         \u_decoder/fir_filter/n754 , \u_decoder/fir_filter/n753 ,
         \u_decoder/fir_filter/n752 , \u_decoder/fir_filter/n751 ,
         \u_decoder/fir_filter/n750 , \u_decoder/fir_filter/n749 ,
         \u_decoder/fir_filter/n748 , \u_decoder/fir_filter/n747 ,
         \u_decoder/fir_filter/n746 , \u_decoder/fir_filter/n745 ,
         \u_decoder/fir_filter/n744 , \u_decoder/fir_filter/n743 ,
         \u_decoder/fir_filter/n742 , \u_decoder/fir_filter/n741 ,
         \u_decoder/fir_filter/n740 , \u_decoder/fir_filter/n738 ,
         \u_decoder/fir_filter/n737 , \u_decoder/fir_filter/n736 ,
         \u_decoder/fir_filter/n735 , \u_decoder/fir_filter/n734 ,
         \u_decoder/fir_filter/n733 , \u_decoder/fir_filter/n732 ,
         \u_decoder/fir_filter/n731 , \u_decoder/fir_filter/n730 ,
         \u_decoder/fir_filter/n729 , \u_decoder/fir_filter/n728 ,
         \u_decoder/fir_filter/n727 , \u_decoder/fir_filter/n726 ,
         \u_decoder/fir_filter/n725 , \u_decoder/fir_filter/n724 ,
         \u_decoder/fir_filter/n723 , \u_decoder/fir_filter/n722 ,
         \u_decoder/fir_filter/n721 , \u_decoder/fir_filter/n713 ,
         \u_decoder/fir_filter/n712 , \u_decoder/fir_filter/n711 ,
         \u_decoder/fir_filter/n710 , \u_decoder/fir_filter/n709 ,
         \u_decoder/fir_filter/n708 , \u_decoder/fir_filter/n707 ,
         \u_decoder/fir_filter/n706 , \u_decoder/fir_filter/n705 ,
         \u_decoder/fir_filter/n704 , \u_decoder/fir_filter/n703 ,
         \u_decoder/fir_filter/n702 , \u_decoder/fir_filter/n701 ,
         \u_decoder/fir_filter/n700 , \u_decoder/fir_filter/n699 ,
         \u_decoder/fir_filter/n698 , \u_decoder/fir_filter/n697 ,
         \u_decoder/fir_filter/n696 , \u_decoder/fir_filter/n695 ,
         \u_decoder/fir_filter/n694 , \u_decoder/fir_filter/n693 ,
         \u_decoder/fir_filter/n692 , \u_decoder/fir_filter/n691 ,
         \u_decoder/fir_filter/n690 , \u_decoder/fir_filter/n689 ,
         \u_decoder/fir_filter/n688 , \u_decoder/fir_filter/n687 ,
         \u_decoder/fir_filter/n686 , \u_decoder/fir_filter/n685 ,
         \u_decoder/fir_filter/n684 , \u_decoder/fir_filter/n677 ,
         \u_decoder/fir_filter/n676 , \u_decoder/fir_filter/n675 ,
         \u_decoder/fir_filter/n674 , \u_decoder/fir_filter/n673 ,
         \u_decoder/fir_filter/n672 , \u_decoder/fir_filter/n671 ,
         \u_decoder/fir_filter/n670 , \u_decoder/fir_filter/n669 ,
         \u_decoder/fir_filter/n668 , \u_decoder/fir_filter/n667 ,
         \u_decoder/fir_filter/n666 , \u_decoder/fir_filter/n665 ,
         \u_decoder/fir_filter/n664 , \u_decoder/fir_filter/n663 ,
         \u_decoder/fir_filter/n656 , \u_decoder/fir_filter/n655 ,
         \u_decoder/fir_filter/n654 , \u_decoder/fir_filter/n653 ,
         \u_decoder/fir_filter/n652 , \u_decoder/fir_filter/n651 ,
         \u_decoder/fir_filter/n650 , \u_decoder/fir_filter/n649 ,
         \u_decoder/fir_filter/n648 , \u_decoder/fir_filter/n647 ,
         \u_decoder/fir_filter/n646 , \u_decoder/fir_filter/n645 ,
         \u_decoder/fir_filter/n644 , \u_decoder/fir_filter/n643 ,
         \u_decoder/fir_filter/n642 , \u_decoder/fir_filter/n635 ,
         \u_decoder/fir_filter/n634 , \u_decoder/fir_filter/n633 ,
         \u_decoder/fir_filter/n632 , \u_decoder/fir_filter/n631 ,
         \u_decoder/fir_filter/n630 , \u_decoder/fir_filter/n629 ,
         \u_decoder/fir_filter/n628 , \u_decoder/fir_filter/n627 ,
         \u_decoder/fir_filter/n626 , \u_decoder/fir_filter/n625 ,
         \u_decoder/fir_filter/n624 , \u_decoder/fir_filter/n623 ,
         \u_decoder/fir_filter/n622 , \u_decoder/fir_filter/n621 ,
         \u_decoder/fir_filter/n614 , \u_decoder/fir_filter/n613 ,
         \u_decoder/fir_filter/n612 , \u_decoder/fir_filter/n611 ,
         \u_decoder/fir_filter/n610 , \u_decoder/fir_filter/n609 ,
         \u_decoder/fir_filter/n608 , \u_decoder/fir_filter/n607 ,
         \u_decoder/fir_filter/n606 , \u_decoder/fir_filter/n605 ,
         \u_decoder/fir_filter/n604 , \u_decoder/fir_filter/n603 ,
         \u_decoder/fir_filter/n602 , \u_decoder/fir_filter/n601 ,
         \u_decoder/fir_filter/n600 , \u_decoder/fir_filter/n593 ,
         \u_decoder/fir_filter/n592 , \u_decoder/fir_filter/n591 ,
         \u_decoder/fir_filter/n590 , \u_decoder/fir_filter/n589 ,
         \u_decoder/fir_filter/n588 , \u_decoder/fir_filter/n587 ,
         \u_decoder/fir_filter/n586 , \u_decoder/fir_filter/n585 ,
         \u_decoder/fir_filter/n584 , \u_decoder/fir_filter/n583 ,
         \u_decoder/fir_filter/n582 , \u_decoder/fir_filter/n581 ,
         \u_decoder/fir_filter/n580 , \u_decoder/fir_filter/n579 ,
         \u_decoder/fir_filter/n572 , \u_decoder/fir_filter/n571 ,
         \u_decoder/fir_filter/n570 , \u_decoder/fir_filter/n569 ,
         \u_decoder/fir_filter/n568 , \u_decoder/fir_filter/n567 ,
         \u_decoder/fir_filter/n566 , \u_decoder/fir_filter/n565 ,
         \u_decoder/fir_filter/n564 , \u_decoder/fir_filter/n563 ,
         \u_decoder/fir_filter/n562 , \u_decoder/fir_filter/n561 ,
         \u_decoder/fir_filter/n560 , \u_decoder/fir_filter/n559 ,
         \u_decoder/fir_filter/n558 , \u_decoder/fir_filter/n557 ,
         \u_decoder/fir_filter/n556 , \u_decoder/fir_filter/n555 ,
         \u_decoder/fir_filter/n554 , \u_decoder/fir_filter/n553 ,
         \u_decoder/fir_filter/n442 , \u_decoder/fir_filter/n441 ,
         \u_decoder/fir_filter/n440 , \u_decoder/fir_filter/n439 ,
         \u_decoder/fir_filter/n438 , \u_decoder/fir_filter/n437 ,
         \u_decoder/fir_filter/n436 , \u_decoder/fir_filter/n435 ,
         \u_decoder/fir_filter/n434 , \u_decoder/fir_filter/n433 ,
         \u_decoder/fir_filter/n432 , \u_decoder/fir_filter/n431 ,
         \u_decoder/fir_filter/n430 , \u_decoder/fir_filter/n429 ,
         \u_decoder/fir_filter/n428 , \u_decoder/fir_filter/n426 ,
         \u_decoder/fir_filter/n425 , \u_decoder/fir_filter/n424 ,
         \u_decoder/fir_filter/n423 , \u_decoder/fir_filter/n422 ,
         \u_decoder/fir_filter/n421 , \u_decoder/fir_filter/n420 ,
         \u_decoder/fir_filter/n419 , \u_decoder/fir_filter/n418 ,
         \u_decoder/fir_filter/n417 , \u_decoder/fir_filter/n416 ,
         \u_decoder/fir_filter/n415 , \u_decoder/fir_filter/n414 ,
         \u_decoder/fir_filter/n413 , \u_decoder/fir_filter/n412 ,
         \u_decoder/fir_filter/n410 , \u_decoder/fir_filter/Q_data_mult_2[8] ,
         \u_decoder/fir_filter/Q_data_mult_2_15 ,
         \u_decoder/fir_filter/Q_data_mult_1[4] ,
         \u_decoder/fir_filter/Q_data_mult_1_15 ,
         \u_decoder/fir_filter/Q_data_mult_0_15 ,
         \u_decoder/fir_filter/I_data_mult_2[8] ,
         \u_decoder/fir_filter/I_data_mult_2_15 ,
         \u_decoder/fir_filter/I_data_mult_1[4] ,
         \u_decoder/fir_filter/I_data_mult_1_15 ,
         \u_decoder/fir_filter/I_data_mult_0_15 , \u_decoder/fir_filter/N12 ,
         \u_decoder/fir_filter/N11 , \u_cordic/mycordic/n587 ,
         \u_cordic/mycordic/n586 , \u_cordic/mycordic/n585 ,
         \u_cordic/mycordic/n584 , \u_cordic/mycordic/n583 ,
         \u_cordic/mycordic/n582 , \u_cordic/mycordic/n581 ,
         \u_cordic/mycordic/n580 , \u_cordic/mycordic/n579 ,
         \u_cordic/mycordic/n578 , \u_cordic/mycordic/n577 ,
         \u_cordic/mycordic/n576 , \u_cordic/mycordic/n575 ,
         \u_cordic/mycordic/n574 , \u_cordic/mycordic/n573 ,
         \u_cordic/mycordic/n572 , \u_cordic/mycordic/n571 ,
         \u_cordic/mycordic/n570 , \u_cordic/mycordic/n569 ,
         \u_cordic/mycordic/n568 , \u_cordic/mycordic/n567 ,
         \u_cordic/mycordic/n566 , \u_cordic/mycordic/n565 ,
         \u_cordic/mycordic/n564 , \u_cordic/mycordic/n563 ,
         \u_cordic/mycordic/n562 , \u_cordic/mycordic/n561 ,
         \u_cordic/mycordic/n560 , \u_cordic/mycordic/n559 ,
         \u_cordic/mycordic/n558 , \u_cordic/mycordic/n557 ,
         \u_cordic/mycordic/n556 , \u_cordic/mycordic/n555 ,
         \u_cordic/mycordic/n554 , \u_cordic/mycordic/n553 ,
         \u_cordic/mycordic/n552 , \u_cordic/mycordic/n551 ,
         \u_cordic/mycordic/n550 , \u_cordic/mycordic/n549 ,
         \u_cordic/mycordic/n548 , \u_cordic/mycordic/n547 ,
         \u_cordic/mycordic/n546 , \u_cordic/mycordic/n545 ,
         \u_cordic/mycordic/n544 , \u_cordic/mycordic/n543 ,
         \u_cordic/mycordic/n542 , \u_cordic/mycordic/n541 ,
         \u_cordic/mycordic/n540 , \u_cordic/mycordic/n539 ,
         \u_cordic/mycordic/n538 , \u_cordic/mycordic/n537 ,
         \u_cordic/mycordic/n536 , \u_cordic/mycordic/n520 ,
         \u_cordic/mycordic/n519 , \u_cordic/mycordic/n518 ,
         \u_cordic/mycordic/n517 , \u_cordic/mycordic/n516 ,
         \u_cordic/mycordic/n515 , \u_cordic/mycordic/n514 ,
         \u_cordic/mycordic/n513 , \u_cordic/mycordic/n512 ,
         \u_cordic/mycordic/n511 , \u_cordic/mycordic/n510 ,
         \u_cordic/mycordic/n509 , \u_cordic/mycordic/n508 ,
         \u_cordic/mycordic/n507 , \u_cordic/mycordic/n506 ,
         \u_cordic/mycordic/n505 , \u_cordic/mycordic/n504 ,
         \u_cordic/mycordic/n503 , \u_cordic/mycordic/n502 ,
         \u_cordic/mycordic/n501 , \u_cordic/mycordic/n500 ,
         \u_cordic/mycordic/n499 , \u_cordic/mycordic/n498 ,
         \u_cordic/mycordic/n497 , \u_cordic/mycordic/n496 ,
         \u_cordic/mycordic/n495 , \u_cordic/mycordic/n494 ,
         \u_cordic/mycordic/n493 , \u_cordic/mycordic/n492 ,
         \u_cordic/mycordic/n491 , \u_cordic/mycordic/n490 ,
         \u_cordic/mycordic/n489 , \u_cordic/mycordic/n488 ,
         \u_cordic/mycordic/n487 , \u_cordic/mycordic/n486 ,
         \u_cordic/mycordic/n485 , \u_cordic/mycordic/n484 ,
         \u_cordic/mycordic/n483 , \u_cordic/mycordic/n482 ,
         \u_cordic/mycordic/n481 , \u_cordic/mycordic/n480 ,
         \u_cordic/mycordic/n479 , \u_cordic/mycordic/n478 ,
         \u_cordic/mycordic/n477 , \u_cordic/mycordic/n476 ,
         \u_cordic/mycordic/n475 , \u_cordic/mycordic/n474 ,
         \u_cordic/mycordic/n473 , \u_cordic/mycordic/n472 ,
         \u_cordic/mycordic/n471 , \u_cordic/mycordic/n470 ,
         \u_cordic/mycordic/n469 , \u_cordic/mycordic/n468 ,
         \u_cordic/mycordic/n467 , \u_cordic/mycordic/n466 ,
         \u_cordic/mycordic/n465 , \u_cordic/mycordic/n464 ,
         \u_cordic/mycordic/n463 , \u_cordic/mycordic/n462 ,
         \u_cordic/mycordic/n461 , \u_cordic/mycordic/n460 ,
         \u_cordic/mycordic/n459 , \u_cordic/mycordic/n458 ,
         \u_cordic/mycordic/n457 , \u_cordic/mycordic/n456 ,
         \u_cordic/mycordic/n455 , \u_cordic/mycordic/n454 ,
         \u_cordic/mycordic/n453 , \u_cordic/mycordic/n452 ,
         \u_cordic/mycordic/n451 , \u_cordic/mycordic/n450 ,
         \u_cordic/mycordic/n449 , \u_cordic/mycordic/n448 ,
         \u_cordic/mycordic/n447 , \u_cordic/mycordic/n446 ,
         \u_cordic/mycordic/n445 , \u_cordic/mycordic/n444 ,
         \u_cordic/mycordic/n443 , \u_cordic/mycordic/n442 ,
         \u_cordic/mycordic/n441 , \u_cordic/mycordic/n440 ,
         \u_cordic/mycordic/n439 , \u_cordic/mycordic/n438 ,
         \u_cordic/mycordic/n437 , \u_cordic/mycordic/n436 ,
         \u_cordic/mycordic/n435 , \u_cordic/mycordic/n433 ,
         \u_cordic/mycordic/n432 , \u_cordic/mycordic/n431 ,
         \u_cordic/mycordic/n430 , \u_cordic/mycordic/n429 ,
         \u_cordic/mycordic/n428 , \u_cordic/mycordic/n427 ,
         \u_cordic/mycordic/n426 , \u_cordic/mycordic/n425 ,
         \u_cordic/mycordic/n424 , \u_cordic/mycordic/n423 ,
         \u_cordic/mycordic/n422 , \u_cordic/mycordic/n421 ,
         \u_cordic/mycordic/n420 , \u_cordic/mycordic/n419 ,
         \u_cordic/mycordic/n418 , \u_cordic/mycordic/n417 ,
         \u_cordic/mycordic/n416 , \u_cordic/mycordic/n415 ,
         \u_cordic/mycordic/n414 , \u_cordic/mycordic/n413 ,
         \u_cordic/mycordic/n412 , \u_cordic/mycordic/n411 ,
         \u_cordic/mycordic/n410 , \u_cordic/mycordic/n409 ,
         \u_cordic/mycordic/n408 , \u_cordic/mycordic/n407 ,
         \u_cordic/mycordic/n406 , \u_cordic/mycordic/n405 ,
         \u_cordic/mycordic/n404 , \u_cordic/mycordic/n403 ,
         \u_cordic/mycordic/n402 , \u_cordic/mycordic/n401 ,
         \u_cordic/mycordic/n400 , \u_cordic/mycordic/n399 ,
         \u_cordic/mycordic/n395 , \u_cordic/mycordic/n394 ,
         \u_cordic/mycordic/n393 , \u_cordic/mycordic/n392 ,
         \u_cordic/mycordic/n391 , \u_cordic/mycordic/n387 ,
         \u_cordic/mycordic/n386 , \u_cordic/mycordic/n385 ,
         \u_cordic/mycordic/n384 , \u_cordic/mycordic/n383 ,
         \u_cordic/mycordic/n382 , \u_cordic/mycordic/n381 ,
         \u_cordic/mycordic/n380 , \u_cordic/mycordic/n379 ,
         \u_cordic/mycordic/n378 , \u_cordic/mycordic/n377 ,
         \u_cordic/mycordic/n376 , \u_cordic/mycordic/n375 ,
         \u_cordic/mycordic/n374 , \u_cordic/mycordic/n373 ,
         \u_cordic/mycordic/n372 , \u_cordic/mycordic/n371 ,
         \u_cordic/mycordic/n370 , \u_cordic/mycordic/n369 ,
         \u_cordic/mycordic/n368 , \u_cordic/mycordic/n367 ,
         \u_cordic/mycordic/n366 , \u_cordic/mycordic/n365 ,
         \u_cordic/mycordic/n364 , \u_cordic/mycordic/n363 ,
         \u_cordic/mycordic/n362 , \u_cordic/mycordic/n358 ,
         \u_cordic/mycordic/n357 , \u_cordic/mycordic/n356 ,
         \u_cordic/mycordic/n355 , \u_cordic/mycordic/n354 ,
         \u_cordic/mycordic/n353 , \u_cordic/mycordic/n349 ,
         \u_cordic/mycordic/n348 , \u_cordic/mycordic/n347 ,
         \u_cordic/mycordic/n346 , \u_cordic/mycordic/n345 ,
         \u_cordic/mycordic/n344 , \u_cordic/mycordic/n343 ,
         \u_cordic/mycordic/n342 , \u_cordic/mycordic/n341 ,
         \u_cordic/mycordic/n340 , \u_cordic/mycordic/n339 ,
         \u_cordic/mycordic/n338 , \u_cordic/mycordic/n337 ,
         \u_cordic/mycordic/n336 , \u_cordic/mycordic/n335 ,
         \u_cordic/mycordic/n334 , \u_cordic/mycordic/n333 ,
         \u_cordic/mycordic/n332 , \u_cordic/mycordic/n331 ,
         \u_cordic/mycordic/n110 , \u_cordic/mycordic/n108 ,
         \u_cordic/mycordic/N630 , \u_cordic/mycordic/N629 ,
         \u_cordic/mycordic/N628 , \u_cordic/mycordic/N627 ,
         \u_cordic/mycordic/N626 , \u_cordic/mycordic/N625 ,
         \u_cordic/mycordic/N624 , \u_cordic/mycordic/N623 ,
         \u_cordic/mycordic/N622 , \u_cordic/mycordic/N621 ,
         \u_cordic/mycordic/N620 , \u_cordic/mycordic/N619 ,
         \u_cordic/mycordic/N615 , \u_cordic/mycordic/N565 ,
         \u_cordic/mycordic/N564 , \u_cordic/mycordic/N563 ,
         \u_cordic/mycordic/N562 , \u_cordic/mycordic/N561 ,
         \u_cordic/mycordic/N560 , \u_cordic/mycordic/N559 ,
         \u_cordic/mycordic/N558 , \u_cordic/mycordic/N557 ,
         \u_cordic/mycordic/N556 , \u_cordic/mycordic/N555 ,
         \u_cordic/mycordic/N554 , \u_cordic/mycordic/N553 ,
         \u_cordic/mycordic/N552 , \u_cordic/mycordic/N550 ,
         \u_cordic/mycordic/N549 , \u_cordic/mycordic/N548 ,
         \u_cordic/mycordic/N547 , \u_cordic/mycordic/N546 ,
         \u_cordic/mycordic/N545 , \u_cordic/mycordic/N544 ,
         \u_cordic/mycordic/N543 , \u_cordic/mycordic/N542 ,
         \u_cordic/mycordic/N541 , \u_cordic/mycordic/N540 ,
         \u_cordic/mycordic/N539 , \u_cordic/mycordic/N538 ,
         \u_cordic/mycordic/N537 , \u_cordic/mycordic/N536 ,
         \u_cordic/mycordic/N533 , \u_cordic/mycordic/N532 ,
         \u_cordic/mycordic/N531 , \u_cordic/mycordic/N530 ,
         \u_cordic/mycordic/N529 , \u_cordic/mycordic/N528 ,
         \u_cordic/mycordic/N527 , \u_cordic/mycordic/N526 ,
         \u_cordic/mycordic/N525 , \u_cordic/mycordic/N524 ,
         \u_cordic/mycordic/N523 , \u_cordic/mycordic/N522 ,
         \u_cordic/mycordic/N521 , \u_cordic/mycordic/N520 ,
         \u_cordic/mycordic/N519 , \u_cordic/mycordic/N517 ,
         \u_cordic/mycordic/N516 , \u_cordic/mycordic/N515 ,
         \u_cordic/mycordic/N514 , \u_cordic/mycordic/N513 ,
         \u_cordic/mycordic/N512 , \u_cordic/mycordic/N511 ,
         \u_cordic/mycordic/N510 , \u_cordic/mycordic/N509 ,
         \u_cordic/mycordic/N508 , \u_cordic/mycordic/N507 ,
         \u_cordic/mycordic/N506 , \u_cordic/mycordic/N505 ,
         \u_cordic/mycordic/N504 , \u_cordic/mycordic/N503 ,
         \u_cordic/mycordic/N502 , \u_cordic/mycordic/N500 ,
         \u_cordic/mycordic/N499 , \u_cordic/mycordic/N498 ,
         \u_cordic/mycordic/N497 , \u_cordic/mycordic/N496 ,
         \u_cordic/mycordic/N495 , \u_cordic/mycordic/N494 ,
         \u_cordic/mycordic/N493 , \u_cordic/mycordic/N492 ,
         \u_cordic/mycordic/N491 , \u_cordic/mycordic/N490 ,
         \u_cordic/mycordic/N489 , \u_cordic/mycordic/N488 ,
         \u_cordic/mycordic/N487 , \u_cordic/mycordic/N486 ,
         \u_cordic/mycordic/N485 , \u_cordic/mycordic/N483 ,
         \u_cordic/mycordic/N482 , \u_cordic/mycordic/N481 ,
         \u_cordic/mycordic/N480 , \u_cordic/mycordic/N479 ,
         \u_cordic/mycordic/N478 , \u_cordic/mycordic/N477 ,
         \u_cordic/mycordic/N476 , \u_cordic/mycordic/N475 ,
         \u_cordic/mycordic/N474 , \u_cordic/mycordic/N473 ,
         \u_cordic/mycordic/N472 , \u_cordic/mycordic/N471 ,
         \u_cordic/mycordic/N470 , \u_cordic/mycordic/N469 ,
         \u_cordic/mycordic/N468 , \u_cordic/mycordic/N467 ,
         \u_cordic/mycordic/N466 , \u_cordic/mycordic/N465 ,
         \u_cordic/mycordic/N464 , \u_cordic/mycordic/N463 ,
         \u_cordic/mycordic/N462 , \u_cordic/mycordic/N461 ,
         \u_cordic/mycordic/N460 , \u_cordic/mycordic/N459 ,
         \u_cordic/mycordic/N458 , \u_cordic/mycordic/N457 ,
         \u_cordic/mycordic/N455 , \u_cordic/mycordic/N454 ,
         \u_cordic/mycordic/N453 , \u_cordic/mycordic/N452 ,
         \u_cordic/mycordic/N451 , \u_cordic/mycordic/N450 ,
         \u_cordic/mycordic/N449 , \u_cordic/mycordic/N448 ,
         \u_cordic/mycordic/N447 , \u_cordic/mycordic/N446 ,
         \u_cordic/mycordic/N445 , \u_cordic/mycordic/N444 ,
         \u_cordic/mycordic/N443 , \u_cordic/mycordic/N442 ,
         \u_cordic/mycordic/N441 , \u_cordic/mycordic/N440 ,
         \u_cordic/mycordic/N439 , \u_cordic/mycordic/N438 ,
         \u_cordic/mycordic/N437 , \u_cordic/mycordic/N436 ,
         \u_cordic/mycordic/N435 , \u_cordic/mycordic/N434 ,
         \u_cordic/mycordic/N433 , \u_cordic/mycordic/N432 ,
         \u_cordic/mycordic/N431 , \u_cordic/mycordic/N430 ,
         \u_cordic/mycordic/N428 , \u_cordic/mycordic/N427 ,
         \u_cordic/mycordic/N426 , \u_cordic/mycordic/N425 ,
         \u_cordic/mycordic/N424 , \u_cordic/mycordic/N423 ,
         \u_cordic/mycordic/N422 , \u_cordic/mycordic/N421 ,
         \u_cordic/mycordic/N420 , \u_cordic/mycordic/N419 ,
         \u_cordic/mycordic/N418 , \u_cordic/mycordic/N417 ,
         \u_cordic/mycordic/N416 , \u_cordic/mycordic/N415 ,
         \u_cordic/mycordic/N414 , \u_cordic/mycordic/N413 ,
         \u_cordic/mycordic/N412 , \u_cordic/mycordic/N411 ,
         \u_cordic/mycordic/N410 , \u_cordic/mycordic/N409 ,
         \u_cordic/mycordic/N408 , \u_cordic/mycordic/N407 ,
         \u_cordic/mycordic/N406 , \u_cordic/mycordic/N405 ,
         \u_cordic/mycordic/N404 , \u_cordic/mycordic/N403 ,
         \u_cordic/mycordic/N402 , \u_cordic/mycordic/N401 ,
         \u_cordic/mycordic/N400 , \u_cordic/mycordic/N399 ,
         \u_cordic/mycordic/N398 , \u_cordic/mycordic/N395 ,
         \u_cordic/mycordic/N394 , \u_cordic/mycordic/N393 ,
         \u_cordic/mycordic/N392 , \u_cordic/mycordic/N391 ,
         \u_cordic/mycordic/N390 , \u_cordic/mycordic/N389 ,
         \u_cordic/mycordic/N388 , \u_cordic/mycordic/N387 ,
         \u_cordic/mycordic/N386 , \u_cordic/mycordic/N385 ,
         \u_cordic/mycordic/N384 , \u_cordic/mycordic/N383 ,
         \u_cordic/mycordic/N382 , \u_cordic/mycordic/N381 ,
         \u_cordic/mycordic/N380 , \u_cordic/mycordic/N379 ,
         \u_cordic/mycordic/N378 , \u_cordic/mycordic/N377 ,
         \u_cordic/mycordic/N376 , \u_cordic/mycordic/N375 ,
         \u_cordic/mycordic/N374 , \u_cordic/mycordic/N373 ,
         \u_cordic/mycordic/N372 , \u_cordic/mycordic/N371 ,
         \u_cordic/mycordic/N370 , \u_cordic/mycordic/N369 ,
         \u_cordic/mycordic/N368 , \u_cordic/mycordic/N367 ,
         \u_cordic/mycordic/N366 , \u_cordic/mycordic/N365 ,
         \u_cordic/mycordic/N363 , \u_cordic/mycordic/N362 ,
         \u_cordic/mycordic/N361 , \u_cordic/mycordic/N360 ,
         \u_cordic/mycordic/N359 , \u_cordic/mycordic/N358 ,
         \u_cordic/mycordic/N357 , \u_cordic/mycordic/N356 ,
         \u_cordic/mycordic/N355 , \u_cordic/mycordic/N354 ,
         \u_cordic/mycordic/N353 , \u_cordic/mycordic/N352 ,
         \u_cordic/mycordic/N351 , \u_cordic/mycordic/N350 ,
         \u_cordic/mycordic/N349 , \u_cordic/mycordic/N348 ,
         \u_cordic/mycordic/N347 , \u_cordic/mycordic/N346 ,
         \u_cordic/mycordic/N345 , \u_cordic/mycordic/N344 ,
         \u_cordic/mycordic/N343 , \u_cordic/mycordic/N342 ,
         \u_cordic/mycordic/N341 , \u_cordic/mycordic/N340 ,
         \u_cordic/mycordic/N339 , \u_cordic/mycordic/N338 ,
         \u_cordic/mycordic/N337 , \u_cordic/mycordic/N336 ,
         \u_cordic/mycordic/N335 , \u_cordic/mycordic/N334 ,
         \u_cordic/mycordic/N333 , \u_cordic/mycordic/N331 ,
         \u_cordic/mycordic/N330 , \u_cordic/mycordic/N329 ,
         \u_cordic/mycordic/N328 , \u_cordic/mycordic/N327 ,
         \u_cordic/mycordic/N326 , \u_cordic/mycordic/N325 ,
         \u_cordic/mycordic/N324 , \u_cordic/mycordic/N323 ,
         \u_cordic/mycordic/N322 , \u_cordic/mycordic/N321 ,
         \u_cordic/mycordic/N320 , \u_cordic/mycordic/N319 ,
         \u_cordic/mycordic/N318 , \u_cordic/mycordic/N317 ,
         \u_cordic/mycordic/N316 , \u_cordic/mycordic/N291 ,
         \u_cordic/mycordic/N290 , \u_cordic/mycordic/N289 ,
         \u_cordic/mycordic/N288 , \u_cordic/mycordic/N287 ,
         \u_cordic/mycordic/N267 , \u_cordic/mycordic/N266 ,
         \u_cordic/mycordic/N265 , \u_cordic/mycordic/N264 ,
         \u_cordic/mycordic/N263 , \u_cordic/mycordic/N259 ,
         \u_cordic/mycordic/N258 , \u_cordic/mycordic/N257 ,
         \u_cordic/mycordic/N256 , \u_cordic/mycordic/N255 ,
         \u_cordic/mycordic/N247 , \u_cordic/mycordic/N246 ,
         \u_cordic/mycordic/N245 , \u_cordic/mycordic/N244 ,
         \u_cordic/mycordic/N238 , \u_cordic/mycordic/N237 ,
         \u_cordic/mycordic/N236 , \u_cordic/mycordic/N212 ,
         \u_cordic/mycordic/N211 , \u_cordic/mycordic/N44 ,
         \u_cordic/mycordic/next_ANGLE_table[6][15] ,
         \u_cordic/mycordic/next_ANGLE_table[6][14] ,
         \u_cordic/mycordic/next_ANGLE_table[6][13] ,
         \u_cordic/mycordic/next_ANGLE_table[6][12] ,
         \u_cordic/mycordic/next_ANGLE_table[6][11] ,
         \u_cordic/mycordic/next_ANGLE_table[6][10] ,
         \u_cordic/mycordic/next_ANGLE_table[6][9] ,
         \u_cordic/mycordic/next_ANGLE_table[6][8] ,
         \u_cordic/mycordic/next_ANGLE_table[6][7] ,
         \u_cordic/mycordic/next_ANGLE_table[6][6] ,
         \u_cordic/mycordic/next_ANGLE_table[6][5] ,
         \u_cordic/mycordic/next_ANGLE_table[6][4] ,
         \u_cordic/mycordic/next_ANGLE_table[6][3] ,
         \u_cordic/mycordic/next_ANGLE_table[6][2] ,
         \u_cordic/mycordic/next_ANGLE_table[6][1] ,
         \u_cordic/mycordic/next_ANGLE_table[6][0] ,
         \u_cordic/mycordic/present_C_table[1][0] ,
         \u_cordic/mycordic/present_C_table[1][1] ,
         \u_cordic/mycordic/present_C_table[1][2] ,
         \u_cordic/mycordic/present_C_table[2][0] ,
         \u_cordic/mycordic/present_C_table[2][1] ,
         \u_cordic/mycordic/present_C_table[2][2] ,
         \u_cordic/mycordic/present_C_table[3][0] ,
         \u_cordic/mycordic/present_C_table[3][1] ,
         \u_cordic/mycordic/present_C_table[3][2] ,
         \u_cordic/mycordic/present_C_table[4][0] ,
         \u_cordic/mycordic/present_C_table[4][1] ,
         \u_cordic/mycordic/present_C_table[4][2] ,
         \u_cordic/mycordic/present_C_table[5][0] ,
         \u_cordic/mycordic/present_C_table[5][1] ,
         \u_cordic/mycordic/present_C_table[5][2] ,
         \u_cordic/mycordic/present_C_table[6][0] ,
         \u_cordic/mycordic/present_C_table[6][1] ,
         \u_cordic/mycordic/present_C_table[6][2] ,
         \u_cordic/mycordic/present_C_table[7][0] ,
         \u_cordic/mycordic/present_C_table[7][1] ,
         \u_cordic/mycordic/present_ANGLE_table[6][15] ,
         \u_cordic/mycordic/present_ANGLE_table[6][14] ,
         \u_cordic/mycordic/present_ANGLE_table[6][13] ,
         \u_cordic/mycordic/present_ANGLE_table[6][12] ,
         \u_cordic/mycordic/present_ANGLE_table[6][11] ,
         \u_cordic/mycordic/present_ANGLE_table[6][10] ,
         \u_cordic/mycordic/present_ANGLE_table[6][9] ,
         \u_cordic/mycordic/present_ANGLE_table[6][8] ,
         \u_cordic/mycordic/present_ANGLE_table[6][7] ,
         \u_cordic/mycordic/present_ANGLE_table[6][6] ,
         \u_cordic/mycordic/present_ANGLE_table[6][5] ,
         \u_cordic/mycordic/present_ANGLE_table[6][4] ,
         \u_cordic/mycordic/present_ANGLE_table[6][3] ,
         \u_cordic/mycordic/present_ANGLE_table[6][2] ,
         \u_cordic/mycordic/present_ANGLE_table[6][1] ,
         \u_cordic/mycordic/present_ANGLE_table[5][15] ,
         \u_cordic/mycordic/present_ANGLE_table[5][14] ,
         \u_cordic/mycordic/present_ANGLE_table[5][13] ,
         \u_cordic/mycordic/present_ANGLE_table[5][12] ,
         \u_cordic/mycordic/present_ANGLE_table[5][11] ,
         \u_cordic/mycordic/present_ANGLE_table[5][10] ,
         \u_cordic/mycordic/present_ANGLE_table[5][9] ,
         \u_cordic/mycordic/present_ANGLE_table[5][8] ,
         \u_cordic/mycordic/present_ANGLE_table[5][7] ,
         \u_cordic/mycordic/present_ANGLE_table[5][6] ,
         \u_cordic/mycordic/present_ANGLE_table[5][5] ,
         \u_cordic/mycordic/present_ANGLE_table[5][4] ,
         \u_cordic/mycordic/present_ANGLE_table[5][3] ,
         \u_cordic/mycordic/present_ANGLE_table[5][2] ,
         \u_cordic/mycordic/present_ANGLE_table[5][1] ,
         \u_cordic/mycordic/present_ANGLE_table[4][15] ,
         \u_cordic/mycordic/present_ANGLE_table[4][14] ,
         \u_cordic/mycordic/present_ANGLE_table[4][13] ,
         \u_cordic/mycordic/present_ANGLE_table[4][12] ,
         \u_cordic/mycordic/present_ANGLE_table[4][11] ,
         \u_cordic/mycordic/present_ANGLE_table[4][10] ,
         \u_cordic/mycordic/present_ANGLE_table[4][9] ,
         \u_cordic/mycordic/present_ANGLE_table[4][8] ,
         \u_cordic/mycordic/present_ANGLE_table[4][7] ,
         \u_cordic/mycordic/present_ANGLE_table[4][6] ,
         \u_cordic/mycordic/present_ANGLE_table[4][5] ,
         \u_cordic/mycordic/present_ANGLE_table[4][4] ,
         \u_cordic/mycordic/present_ANGLE_table[4][3] ,
         \u_cordic/mycordic/present_ANGLE_table[4][2] ,
         \u_cordic/mycordic/present_ANGLE_table[4][1] ,
         \u_cordic/mycordic/present_ANGLE_table[4][0] ,
         \u_cordic/mycordic/present_ANGLE_table[3][15] ,
         \u_cordic/mycordic/present_ANGLE_table[3][14] ,
         \u_cordic/mycordic/present_ANGLE_table[3][13] ,
         \u_cordic/mycordic/present_ANGLE_table[3][12] ,
         \u_cordic/mycordic/present_ANGLE_table[3][11] ,
         \u_cordic/mycordic/present_ANGLE_table[3][10] ,
         \u_cordic/mycordic/present_ANGLE_table[3][9] ,
         \u_cordic/mycordic/present_ANGLE_table[3][8] ,
         \u_cordic/mycordic/present_ANGLE_table[3][7] ,
         \u_cordic/mycordic/present_ANGLE_table[3][6] ,
         \u_cordic/mycordic/present_ANGLE_table[3][5] ,
         \u_cordic/mycordic/present_ANGLE_table[3][4] ,
         \u_cordic/mycordic/present_ANGLE_table[3][3] ,
         \u_cordic/mycordic/present_ANGLE_table[3][2] ,
         \u_cordic/mycordic/present_ANGLE_table[3][1] ,
         \u_cordic/mycordic/present_ANGLE_table[3][0] ,
         \u_cordic/mycordic/present_ANGLE_table[2][15] ,
         \u_cordic/mycordic/present_ANGLE_table[2][14] ,
         \u_cordic/mycordic/present_ANGLE_table[2][13] ,
         \u_cordic/mycordic/present_ANGLE_table[2][12] ,
         \u_cordic/mycordic/present_ANGLE_table[2][11] ,
         \u_cordic/mycordic/present_ANGLE_table[2][10] ,
         \u_cordic/mycordic/present_ANGLE_table[2][9] ,
         \u_cordic/mycordic/present_ANGLE_table[2][8] ,
         \u_cordic/mycordic/present_ANGLE_table[2][7] ,
         \u_cordic/mycordic/present_ANGLE_table[2][6] ,
         \u_cordic/mycordic/present_ANGLE_table[2][5] ,
         \u_cordic/mycordic/present_ANGLE_table[2][4] ,
         \u_cordic/mycordic/present_ANGLE_table[2][3] ,
         \u_cordic/mycordic/present_ANGLE_table[2][2] ,
         \u_cordic/mycordic/present_ANGLE_table[2][1] ,
         \u_cordic/mycordic/present_ANGLE_table[1][15] ,
         \u_cordic/mycordic/present_ANGLE_table[1][14] ,
         \u_cordic/mycordic/present_ANGLE_table[1][13] ,
         \u_cordic/mycordic/present_ANGLE_table[1][12] ,
         \u_cordic/mycordic/present_ANGLE_table[1][11] ,
         \u_cordic/mycordic/present_ANGLE_table[1][10] ,
         \u_cordic/mycordic/present_ANGLE_table[1][9] ,
         \u_cordic/mycordic/present_ANGLE_table[1][8] ,
         \u_cordic/mycordic/present_ANGLE_table[1][7] ,
         \u_cordic/mycordic/present_ANGLE_table[1][6] ,
         \u_cordic/mycordic/present_ANGLE_table[1][5] ,
         \u_cordic/mycordic/present_ANGLE_table[1][4] ,
         \u_cordic/mycordic/present_ANGLE_table[1][3] ,
         \u_cordic/mycordic/present_ANGLE_table[1][2] ,
         \u_cordic/mycordic/present_ANGLE_table[1][1] ,
         \u_cordic/mycordic/present_ANGLE_table[1][0] ,
         \u_cordic/mycordic/present_Q_table[0][3] ,
         \u_cordic/mycordic/present_Q_table[0][4] ,
         \u_cordic/mycordic/present_Q_table[0][5] ,
         \u_cordic/mycordic/present_Q_table[0][6] ,
         \u_cordic/mycordic/present_Q_table[0][7] ,
         \u_cordic/mycordic/present_Q_table[1][3] ,
         \u_cordic/mycordic/present_Q_table[1][4] ,
         \u_cordic/mycordic/present_Q_table[1][5] ,
         \u_cordic/mycordic/present_Q_table[1][6] ,
         \u_cordic/mycordic/present_Q_table[1][7] ,
         \u_cordic/mycordic/present_Q_table[2][0] ,
         \u_cordic/mycordic/present_Q_table[2][1] ,
         \u_cordic/mycordic/present_Q_table[2][2] ,
         \u_cordic/mycordic/present_Q_table[2][3] ,
         \u_cordic/mycordic/present_Q_table[2][4] ,
         \u_cordic/mycordic/present_Q_table[2][5] ,
         \u_cordic/mycordic/present_Q_table[2][6] ,
         \u_cordic/mycordic/present_Q_table[2][7] ,
         \u_cordic/mycordic/present_Q_table[3][0] ,
         \u_cordic/mycordic/present_Q_table[3][1] ,
         \u_cordic/mycordic/present_Q_table[3][2] ,
         \u_cordic/mycordic/present_Q_table[3][3] ,
         \u_cordic/mycordic/present_Q_table[3][4] ,
         \u_cordic/mycordic/present_Q_table[3][5] ,
         \u_cordic/mycordic/present_Q_table[3][6] ,
         \u_cordic/mycordic/present_Q_table[3][7] ,
         \u_cordic/mycordic/present_Q_table[4][0] ,
         \u_cordic/mycordic/present_Q_table[4][1] ,
         \u_cordic/mycordic/present_Q_table[4][2] ,
         \u_cordic/mycordic/present_Q_table[4][3] ,
         \u_cordic/mycordic/present_Q_table[4][4] ,
         \u_cordic/mycordic/present_Q_table[4][5] ,
         \u_cordic/mycordic/present_Q_table[4][6] ,
         \u_cordic/mycordic/present_Q_table[4][7] ,
         \u_cordic/mycordic/present_Q_table[5][0] ,
         \u_cordic/mycordic/present_Q_table[5][1] ,
         \u_cordic/mycordic/present_Q_table[5][2] ,
         \u_cordic/mycordic/present_Q_table[5][3] ,
         \u_cordic/mycordic/present_Q_table[5][4] ,
         \u_cordic/mycordic/present_Q_table[5][5] ,
         \u_cordic/mycordic/present_Q_table[5][6] ,
         \u_cordic/mycordic/present_Q_table[5][7] ,
         \u_cordic/mycordic/present_Q_table[6][7] ,
         \u_cordic/mycordic/present_I_table[0][3] ,
         \u_cordic/mycordic/present_I_table[0][4] ,
         \u_cordic/mycordic/present_I_table[0][5] ,
         \u_cordic/mycordic/present_I_table[0][6] ,
         \u_cordic/mycordic/present_I_table[0][7] ,
         \u_cordic/mycordic/present_I_table[1][3] ,
         \u_cordic/mycordic/present_I_table[1][4] ,
         \u_cordic/mycordic/present_I_table[1][5] ,
         \u_cordic/mycordic/present_I_table[1][6] ,
         \u_cordic/mycordic/present_I_table[1][7] ,
         \u_cordic/mycordic/present_I_table[2][0] ,
         \u_cordic/mycordic/present_I_table[2][1] ,
         \u_cordic/mycordic/present_I_table[2][2] ,
         \u_cordic/mycordic/present_I_table[2][3] ,
         \u_cordic/mycordic/present_I_table[2][4] ,
         \u_cordic/mycordic/present_I_table[2][5] ,
         \u_cordic/mycordic/present_I_table[2][6] ,
         \u_cordic/mycordic/present_I_table[2][7] ,
         \u_cordic/mycordic/present_I_table[3][0] ,
         \u_cordic/mycordic/present_I_table[3][1] ,
         \u_cordic/mycordic/present_I_table[3][2] ,
         \u_cordic/mycordic/present_I_table[3][3] ,
         \u_cordic/mycordic/present_I_table[3][4] ,
         \u_cordic/mycordic/present_I_table[3][5] ,
         \u_cordic/mycordic/present_I_table[3][6] ,
         \u_cordic/mycordic/present_I_table[3][7] ,
         \u_cordic/mycordic/present_I_table[4][0] ,
         \u_cordic/mycordic/present_I_table[4][1] ,
         \u_cordic/mycordic/present_I_table[4][2] ,
         \u_cordic/mycordic/present_I_table[4][3] ,
         \u_cordic/mycordic/present_I_table[4][4] ,
         \u_cordic/mycordic/present_I_table[4][5] ,
         \u_cordic/mycordic/present_I_table[4][6] ,
         \u_cordic/mycordic/present_I_table[4][7] ,
         \u_cordic/mycordic/present_I_table[5][4] ,
         \u_cordic/mycordic/present_I_table[5][5] ,
         \u_cordic/mycordic/present_I_table[5][6] ,
         \u_cordic/mycordic/present_I_table[5][7] , \u_cordic/my_rotation/n85 ,
         \u_cordic/my_rotation/n84 , \u_cordic/my_rotation/n83 ,
         \u_cordic/my_rotation/n82 , \u_cordic/my_rotation/n81 ,
         \u_cordic/my_rotation/n80 , \u_cordic/my_rotation/n79 ,
         \u_cordic/my_rotation/n78 , \u_cordic/my_rotation/n77 ,
         \u_cordic/my_rotation/n76 , \u_cordic/my_rotation/n75 ,
         \u_cordic/my_rotation/n74 , \u_cordic/my_rotation/n73 ,
         \u_cordic/my_rotation/n72 , \u_cordic/my_rotation/n71 ,
         \u_cordic/my_rotation/n70 , \u_cordic/my_rotation/n69 ,
         \u_cordic/my_rotation/n68 , \u_cordic/my_rotation/n67 ,
         \u_cordic/my_rotation/n66 , \u_cordic/my_rotation/n65 ,
         \u_cordic/my_rotation/n64 , \u_cordic/my_rotation/n63 ,
         \u_cordic/my_rotation/n62 , \u_cordic/my_rotation/n61 ,
         \u_cordic/my_rotation/n60 , \u_cordic/my_rotation/n59 ,
         \u_cordic/my_rotation/n58 , \u_cordic/my_rotation/n57 ,
         \u_cordic/my_rotation/n56 , \u_cordic/my_rotation/n55 ,
         \u_cordic/my_rotation/n54 , \u_cordic/my_rotation/n53 ,
         \u_cordic/my_rotation/n52 , \u_cordic/my_rotation/n51 ,
         \u_cordic/my_rotation/n50 , \u_cordic/my_rotation/n49 ,
         \u_cordic/my_rotation/n48 , \u_cordic/my_rotation/n47 ,
         \u_cordic/my_rotation/N40 , \u_cordic/my_rotation/N39 ,
         \u_cordic/my_rotation/N38 , \u_cordic/my_rotation/N37 ,
         \u_cordic/my_rotation/N36 , \u_cordic/my_rotation/N35 ,
         \u_cordic/my_rotation/N34 , \u_cordic/my_rotation/N33 ,
         \u_cordic/my_rotation/N32 , \u_cordic/my_rotation/N31 ,
         \u_cordic/my_rotation/N30 , \u_cordic/my_rotation/N29 ,
         \u_cordic/my_rotation/N25 , \u_cordic/my_rotation/N23 ,
         \u_cordic/my_rotation/present_angle[0][15] ,
         \u_cordic/my_rotation/present_angle[0][14] ,
         \u_cordic/my_rotation/present_angle[0][13] ,
         \u_cordic/my_rotation/present_angle[0][12] ,
         \u_cordic/my_rotation/present_angle[0][11] ,
         \u_cordic/my_rotation/present_angle[0][10] ,
         \u_cordic/my_rotation/present_angle[0][9] ,
         \u_cordic/my_rotation/present_angle[0][8] ,
         \u_cordic/my_rotation/present_angle[0][7] ,
         \u_cordic/my_rotation/present_angle[0][6] ,
         \u_cordic/my_rotation/present_angle[0][5] ,
         \u_cordic/my_rotation/present_angle[0][4] ,
         \u_cordic/my_rotation/present_angle[0][3] ,
         \u_cordic/my_rotation/present_angle[0][2] ,
         \u_cordic/my_rotation/present_angle[0][1] ,
         \u_cordic/my_rotation/present_angle[0][0] , \u_cdr/div1/n40 ,
         \u_cdr/div1/n39 , \u_cdr/div1/n38 , \u_cdr/div1/n37 ,
         \u_cdr/div1/n36 , \u_cdr/div1/n35 , \u_cdr/div1/n32 ,
         \u_cdr/div1/n31 , \u_cdr/div1/n27 , \u_cdr/div1/n10 , \u_cdr/div1/n9 ,
         \u_cdr/div1/n8 , \u_cdr/div1/n7 , \u_cdr/div1/N35 ,
         \u_cdr/div1/w_en_freq_synch , \u_cdr/phd1/n23 , \u_cdr/phd1/n22 ,
         \u_cdr/phd1/n21 , \u_cdr/phd1/n20 , \u_cdr/phd1/n19 ,
         \u_cdr/phd1/n18 , \u_cdr/phd1/n17 , \u_cdr/phd1/n16 ,
         \u_cdr/phd1/n15 , \u_cdr/phd1/n14 , \u_cdr/phd1/n13 ,
         \u_cdr/phd1/n12 , \u_cdr/phd1/n11 , \u_cdr/phd1/w_s4 ,
         \u_cdr/phd1/w_s3 , \u_cdr/phd1/w_s2 , \u_cdr/phd1/w_s1 ,
         \u_cdr/phd1/w_en_f , \u_cdr/phd1/w_en_m , \u_cdr/phd1/w_en_d ,
         \u_cdr/dec1/n33 , \u_cdr/dec1/n32 , \u_cdr/dec1/n31 ,
         \u_cdr/dec1/n30 , \u_cdr/dec1/n29 , \u_cdr/dec1/n26 ,
         \u_cdr/dec1/n25 , \u_cdr/dec1/n24 , \u_cdr/dec1/n20 ,
         \u_cdr/dec1/w_en_dec , \u_cdr/dec1/N73 , \u_cdr/dec1/N65 ,
         \u_cdr/dec1/N64 , \u_cdr/dec1/N63 , \u_cdr/dec1/N62 ,
         \u_cdr/dec1/N61 , \u_cdr/dec1/w_s_r , \u_inFIFO/os1/dff1/n2 ,
         \u_decoder/iq_demod/cossin_dig/n56 ,
         \u_decoder/iq_demod/cossin_dig/n55 ,
         \u_decoder/iq_demod/cossin_dig/n54 ,
         \u_decoder/iq_demod/cossin_dig/n53 ,
         \u_decoder/iq_demod/cossin_dig/n52 ,
         \u_decoder/iq_demod/cossin_dig/n51 ,
         \u_decoder/iq_demod/cossin_dig/n50 ,
         \u_decoder/iq_demod/cossin_dig/n49 ,
         \u_decoder/iq_demod/cossin_dig/n48 ,
         \u_decoder/iq_demod/cossin_dig/n47 ,
         \u_decoder/iq_demod/cossin_dig/n46 ,
         \u_decoder/iq_demod/cossin_dig/n45 ,
         \u_decoder/iq_demod/cossin_dig/n44 ,
         \u_decoder/iq_demod/cossin_dig/n43 ,
         \u_decoder/iq_demod/cossin_dig/n42 ,
         \u_decoder/iq_demod/cossin_dig/n41 ,
         \u_decoder/iq_demod/cossin_dig/n40 ,
         \u_decoder/iq_demod/cossin_dig/n39 ,
         \u_decoder/iq_demod/cossin_dig/n38 ,
         \u_decoder/iq_demod/cossin_dig/n37 ,
         \u_decoder/iq_demod/cossin_dig/n36 ,
         \u_decoder/iq_demod/cossin_dig/n35 ,
         \u_decoder/iq_demod/cossin_dig/n34 ,
         \u_decoder/iq_demod/cossin_dig/n33 ,
         \u_decoder/iq_demod/cossin_dig/n32 ,
         \u_decoder/iq_demod/cossin_dig/n31 ,
         \u_decoder/iq_demod/cossin_dig/n30 ,
         \u_decoder/iq_demod/cossin_dig/n29 ,
         \u_decoder/iq_demod/cossin_dig/n28 ,
         \u_decoder/iq_demod/cossin_dig/n27 ,
         \u_decoder/iq_demod/cossin_dig/n26 ,
         \u_decoder/iq_demod/cossin_dig/n25 ,
         \u_decoder/iq_demod/cossin_dig/n23 ,
         \u_decoder/iq_demod/cossin_dig/n21 ,
         \u_decoder/iq_demod/cossin_dig/n19 ,
         \u_decoder/iq_demod/cossin_dig/n10 ,
         \u_decoder/iq_demod/cossin_dig/N60 ,
         \u_decoder/iq_demod/cossin_dig/N55 ,
         \u_decoder/iq_demod/cossin_dig/N52 ,
         \u_decoder/iq_demod/cossin_dig/N42 ,
         \u_decoder/iq_demod/cossin_dig/N41 ,
         \u_decoder/iq_demod/cossin_dig/N22 ,
         \u_decoder/iq_demod/cossin_dig/N21 ,
         \u_decoder/iq_demod/cossin_dig/N20 ,
         \u_decoder/iq_demod/cossin_dig/state[0] , \u_cdr/div1/cnt_div/n41 ,
         \u_cdr/div1/cnt_div/n40 , \u_cdr/div1/cnt_div/n39 ,
         \u_cdr/div1/cnt_div/n38 , \u_cdr/div1/cnt_div/n37 ,
         \u_cdr/div1/cnt_div/n36 , \u_cdr/div1/cnt_div/n35 ,
         \u_cdr/div1/cnt_div/n34 , \u_cdr/div1/cnt_div/n33 ,
         \u_cdr/div1/cnt_div/N88 , \u_cdr/div1/cnt_div/N76 ,
         \u_cdr/div1/cnt_div/N75 , \u_cdr/div1/cnt_div/N74 ,
         \u_cdr/div1/cnt_div/N73 , \u_cdr/div1/cnt_div/N72 ,
         \u_cdr/phd1/f1/n2 , \u_cdr/dec1/cnt_dec/n24 ,
         \u_cdr/dec1/cnt_dec/n23 , \u_cdr/dec1/cnt_dec/n22 ,
         \u_cdr/dec1/cnt_dec/n21 , \u_cdr/dec1/cnt_dec/n20 ,
         \u_cdr/dec1/cnt_dec/n19 , \u_cdr/dec1/cnt_dec/n18 ,
         \u_cdr/dec1/cnt_dec/n17 , \u_cdr/dec1/cnt_dec/n16 ,
         \u_cdr/dec1/cnt_dec/N33 , \u_cdr/dec1/cnt_dec/N9 ,
         \u_cdr/dec1/cnt_dec/N8 , \u_cdr/dec1/cnt_dec/N7 ,
         \u_cdr/dec1/cnt_dec/N6 , \u_cdr/dec1/cnt_dec/N5 ,
         \u_outFIFO/os2/sigQout2 , \u_outFIFO/os2/sigQout1 ,
         \u_outFIFO/os1/sigQout2 , \u_outFIFO/os1/sigQout1 ,
         \u_inFIFO/os2/sigQout2 , \u_inFIFO/os2/sigQout1 ,
         \u_cdr/phd1/cnt_phd/N84 , \u_cdr/phd1/cnt_phd/N76 ,
         \u_cdr/phd1/cnt_phd/N75 , \u_cdr/phd1/cnt_phd/N74 ,
         \u_cdr/phd1/cnt_phd/N73 , \u_cdr/phd1/cnt_phd/N72 ,
         \u_cdr/phd1/cnt_phd/N58 , \u_cdr/phd1/cnt_phd/N50 ,
         \u_cdr/phd1/cnt_phd/N42 , \u_cdr/phd1/cnt_phd/N41 ,
         \u_cdr/phd1/cnt_phd/N14 , \u_cdr/phd1/cnt_phd/N13 ,
         \u_cdr/phd1/cnt_phd/N12 , \u_cordic/mycordic/add_191/carry[2] ,
         \u_cordic/mycordic/add_191/carry[3] ,
         \u_cordic/mycordic/add_191/carry[4] ,
         \u_cordic/mycordic/add_191/carry[5] ,
         \u_cordic/mycordic/add_191/carry[6] ,
         \u_cordic/mycordic/add_191/carry[7] ,
         \u_cordic/mycordic/add_191/carry[8] ,
         \u_cordic/mycordic/add_191/carry[9] ,
         \u_cordic/mycordic/add_191/carry[10] ,
         \u_cordic/mycordic/add_191/carry[11] ,
         \u_cordic/mycordic/add_191/carry[12] ,
         \u_cordic/mycordic/add_191/carry[13] ,
         \u_cordic/mycordic/add_191/carry[14] ,
         \u_cordic/mycordic/add_191/carry[15] ,
         \u_cordic/mycordic/sub_196/carry[2] ,
         \u_cordic/mycordic/sub_196/carry[3] ,
         \u_cordic/mycordic/sub_196/carry[4] ,
         \u_cordic/mycordic/sub_196/carry[5] ,
         \u_cordic/mycordic/sub_196/carry[6] ,
         \u_cordic/mycordic/sub_196/carry[7] ,
         \u_cordic/mycordic/sub_196/carry[8] ,
         \u_cordic/mycordic/sub_196/carry[9] ,
         \u_cordic/mycordic/sub_196/carry[10] ,
         \u_cordic/mycordic/sub_196/carry[11] ,
         \u_cordic/mycordic/sub_196/carry[12] ,
         \u_cordic/mycordic/sub_196/carry[13] ,
         \u_cordic/mycordic/sub_196/carry[14] ,
         \u_cordic/mycordic/sub_196/carry[15] ,
         \u_cordic/mycordic/add_213/carry[2] ,
         \u_cordic/mycordic/add_213/carry[3] ,
         \u_cordic/mycordic/add_213/carry[4] ,
         \u_cordic/mycordic/add_213/carry[5] ,
         \u_cordic/mycordic/add_213/carry[6] ,
         \u_cordic/mycordic/add_213/carry[7] ,
         \u_cordic/mycordic/add_213/carry[8] ,
         \u_cordic/mycordic/add_213/carry[9] ,
         \u_cordic/mycordic/add_213/carry[10] ,
         \u_cordic/mycordic/add_213/carry[11] ,
         \u_cordic/mycordic/add_213/carry[12] ,
         \u_cordic/mycordic/add_213/carry[13] ,
         \u_cordic/mycordic/add_213/carry[14] ,
         \u_cordic/mycordic/add_213/carry[15] ,
         \u_cordic/mycordic/sub_218/carry[2] ,
         \u_cordic/mycordic/sub_218/carry[3] ,
         \u_cordic/mycordic/sub_218/carry[4] ,
         \u_cordic/mycordic/sub_218/carry[5] ,
         \u_cordic/mycordic/sub_218/carry[6] ,
         \u_cordic/mycordic/sub_218/carry[7] ,
         \u_cordic/mycordic/sub_218/carry[8] ,
         \u_cordic/mycordic/sub_218/carry[9] ,
         \u_cordic/mycordic/sub_218/carry[10] ,
         \u_cordic/mycordic/sub_218/carry[11] ,
         \u_cordic/mycordic/sub_218/carry[12] ,
         \u_cordic/mycordic/sub_218/carry[13] ,
         \u_cordic/mycordic/sub_218/carry[14] ,
         \u_cordic/mycordic/sub_218/carry[15] ,
         \u_cordic/mycordic/sub_223/carry[7] ,
         \u_cordic/mycordic/add_224/carry[2] ,
         \u_cordic/mycordic/add_224/carry[3] ,
         \u_cordic/mycordic/add_224/carry[4] ,
         \u_cordic/mycordic/add_224/carry[5] ,
         \u_cordic/mycordic/add_224/carry[6] ,
         \u_cordic/mycordic/add_224/carry[7] ,
         \u_cordic/mycordic/add_224/carry[8] ,
         \u_cordic/mycordic/add_224/carry[9] ,
         \u_cordic/mycordic/add_224/carry[10] ,
         \u_cordic/mycordic/add_224/carry[11] ,
         \u_cordic/mycordic/add_224/carry[12] ,
         \u_cordic/mycordic/add_224/carry[13] ,
         \u_cordic/mycordic/add_224/carry[14] ,
         \u_cordic/mycordic/add_224/carry[15] ,
         \u_cordic/mycordic/add_228/carry[7] ,
         \u_cordic/mycordic/sub_229/carry[2] ,
         \u_cordic/mycordic/sub_229/carry[3] ,
         \u_cordic/mycordic/sub_229/carry[4] ,
         \u_cordic/mycordic/sub_229/carry[5] ,
         \u_cordic/mycordic/sub_229/carry[6] ,
         \u_cordic/mycordic/sub_229/carry[7] ,
         \u_cordic/mycordic/sub_229/carry[8] ,
         \u_cordic/mycordic/sub_229/carry[9] ,
         \u_cordic/mycordic/sub_229/carry[10] ,
         \u_cordic/mycordic/sub_229/carry[11] ,
         \u_cordic/mycordic/sub_229/carry[12] ,
         \u_cordic/mycordic/sub_229/carry[13] ,
         \u_cordic/mycordic/sub_229/carry[14] ,
         \u_cordic/mycordic/sub_229/carry[15] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_276/A2[7] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_276/A2[8] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_276/A2[9] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_276/A2[10] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_276/A2[11] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_276/A1[7] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_276/A1[8] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_276/A1[9] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_276/A1[10] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_276/SUMB[1][5] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_276/SUMB[2][3] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_276/SUMB[2][5] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_276/SUMB[3][3] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_276/SUMB[3][5] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_276/SUMB[4][3] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_276/SUMB[4][5] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_276/SUMB[5][3] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_276/SUMB[5][5] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_276/SUMB[6][3] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_276/SUMB[6][5] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_276/SUMB[7][0] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_276/SUMB[7][1] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_276/SUMB[7][2] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_276/SUMB[7][3] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_276/SUMB[7][4] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_276/SUMB[7][5] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[1][5] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[2][3] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[2][5] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[3][0] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[3][3] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[3][5] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[4][0] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[4][3] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[4][5] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[5][0] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[5][3] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[5][5] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[6][0] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[6][3] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[6][5] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[7][0] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[7][1] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[7][2] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[7][3] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[7][4] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[7][5] ,
         \u_decoder/fir_filter/dp_cluster_0/r167/A2[7] ,
         \u_decoder/fir_filter/dp_cluster_0/r167/A2[8] ,
         \u_decoder/fir_filter/dp_cluster_0/r167/A2[9] ,
         \u_decoder/fir_filter/dp_cluster_0/r167/A2[10] ,
         \u_decoder/fir_filter/dp_cluster_0/r167/A2[11] ,
         \u_decoder/fir_filter/dp_cluster_0/r167/A1[7] ,
         \u_decoder/fir_filter/dp_cluster_0/r167/A1[8] ,
         \u_decoder/fir_filter/dp_cluster_0/r167/A1[9] ,
         \u_decoder/fir_filter/dp_cluster_0/r167/A1[10] ,
         \u_decoder/fir_filter/dp_cluster_0/r167/SUMB[2][1] ,
         \u_decoder/fir_filter/dp_cluster_0/r167/SUMB[3][1] ,
         \u_decoder/fir_filter/dp_cluster_0/r167/SUMB[3][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r167/SUMB[4][1] ,
         \u_decoder/fir_filter/dp_cluster_0/r167/SUMB[4][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r167/SUMB[5][1] ,
         \u_decoder/fir_filter/dp_cluster_0/r167/SUMB[5][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r167/SUMB[6][1] ,
         \u_decoder/fir_filter/dp_cluster_0/r167/SUMB[6][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r167/SUMB[7][0] ,
         \u_decoder/fir_filter/dp_cluster_0/r167/SUMB[7][1] ,
         \u_decoder/fir_filter/dp_cluster_0/r167/SUMB[7][2] ,
         \u_decoder/fir_filter/dp_cluster_0/r167/SUMB[7][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r167/SUMB[7][4] ,
         \u_decoder/fir_filter/dp_cluster_0/r167/SUMB[7][5] ,
         \u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[1][0] ,
         \u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[2][0] ,
         \u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[2][1] ,
         \u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[3][0] ,
         \u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[3][1] ,
         \u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[3][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[4][0] ,
         \u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[4][1] ,
         \u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[4][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[5][0] ,
         \u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[5][1] ,
         \u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[5][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[6][0] ,
         \u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[6][1] ,
         \u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[6][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[7][0] ,
         \u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[7][1] ,
         \u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[7][2] ,
         \u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[7][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[7][4] ,
         \u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[7][5] ,
         \u_decoder/fir_filter/dp_cluster_0/r166/A2[6] ,
         \u_decoder/fir_filter/dp_cluster_0/r166/A2[7] ,
         \u_decoder/fir_filter/dp_cluster_0/r166/A2[8] ,
         \u_decoder/fir_filter/dp_cluster_0/r166/A2[9] ,
         \u_decoder/fir_filter/dp_cluster_0/r166/A1[6] ,
         \u_decoder/fir_filter/dp_cluster_0/r166/A1[7] ,
         \u_decoder/fir_filter/dp_cluster_0/r166/A1[8] ,
         \u_decoder/fir_filter/dp_cluster_0/r166/SUMB[1][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r166/SUMB[2][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r166/SUMB[3][1] ,
         \u_decoder/fir_filter/dp_cluster_0/r166/SUMB[3][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r166/SUMB[4][1] ,
         \u_decoder/fir_filter/dp_cluster_0/r166/SUMB[4][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r166/SUMB[5][1] ,
         \u_decoder/fir_filter/dp_cluster_0/r166/SUMB[5][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r166/SUMB[6][1] ,
         \u_decoder/fir_filter/dp_cluster_0/r166/SUMB[6][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r166/SUMB[7][0] ,
         \u_decoder/fir_filter/dp_cluster_0/r166/SUMB[7][1] ,
         \u_decoder/fir_filter/dp_cluster_0/r166/SUMB[7][2] ,
         \u_decoder/fir_filter/dp_cluster_0/r166/SUMB[7][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r166/CARRYB[1][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r166/CARRYB[2][1] ,
         \u_decoder/fir_filter/dp_cluster_0/r166/CARRYB[2][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r166/CARRYB[3][1] ,
         \u_decoder/fir_filter/dp_cluster_0/r166/CARRYB[3][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r166/CARRYB[4][1] ,
         \u_decoder/fir_filter/dp_cluster_0/r166/CARRYB[4][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r166/CARRYB[5][1] ,
         \u_decoder/fir_filter/dp_cluster_0/r166/CARRYB[5][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r166/CARRYB[6][1] ,
         \u_decoder/fir_filter/dp_cluster_0/r166/CARRYB[6][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r166/CARRYB[7][0] ,
         \u_decoder/fir_filter/dp_cluster_0/r166/CARRYB[7][1] ,
         \u_decoder/fir_filter/dp_cluster_0/r166/CARRYB[7][2] ,
         \u_decoder/fir_filter/dp_cluster_0/r166/CARRYB[7][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r165/A2[6] ,
         \u_decoder/fir_filter/dp_cluster_0/r165/A2[7] ,
         \u_decoder/fir_filter/dp_cluster_0/r165/A2[8] ,
         \u_decoder/fir_filter/dp_cluster_0/r165/A2[9] ,
         \u_decoder/fir_filter/dp_cluster_0/r165/A2[10] ,
         \u_decoder/fir_filter/dp_cluster_0/r165/A1[4] ,
         \u_decoder/fir_filter/dp_cluster_0/r165/A1[5] ,
         \u_decoder/fir_filter/dp_cluster_0/r165/A1[6] ,
         \u_decoder/fir_filter/dp_cluster_0/r165/A1[7] ,
         \u_decoder/fir_filter/dp_cluster_0/r165/A1[8] ,
         \u_decoder/fir_filter/dp_cluster_0/r165/A1[9] ,
         \u_decoder/fir_filter/dp_cluster_0/r165/PROD1[5] ,
         \u_decoder/fir_filter/dp_cluster_0/r165/SUMB[2][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r165/SUMB[3][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r165/SUMB[4][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r165/SUMB[5][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r165/SUMB[6][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r165/SUMB[7][0] ,
         \u_decoder/fir_filter/dp_cluster_0/r165/SUMB[7][1] ,
         \u_decoder/fir_filter/dp_cluster_0/r165/SUMB[7][2] ,
         \u_decoder/fir_filter/dp_cluster_0/r165/SUMB[7][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r165/SUMB[7][4] ,
         \u_decoder/fir_filter/dp_cluster_0/r165/CARRYB[2][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r165/CARRYB[3][0] ,
         \u_decoder/fir_filter/dp_cluster_0/r165/CARRYB[3][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r165/CARRYB[4][0] ,
         \u_decoder/fir_filter/dp_cluster_0/r165/CARRYB[4][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r165/CARRYB[5][0] ,
         \u_decoder/fir_filter/dp_cluster_0/r165/CARRYB[5][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r165/CARRYB[6][0] ,
         \u_decoder/fir_filter/dp_cluster_0/r165/CARRYB[6][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r165/CARRYB[7][0] ,
         \u_decoder/fir_filter/dp_cluster_0/r165/CARRYB[7][1] ,
         \u_decoder/fir_filter/dp_cluster_0/r165/CARRYB[7][2] ,
         \u_decoder/fir_filter/dp_cluster_0/r165/CARRYB[7][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r165/CARRYB[7][4] ,
         \u_decoder/fir_filter/dp_cluster_0/r164/A2[6] ,
         \u_decoder/fir_filter/dp_cluster_0/r164/A2[7] ,
         \u_decoder/fir_filter/dp_cluster_0/r164/A2[8] ,
         \u_decoder/fir_filter/dp_cluster_0/r164/A2[9] ,
         \u_decoder/fir_filter/dp_cluster_0/r164/A1[3] ,
         \u_decoder/fir_filter/dp_cluster_0/r164/A1[4] ,
         \u_decoder/fir_filter/dp_cluster_0/r164/A1[5] ,
         \u_decoder/fir_filter/dp_cluster_0/r164/A1[6] ,
         \u_decoder/fir_filter/dp_cluster_0/r164/A1[7] ,
         \u_decoder/fir_filter/dp_cluster_0/r164/A1[8] ,
         \u_decoder/fir_filter/dp_cluster_0/r164/PROD1[4] ,
         \u_decoder/fir_filter/dp_cluster_0/r164/SUMB[2][2] ,
         \u_decoder/fir_filter/dp_cluster_0/r164/SUMB[3][2] ,
         \u_decoder/fir_filter/dp_cluster_0/r164/SUMB[4][2] ,
         \u_decoder/fir_filter/dp_cluster_0/r164/SUMB[5][2] ,
         \u_decoder/fir_filter/dp_cluster_0/r164/SUMB[6][2] ,
         \u_decoder/fir_filter/dp_cluster_0/r164/SUMB[7][0] ,
         \u_decoder/fir_filter/dp_cluster_0/r164/SUMB[7][1] ,
         \u_decoder/fir_filter/dp_cluster_0/r164/SUMB[7][2] ,
         \u_decoder/fir_filter/dp_cluster_0/r164/SUMB[7][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r164/CARRYB[2][0] ,
         \u_decoder/fir_filter/dp_cluster_0/r164/CARRYB[2][2] ,
         \u_decoder/fir_filter/dp_cluster_0/r164/CARRYB[3][0] ,
         \u_decoder/fir_filter/dp_cluster_0/r164/CARRYB[3][2] ,
         \u_decoder/fir_filter/dp_cluster_0/r164/CARRYB[4][0] ,
         \u_decoder/fir_filter/dp_cluster_0/r164/CARRYB[4][2] ,
         \u_decoder/fir_filter/dp_cluster_0/r164/CARRYB[5][0] ,
         \u_decoder/fir_filter/dp_cluster_0/r164/CARRYB[5][2] ,
         \u_decoder/fir_filter/dp_cluster_0/r164/CARRYB[6][0] ,
         \u_decoder/fir_filter/dp_cluster_0/r164/CARRYB[6][2] ,
         \u_decoder/fir_filter/dp_cluster_0/r164/CARRYB[7][0] ,
         \u_decoder/fir_filter/dp_cluster_0/r164/CARRYB[7][1] ,
         \u_decoder/fir_filter/dp_cluster_0/r164/CARRYB[7][2] ,
         \u_decoder/fir_filter/dp_cluster_0/r164/CARRYB[7][3] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_308/A2[7] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_308/A2[8] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_308/A2[9] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_308/A2[10] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_308/A2[11] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_308/A1[7] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_308/A1[8] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_308/A1[9] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_308/A1[10] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_308/SUMB[1][5] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_308/SUMB[2][3] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_308/SUMB[2][5] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_308/SUMB[3][3] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_308/SUMB[3][5] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_308/SUMB[4][3] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_308/SUMB[4][5] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_308/SUMB[5][3] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_308/SUMB[5][5] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_308/SUMB[6][3] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_308/SUMB[6][5] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_308/SUMB[7][0] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_308/SUMB[7][1] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_308/SUMB[7][2] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_308/SUMB[7][3] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_308/SUMB[7][4] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_308/SUMB[7][5] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[1][5] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[2][3] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[2][5] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[3][0] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[3][3] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[3][5] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[4][0] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[4][3] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[4][5] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[5][0] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[5][3] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[5][5] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[6][0] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[6][3] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[6][5] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[7][0] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[7][1] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[7][2] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[7][3] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[7][4] ,
         \u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[7][5] ,
         \u_decoder/fir_filter/dp_cluster_0/r180/A2[7] ,
         \u_decoder/fir_filter/dp_cluster_0/r180/A2[8] ,
         \u_decoder/fir_filter/dp_cluster_0/r180/A2[9] ,
         \u_decoder/fir_filter/dp_cluster_0/r180/A2[10] ,
         \u_decoder/fir_filter/dp_cluster_0/r180/A2[11] ,
         \u_decoder/fir_filter/dp_cluster_0/r180/A1[7] ,
         \u_decoder/fir_filter/dp_cluster_0/r180/A1[8] ,
         \u_decoder/fir_filter/dp_cluster_0/r180/A1[9] ,
         \u_decoder/fir_filter/dp_cluster_0/r180/A1[10] ,
         \u_decoder/fir_filter/dp_cluster_0/r180/SUMB[2][1] ,
         \u_decoder/fir_filter/dp_cluster_0/r180/SUMB[3][1] ,
         \u_decoder/fir_filter/dp_cluster_0/r180/SUMB[3][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r180/SUMB[4][1] ,
         \u_decoder/fir_filter/dp_cluster_0/r180/SUMB[4][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r180/SUMB[5][1] ,
         \u_decoder/fir_filter/dp_cluster_0/r180/SUMB[5][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r180/SUMB[6][1] ,
         \u_decoder/fir_filter/dp_cluster_0/r180/SUMB[6][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r180/SUMB[7][0] ,
         \u_decoder/fir_filter/dp_cluster_0/r180/SUMB[7][1] ,
         \u_decoder/fir_filter/dp_cluster_0/r180/SUMB[7][2] ,
         \u_decoder/fir_filter/dp_cluster_0/r180/SUMB[7][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r180/SUMB[7][4] ,
         \u_decoder/fir_filter/dp_cluster_0/r180/SUMB[7][5] ,
         \u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[1][0] ,
         \u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[2][0] ,
         \u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[2][1] ,
         \u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[3][0] ,
         \u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[3][1] ,
         \u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[3][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[4][0] ,
         \u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[4][1] ,
         \u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[4][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[5][0] ,
         \u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[5][1] ,
         \u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[5][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[6][0] ,
         \u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[6][1] ,
         \u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[6][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[7][0] ,
         \u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[7][1] ,
         \u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[7][2] ,
         \u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[7][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[7][4] ,
         \u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[7][5] ,
         \u_decoder/fir_filter/dp_cluster_0/r179/A2[6] ,
         \u_decoder/fir_filter/dp_cluster_0/r179/A2[7] ,
         \u_decoder/fir_filter/dp_cluster_0/r179/A2[8] ,
         \u_decoder/fir_filter/dp_cluster_0/r179/A2[9] ,
         \u_decoder/fir_filter/dp_cluster_0/r179/A1[6] ,
         \u_decoder/fir_filter/dp_cluster_0/r179/A1[7] ,
         \u_decoder/fir_filter/dp_cluster_0/r179/A1[8] ,
         \u_decoder/fir_filter/dp_cluster_0/r179/SUMB[1][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r179/SUMB[2][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r179/SUMB[3][1] ,
         \u_decoder/fir_filter/dp_cluster_0/r179/SUMB[3][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r179/SUMB[4][1] ,
         \u_decoder/fir_filter/dp_cluster_0/r179/SUMB[4][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r179/SUMB[5][1] ,
         \u_decoder/fir_filter/dp_cluster_0/r179/SUMB[5][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r179/SUMB[6][1] ,
         \u_decoder/fir_filter/dp_cluster_0/r179/SUMB[6][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r179/SUMB[7][0] ,
         \u_decoder/fir_filter/dp_cluster_0/r179/SUMB[7][1] ,
         \u_decoder/fir_filter/dp_cluster_0/r179/SUMB[7][2] ,
         \u_decoder/fir_filter/dp_cluster_0/r179/SUMB[7][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r179/CARRYB[1][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r179/CARRYB[2][1] ,
         \u_decoder/fir_filter/dp_cluster_0/r179/CARRYB[2][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r179/CARRYB[3][1] ,
         \u_decoder/fir_filter/dp_cluster_0/r179/CARRYB[3][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r179/CARRYB[4][1] ,
         \u_decoder/fir_filter/dp_cluster_0/r179/CARRYB[4][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r179/CARRYB[5][1] ,
         \u_decoder/fir_filter/dp_cluster_0/r179/CARRYB[5][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r179/CARRYB[6][1] ,
         \u_decoder/fir_filter/dp_cluster_0/r179/CARRYB[6][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r179/CARRYB[7][0] ,
         \u_decoder/fir_filter/dp_cluster_0/r179/CARRYB[7][1] ,
         \u_decoder/fir_filter/dp_cluster_0/r179/CARRYB[7][2] ,
         \u_decoder/fir_filter/dp_cluster_0/r179/CARRYB[7][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r178/A2[6] ,
         \u_decoder/fir_filter/dp_cluster_0/r178/A2[7] ,
         \u_decoder/fir_filter/dp_cluster_0/r178/A2[8] ,
         \u_decoder/fir_filter/dp_cluster_0/r178/A2[9] ,
         \u_decoder/fir_filter/dp_cluster_0/r178/A2[10] ,
         \u_decoder/fir_filter/dp_cluster_0/r178/A1[4] ,
         \u_decoder/fir_filter/dp_cluster_0/r178/A1[5] ,
         \u_decoder/fir_filter/dp_cluster_0/r178/A1[6] ,
         \u_decoder/fir_filter/dp_cluster_0/r178/A1[7] ,
         \u_decoder/fir_filter/dp_cluster_0/r178/A1[8] ,
         \u_decoder/fir_filter/dp_cluster_0/r178/A1[9] ,
         \u_decoder/fir_filter/dp_cluster_0/r178/PROD1[5] ,
         \u_decoder/fir_filter/dp_cluster_0/r178/SUMB[2][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r178/SUMB[3][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r178/SUMB[4][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r178/SUMB[5][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r178/SUMB[6][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r178/SUMB[7][0] ,
         \u_decoder/fir_filter/dp_cluster_0/r178/SUMB[7][1] ,
         \u_decoder/fir_filter/dp_cluster_0/r178/SUMB[7][2] ,
         \u_decoder/fir_filter/dp_cluster_0/r178/SUMB[7][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r178/SUMB[7][4] ,
         \u_decoder/fir_filter/dp_cluster_0/r178/CARRYB[2][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r178/CARRYB[3][0] ,
         \u_decoder/fir_filter/dp_cluster_0/r178/CARRYB[3][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r178/CARRYB[4][0] ,
         \u_decoder/fir_filter/dp_cluster_0/r178/CARRYB[4][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r178/CARRYB[5][0] ,
         \u_decoder/fir_filter/dp_cluster_0/r178/CARRYB[5][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r178/CARRYB[6][0] ,
         \u_decoder/fir_filter/dp_cluster_0/r178/CARRYB[6][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r178/CARRYB[7][0] ,
         \u_decoder/fir_filter/dp_cluster_0/r178/CARRYB[7][1] ,
         \u_decoder/fir_filter/dp_cluster_0/r178/CARRYB[7][2] ,
         \u_decoder/fir_filter/dp_cluster_0/r178/CARRYB[7][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r178/CARRYB[7][4] ,
         \u_decoder/fir_filter/dp_cluster_0/r177/A2[6] ,
         \u_decoder/fir_filter/dp_cluster_0/r177/A2[7] ,
         \u_decoder/fir_filter/dp_cluster_0/r177/A2[8] ,
         \u_decoder/fir_filter/dp_cluster_0/r177/A2[9] ,
         \u_decoder/fir_filter/dp_cluster_0/r177/A1[3] ,
         \u_decoder/fir_filter/dp_cluster_0/r177/A1[4] ,
         \u_decoder/fir_filter/dp_cluster_0/r177/A1[5] ,
         \u_decoder/fir_filter/dp_cluster_0/r177/A1[6] ,
         \u_decoder/fir_filter/dp_cluster_0/r177/A1[7] ,
         \u_decoder/fir_filter/dp_cluster_0/r177/A1[8] ,
         \u_decoder/fir_filter/dp_cluster_0/r177/PROD1[4] ,
         \u_decoder/fir_filter/dp_cluster_0/r177/SUMB[2][2] ,
         \u_decoder/fir_filter/dp_cluster_0/r177/SUMB[3][2] ,
         \u_decoder/fir_filter/dp_cluster_0/r177/SUMB[4][2] ,
         \u_decoder/fir_filter/dp_cluster_0/r177/SUMB[5][2] ,
         \u_decoder/fir_filter/dp_cluster_0/r177/SUMB[6][2] ,
         \u_decoder/fir_filter/dp_cluster_0/r177/SUMB[7][0] ,
         \u_decoder/fir_filter/dp_cluster_0/r177/SUMB[7][1] ,
         \u_decoder/fir_filter/dp_cluster_0/r177/SUMB[7][2] ,
         \u_decoder/fir_filter/dp_cluster_0/r177/SUMB[7][3] ,
         \u_decoder/fir_filter/dp_cluster_0/r177/CARRYB[2][0] ,
         \u_decoder/fir_filter/dp_cluster_0/r177/CARRYB[2][2] ,
         \u_decoder/fir_filter/dp_cluster_0/r177/CARRYB[3][0] ,
         \u_decoder/fir_filter/dp_cluster_0/r177/CARRYB[3][2] ,
         \u_decoder/fir_filter/dp_cluster_0/r177/CARRYB[4][0] ,
         \u_decoder/fir_filter/dp_cluster_0/r177/CARRYB[4][2] ,
         \u_decoder/fir_filter/dp_cluster_0/r177/CARRYB[5][0] ,
         \u_decoder/fir_filter/dp_cluster_0/r177/CARRYB[5][2] ,
         \u_decoder/fir_filter/dp_cluster_0/r177/CARRYB[6][0] ,
         \u_decoder/fir_filter/dp_cluster_0/r177/CARRYB[6][2] ,
         \u_decoder/fir_filter/dp_cluster_0/r177/CARRYB[7][0] ,
         \u_decoder/fir_filter/dp_cluster_0/r177/CARRYB[7][1] ,
         \u_decoder/fir_filter/dp_cluster_0/r177/CARRYB[7][2] ,
         \u_decoder/fir_filter/dp_cluster_0/r177/CARRYB[7][3] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_151/A2[2] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_151/A2[3] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_151/A2[4] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_151/A2[5] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_151/A1[2] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_151/A1[3] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_151/A1[4] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_151/SUMB[1][1] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_151/SUMB[1][2] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_151/SUMB[2][1] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_151/SUMB[2][2] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_151/SUMB[3][0] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_151/SUMB[3][1] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_151/SUMB[3][2] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_151/SUMB[3][3] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_151/CARRYB[1][0] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_151/CARRYB[1][1] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_151/CARRYB[1][2] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_151/CARRYB[2][0] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_151/CARRYB[2][1] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_151/CARRYB[2][2] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_151/CARRYB[3][0] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_151/CARRYB[3][1] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_151/CARRYB[3][2] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_151/CARRYB[3][3] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_151/ab[0][1] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_151/ab[0][2] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_151/ab[0][3] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_151/ab[1][0] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_151/ab[1][1] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_151/ab[1][2] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_151/ab[1][3] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_151/ab[2][0] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_151/ab[2][1] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_151/ab[2][2] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_151/ab[2][3] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_151/ab[3][0] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_151/ab[3][1] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_151/ab[3][2] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_151/ab[3][3] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_148/A2[2] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_148/A2[3] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_148/A2[4] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_148/A2[5] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_148/A1[2] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_148/A1[3] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_148/A1[4] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_148/SUMB[1][1] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_148/SUMB[1][2] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_148/SUMB[2][1] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_148/SUMB[2][2] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_148/SUMB[3][0] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_148/SUMB[3][1] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_148/SUMB[3][2] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_148/SUMB[3][3] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_148/CARRYB[1][0] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_148/CARRYB[1][1] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_148/CARRYB[1][2] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_148/CARRYB[2][0] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_148/CARRYB[2][1] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_148/CARRYB[2][2] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_148/CARRYB[3][0] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_148/CARRYB[3][1] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_148/CARRYB[3][2] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_148/CARRYB[3][3] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_148/ab[0][1] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_148/ab[0][2] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_148/ab[0][3] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_148/ab[1][0] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_148/ab[1][1] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_148/ab[1][2] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_148/ab[1][3] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_148/ab[2][0] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_148/ab[2][1] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_148/ab[2][2] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_148/ab[2][3] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_148/ab[3][0] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_148/ab[3][1] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_148/ab[3][2] ,
         \u_decoder/iq_demod/dp_cluster_0/mult_148/ab[3][3] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_150/A2[2] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_150/A2[3] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_150/A2[4] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_150/A2[5] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_150/A1[2] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_150/A1[3] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_150/A1[4] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_150/SUMB[1][1] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_150/SUMB[1][2] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_150/SUMB[2][1] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_150/SUMB[2][2] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_150/SUMB[3][0] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_150/SUMB[3][1] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_150/SUMB[3][2] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_150/SUMB[3][3] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_150/CARRYB[1][0] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_150/CARRYB[1][1] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_150/CARRYB[1][2] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_150/CARRYB[2][0] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_150/CARRYB[2][1] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_150/CARRYB[2][2] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_150/CARRYB[3][0] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_150/CARRYB[3][1] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_150/CARRYB[3][2] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_150/CARRYB[3][3] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_150/ab[0][1] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_150/ab[0][2] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_150/ab[0][3] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_150/ab[1][0] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_150/ab[1][1] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_150/ab[1][2] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_150/ab[1][3] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_150/ab[2][0] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_150/ab[2][1] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_150/ab[2][2] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_150/ab[2][3] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_150/ab[3][0] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_150/ab[3][1] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_150/ab[3][2] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_150/ab[3][3] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_149/A2[2] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_149/A2[3] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_149/A2[4] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_149/A2[5] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_149/A1[2] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_149/A1[3] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_149/A1[4] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_149/SUMB[1][1] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_149/SUMB[1][2] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_149/SUMB[2][1] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_149/SUMB[2][2] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_149/SUMB[3][0] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_149/SUMB[3][1] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_149/SUMB[3][2] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_149/SUMB[3][3] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_149/CARRYB[1][0] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_149/CARRYB[1][1] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_149/CARRYB[1][2] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_149/CARRYB[2][0] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_149/CARRYB[2][1] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_149/CARRYB[2][2] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_149/CARRYB[3][0] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_149/CARRYB[3][1] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_149/CARRYB[3][2] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_149/CARRYB[3][3] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_149/ab[0][1] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_149/ab[0][2] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_149/ab[0][3] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_149/ab[1][0] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_149/ab[1][1] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_149/ab[1][2] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_149/ab[1][3] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_149/ab[2][0] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_149/ab[2][1] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_149/ab[2][2] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_149/ab[2][3] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_149/ab[3][0] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_149/ab[3][1] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_149/ab[3][2] ,
         \u_decoder/iq_demod/dp_cluster_1/mult_149/ab[3][3] ,
         \u_cdr/dp_cluster_0/mult_add_59_aco/PROD_not[0] ,
         \u_cdr/dp_cluster_0/mult_add_59_aco/PROD_not[1] ,
         \u_cdr/dp_cluster_0/mult_add_59_aco/PROD_not[2] ,
         \u_cdr/dp_cluster_0/mult_add_59_aco/PROD_not[3] , n1, n2, n3, n4, n5,
         n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
         n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
         n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
         n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
         n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
         n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
         n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
         n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
         n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
         n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
         n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
         n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
         n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
         n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
         n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
         n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
         n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
         n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
         n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
         n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
         n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
         n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
         n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
         n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
         n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
         n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404,
         n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414,
         n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424,
         n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434,
         n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444,
         n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454,
         n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464,
         n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474,
         n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484,
         n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494,
         n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504,
         n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514,
         n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524,
         n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534,
         n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544,
         n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554,
         n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564,
         n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574,
         n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584,
         n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594,
         n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604,
         n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614,
         n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624,
         n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634,
         n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644,
         n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654,
         n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664,
         n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674,
         n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684,
         n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694,
         n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704,
         n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714,
         n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724,
         n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734,
         n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744,
         n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754,
         n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764,
         n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774,
         n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784,
         n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794,
         n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804,
         n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814,
         n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824,
         n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834,
         n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844,
         n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854,
         n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864,
         n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874,
         n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884,
         n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894,
         n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904,
         n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914,
         n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924,
         n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934,
         n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944,
         n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954,
         n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964,
         n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974,
         n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984,
         n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994,
         n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004,
         n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014,
         n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024,
         n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034,
         n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044,
         n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054,
         n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064,
         n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074,
         n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084,
         n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094,
         n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104,
         n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114,
         n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124,
         n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134,
         n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144,
         n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154,
         n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164,
         n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174,
         n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184,
         n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194,
         n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204,
         n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214,
         n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224,
         n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234,
         n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244,
         n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254,
         n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264,
         n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274,
         n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284,
         n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294,
         n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304,
         n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314,
         n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324,
         n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334,
         n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344,
         n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354,
         n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364,
         n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374,
         n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384,
         n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394,
         n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404,
         n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414,
         n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424,
         n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434,
         n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444,
         n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454,
         n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464,
         n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474,
         n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484,
         n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494,
         n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504,
         n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514,
         n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524,
         n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534,
         n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544,
         n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554,
         n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564,
         n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574,
         n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584,
         n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594,
         n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604,
         n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614,
         n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624,
         n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634,
         n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644,
         n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654,
         n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664,
         n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674,
         n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684,
         n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694,
         n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704,
         n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714,
         n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724,
         n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734,
         n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744,
         n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754,
         n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764,
         n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774,
         n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784,
         n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794,
         n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804,
         n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814,
         n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824,
         n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834,
         n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844,
         n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854,
         n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864,
         n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874,
         n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884,
         n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894,
         n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904,
         n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914,
         n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924,
         n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934,
         n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944,
         n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954,
         n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964,
         n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974,
         n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984,
         n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994,
         n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004,
         n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014,
         n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024,
         n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034,
         n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044,
         n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054,
         n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064,
         n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074,
         n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084,
         n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094,
         n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104,
         n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114,
         n3115, n3116, n3117, n3118;
  wire   [3:0] sig_coder_outSinI;
  wire   [3:0] sig_coder_outSinQ;
  wire   [3:0] sig_coder_outSinIMasked;
  wire   [3:0] sig_coder_outSinQMasked;
  wire   [3:0] sig_decod_outI;
  wire   [3:0] sig_decod_outQ;
  wire   [3:0] sig_outFIFO_outData;
  wire   [7:0] sig_DEMUX_outDEMUX1;
  wire   [7:0] sig_DEMUX_outDEMUX2;
  wire   [7:0] sig_DEMUX_outDEMUX17;
  wire   [7:0] sig_DEMUX_outDEMUX18;
  wire   [3:0] sig_MUX_outMUX6;
  wire   [3:0] sig_MUX_outMUX7;
  wire   [6:0] \u_inFIFO/j_FIFO ;
  wire   [3:0] \u_inFIFO/currentState ;
  wire   [19:0] \u_coder/j ;
  wire   [19:0] \u_coder/i ;
  wire   [19:0] \u_coder/c ;
  wire   [7:0] \u_decoder/Q_prefilter ;
  wire   [7:0] \u_decoder/I_prefilter ;
  wire   [2:0] \u_cordic/present_state ;
  wire   [3:0] \u_cordic/Q ;
  wire   [3:0] \u_cordic/I ;
  wire   [15:0] \u_cordic/cordic_to_rotation ;
  wire   [5:0] \u_cdr/w_nb_P ;
  wire   [2:0] \u_cdr/cnt ;
  wire   [1:0] \u_cdr/cnt_d ;
  wire   [3:0] \u_cdr/cnt_in ;
  wire   [1:0] \u_outFIFO/k_FIFO ;
  wire   [6:0] \u_outFIFO/i_FIFO ;
  wire   [3:0] \u_outFIFO/currentState ;
  wire   [7:0] \u_decoder/iq_demod/dp_cluster_1/mult_I_sin_out ;
  wire   [7:0] \u_decoder/iq_demod/dp_cluster_1/mult_Q_cos_out ;
  wire   [7:0] \u_decoder/iq_demod/dp_cluster_0/mult_I_cos_out ;
  wire   [7:0] \u_decoder/iq_demod/dp_cluster_0/mult_Q_sin_out ;
  wire   [3:0] \u_decoder/iq_demod/Q_if_signed ;
  wire   [3:0] \u_decoder/iq_demod/I_if_signed ;
  wire   [7:0] \u_decoder/iq_demod/add_Q_out ;
  wire   [7:0] \u_decoder/iq_demod/add_I_out ;
  wire   [1:0] \u_decoder/iq_demod/state ;
  wire   [3:0] \u_decoder/iq_demod/sin_out ;
  wire   [3:0] \u_decoder/iq_demod/cos_out ;
  wire   [20:0] \u_decoder/fir_filter/Q_data_mult_8_buff ;
  wire   [15:0] \u_decoder/fir_filter/Q_data_mult_7_buff ;
  wire   [15:0] \u_decoder/fir_filter/Q_data_mult_6_buff ;
  wire   [15:0] \u_decoder/fir_filter/Q_data_mult_5_buff ;
  wire   [15:0] \u_decoder/fir_filter/Q_data_mult_4 ;
  wire   [15:0] \u_decoder/fir_filter/Q_data_mult_4_buff ;
  wire   [15:0] \u_decoder/fir_filter/Q_data_mult_3 ;
  wire   [15:0] \u_decoder/fir_filter/Q_data_mult_3_buff ;
  wire   [15:0] \u_decoder/fir_filter/Q_data_mult_2_buff ;
  wire   [15:0] \u_decoder/fir_filter/Q_data_mult_1_buff ;
  wire   [11:0] \u_decoder/fir_filter/Q_data_mult_0 ;
  wire   [14:0] \u_decoder/fir_filter/Q_data_mult_0_buff ;
  wire   [20:0] \u_decoder/fir_filter/Q_data_add_7 ;
  wire   [20:0] \u_decoder/fir_filter/Q_data_add_7_buff ;
  wire   [20:0] \u_decoder/fir_filter/Q_data_add_6 ;
  wire   [20:0] \u_decoder/fir_filter/Q_data_add_6_buff ;
  wire   [20:0] \u_decoder/fir_filter/Q_data_add_5 ;
  wire   [20:0] \u_decoder/fir_filter/Q_data_add_5_buff ;
  wire   [20:0] \u_decoder/fir_filter/Q_data_add_4 ;
  wire   [20:0] \u_decoder/fir_filter/Q_data_add_4_buff ;
  wire   [20:0] \u_decoder/fir_filter/Q_data_add_3 ;
  wire   [20:0] \u_decoder/fir_filter/Q_data_add_3_buff ;
  wire   [20:0] \u_decoder/fir_filter/Q_data_add_2 ;
  wire   [20:0] \u_decoder/fir_filter/Q_data_add_2_buff ;
  wire   [14:0] \u_decoder/fir_filter/Q_data_add_1 ;
  wire   [14:0] \u_decoder/fir_filter/Q_data_add_1_buff ;
  wire   [20:0] \u_decoder/fir_filter/I_data_mult_8_buff ;
  wire   [15:0] \u_decoder/fir_filter/I_data_mult_7_buff ;
  wire   [15:0] \u_decoder/fir_filter/I_data_mult_6_buff ;
  wire   [15:0] \u_decoder/fir_filter/I_data_mult_5_buff ;
  wire   [15:0] \u_decoder/fir_filter/I_data_mult_4 ;
  wire   [15:0] \u_decoder/fir_filter/I_data_mult_4_buff ;
  wire   [15:0] \u_decoder/fir_filter/I_data_mult_3 ;
  wire   [15:0] \u_decoder/fir_filter/I_data_mult_3_buff ;
  wire   [15:0] \u_decoder/fir_filter/I_data_mult_2_buff ;
  wire   [15:0] \u_decoder/fir_filter/I_data_mult_1_buff ;
  wire   [11:0] \u_decoder/fir_filter/I_data_mult_0 ;
  wire   [14:0] \u_decoder/fir_filter/I_data_mult_0_buff ;
  wire   [20:0] \u_decoder/fir_filter/I_data_add_7 ;
  wire   [20:0] \u_decoder/fir_filter/I_data_add_7_buff ;
  wire   [20:0] \u_decoder/fir_filter/I_data_add_6 ;
  wire   [20:0] \u_decoder/fir_filter/I_data_add_6_buff ;
  wire   [20:0] \u_decoder/fir_filter/I_data_add_5 ;
  wire   [20:0] \u_decoder/fir_filter/I_data_add_5_buff ;
  wire   [20:0] \u_decoder/fir_filter/I_data_add_4 ;
  wire   [20:0] \u_decoder/fir_filter/I_data_add_4_buff ;
  wire   [20:0] \u_decoder/fir_filter/I_data_add_3 ;
  wire   [20:0] \u_decoder/fir_filter/I_data_add_3_buff ;
  wire   [20:0] \u_decoder/fir_filter/I_data_add_2 ;
  wire   [20:0] \u_decoder/fir_filter/I_data_add_2_buff ;
  wire   [14:0] \u_decoder/fir_filter/I_data_add_1 ;
  wire   [14:0] \u_decoder/fir_filter/I_data_add_1_buff ;
  wire   [14:11] \u_decoder/fir_filter/Q_data_add_0 ;
  wire   [14:11] \u_decoder/fir_filter/I_data_add_0 ;
  wire   [1:0] \u_decoder/fir_filter/state ;
  wire   [15:0] \u_cordic/my_rotation/delta ;
  wire   [5:0] \u_cdr/dec1/cnt_r ;
  wire   [2:0] \u_decoder/iq_demod/cossin_dig/val_counter ;
  wire   [2:0] \u_decoder/iq_demod/cossin_dig/counter ;
  wire   [5:0] \u_cdr/div1/cnt_div/cnt ;
  wire   [5:0] \u_cdr/dec1/cnt_dec/cnt_dec ;
  wire   [5:0] \u_cdr/phd1/cnt_phd/cnt ;
  wire   [5:2] \u_cdr/phd1/cnt_phd/add_58/carry ;
  wire   [5:2] \u_cdr/dec1/cnt_dec/add_20/carry ;
  wire   [5:2] \u_cdr/div1/cnt_div/add_58/carry ;
  wire   [5:2] \u_cdr/dec1/add_40/carry ;
  wire   [16:0] \u_cordic/my_rotation/sub_35/carry ;
  wire   [15:1] \u_cordic/my_rotation/add_38/carry ;
  wire   [7:1] \u_cordic/mycordic/r144/carry ;
  wire   [15:1] \u_cordic/mycordic/r173/carry ;
  wire   [8:0] \u_cordic/mycordic/sub_178/carry ;
  wire   [8:0] \u_cordic/mycordic/sub_182/carry ;
  wire   [7:1] \u_cordic/mycordic/add_189/carry ;
  wire   [8:0] \u_cordic/mycordic/sub_190/carry ;
  wire   [8:0] \u_cordic/mycordic/sub_194/carry ;
  wire   [7:1] \u_cordic/mycordic/add_195/carry ;
  wire   [7:1] \u_cordic/mycordic/add_200/carry ;
  wire   [8:0] \u_cordic/mycordic/sub_201/carry ;
  wire   [15:1] \u_cordic/mycordic/add_202/carry ;
  wire   [8:0] \u_cordic/mycordic/sub_205/carry ;
  wire   [7:1] \u_cordic/mycordic/add_206/carry ;
  wire   [16:0] \u_cordic/mycordic/sub_207/carry ;
  wire   [7:1] \u_cordic/mycordic/add_211/carry ;
  wire   [8:0] \u_cordic/mycordic/sub_212/carry ;
  wire   [8:0] \u_cordic/mycordic/sub_216/carry ;
  wire   [7:1] \u_cordic/mycordic/add_217/carry ;
  wire   [15:1] \u_cordic/mycordic/add_233/carry ;
  wire   [16:0] \u_cordic/mycordic/sub_236/carry ;
  wire   [15:1] \u_cordic/mycordic/add_262/carry ;
  wire   [8:0] \u_cordic/mycordic/sub_add_150_b0/carry ;
  wire   [8:0] \u_cordic/mycordic/sub_add_151_b0/carry ;
  wire   [14:1] \u_decoder/fir_filter/add_294/carry ;
  wire   [20:1] \u_decoder/fir_filter/add_295/carry ;
  wire   [20:1] \u_decoder/fir_filter/add_296/carry ;
  wire   [20:1] \u_decoder/fir_filter/add_297/carry ;
  wire   [20:1] \u_decoder/fir_filter/add_298/carry ;
  wire   [20:1] \u_decoder/fir_filter/add_299/carry ;
  wire   [20:1] \u_decoder/fir_filter/add_300/carry ;
  wire   [20:1] \u_decoder/fir_filter/add_301/carry ;
  wire   [14:1] \u_decoder/fir_filter/add_326/carry ;
  wire   [20:1] \u_decoder/fir_filter/add_327/carry ;
  wire   [20:1] \u_decoder/fir_filter/add_328/carry ;
  wire   [20:1] \u_decoder/fir_filter/add_329/carry ;
  wire   [20:1] \u_decoder/fir_filter/add_330/carry ;
  wire   [20:1] \u_decoder/fir_filter/add_331/carry ;
  wire   [20:1] \u_decoder/fir_filter/add_332/carry ;
  wire   [20:1] \u_decoder/fir_filter/add_333/carry ;
  wire   [8:0] \u_decoder/iq_demod/dp_cluster_0/sub_153/carry ;
  wire   [7:1] \u_decoder/iq_demod/dp_cluster_1/add_154/carry ;
  wire   [8:0] \u_outFIFO/r98/carry ;
  wire   [7:2] \u_outFIFO/add_255/carry ;
  wire   [6:2] \u_outFIFO/add_256/carry ;
  wire   [6:2] \u_outFIFO/add_260/carry ;
  wire   [6:2] \u_outFIFO/add_360/carry ;
  wire   [19:2] \u_coder/add_93/carry ;
  wire   [19:2] \u_coder/add_206/carry ;
  wire   [19:2] \u_coder/add_282/carry ;
  wire   [8:0] \u_inFIFO/r96/carry ;
  wire   [6:2] \u_inFIFO/add_252/carry ;
  wire   [6:2] \u_inFIFO/add_253/carry ;
  wire   [7:2] \u_inFIFO/add_263/carry ;
  wire   [6:2] \u_inFIFO/add_357/carry ;

  OAI222 \u_inFIFO/U505  ( .A(n1237), .B(\u_inFIFO/n531 ), .C(
        \u_inFIFO/currentState [0]), .D(\u_inFIFO/n551 ), .Q(\u_inFIFO/n566 )
         );
  OAI212 \u_inFIFO/U504  ( .A(\u_inFIFO/n565 ), .B(n1241), .C(n1829), .Q(
        \u_inFIFO/N48 ) );
  OAI212 \u_inFIFO/U501  ( .A(\u_inFIFO/n562 ), .B(n1236), .C(n1829), .Q(
        \u_inFIFO/N49 ) );
  OAI212 \u_inFIFO/U484  ( .A(n1828), .B(\u_inFIFO/n179 ), .C(\u_inFIFO/n548 ), 
        .Q(\u_inFIFO/n582 ) );
  OAI212 \u_inFIFO/U476  ( .A(n1828), .B(\u_inFIFO/n188 ), .C(\u_inFIFO/n540 ), 
        .Q(\u_inFIFO/n581 ) );
  OAI212 \u_inFIFO/U474  ( .A(n1828), .B(\u_inFIFO/n182 ), .C(\u_inFIFO/n539 ), 
        .Q(\u_inFIFO/n580 ) );
  OAI212 \u_inFIFO/U472  ( .A(n1828), .B(\u_inFIFO/n183 ), .C(\u_inFIFO/n538 ), 
        .Q(\u_inFIFO/n579 ) );
  OAI212 \u_inFIFO/U470  ( .A(n1828), .B(\u_inFIFO/n184 ), .C(\u_inFIFO/n537 ), 
        .Q(\u_inFIFO/n578 ) );
  OAI212 \u_inFIFO/U468  ( .A(n1828), .B(\u_inFIFO/n185 ), .C(\u_inFIFO/n536 ), 
        .Q(\u_inFIFO/n577 ) );
  OAI212 \u_inFIFO/U466  ( .A(n1828), .B(\u_inFIFO/n186 ), .C(\u_inFIFO/n535 ), 
        .Q(\u_inFIFO/n576 ) );
  OAI212 \u_inFIFO/U464  ( .A(n1828), .B(\u_inFIFO/n187 ), .C(\u_inFIFO/n532 ), 
        .Q(\u_inFIFO/n575 ) );
  OAI222 \u_inFIFO/U461  ( .A(\u_inFIFO/n217 ), .B(\u_inFIFO/n198 ), .C(
        \u_inFIFO/N44 ), .D(\u_inFIFO/n216 ), .Q(\u_inFIFO/n574 ) );
  OAI222 \u_inFIFO/U459  ( .A(\u_inFIFO/n217 ), .B(\u_inFIFO/n197 ), .C(
        \u_inFIFO/n530 ), .D(\u_inFIFO/n216 ), .Q(\u_inFIFO/n573 ) );
  OAI212 \u_inFIFO/U434  ( .A(\u_inFIFO/n511 ), .B(n1203), .C(n1209), .Q(
        \u_inFIFO/n510 ) );
  OAI212 \u_inFIFO/U427  ( .A(\u_inFIFO/n509 ), .B(n1203), .C(n1209), .Q(
        \u_inFIFO/n508 ) );
  OAI212 \u_inFIFO/U423  ( .A(\u_inFIFO/n507 ), .B(n1203), .C(n1209), .Q(
        \u_inFIFO/n506 ) );
  OAI212 \u_inFIFO/U419  ( .A(\u_inFIFO/n504 ), .B(n1203), .C(n1209), .Q(
        \u_inFIFO/n503 ) );
  OAI212 \u_inFIFO/U415  ( .A(\u_inFIFO/n502 ), .B(n1203), .C(n1209), .Q(
        \u_inFIFO/n501 ) );
  OAI212 \u_inFIFO/U412  ( .A(\u_inFIFO/n500 ), .B(n1203), .C(n1209), .Q(
        \u_inFIFO/n499 ) );
  OAI212 \u_inFIFO/U409  ( .A(\u_inFIFO/n498 ), .B(n1203), .C(n1209), .Q(
        \u_inFIFO/n497 ) );
  OAI212 \u_inFIFO/U406  ( .A(\u_inFIFO/n495 ), .B(n1203), .C(n1209), .Q(
        \u_inFIFO/n494 ) );
  OAI212 \u_inFIFO/U402  ( .A(\u_inFIFO/n493 ), .B(n1203), .C(n1209), .Q(
        \u_inFIFO/n492 ) );
  OAI212 \u_inFIFO/U399  ( .A(\u_inFIFO/n491 ), .B(n1203), .C(n1209), .Q(
        \u_inFIFO/n490 ) );
  OAI212 \u_inFIFO/U396  ( .A(\u_inFIFO/n489 ), .B(n1203), .C(n1209), .Q(
        \u_inFIFO/n488 ) );
  OAI212 \u_inFIFO/U393  ( .A(\u_inFIFO/n486 ), .B(n1203), .C(n1209), .Q(
        \u_inFIFO/n485 ) );
  OAI212 \u_inFIFO/U389  ( .A(\u_inFIFO/n483 ), .B(n1203), .C(n1209), .Q(
        \u_inFIFO/n482 ) );
  OAI212 \u_inFIFO/U386  ( .A(\u_inFIFO/n480 ), .B(n1203), .C(n1209), .Q(
        \u_inFIFO/n479 ) );
  OAI212 \u_inFIFO/U383  ( .A(\u_inFIFO/n477 ), .B(n1203), .C(n1209), .Q(
        \u_inFIFO/n476 ) );
  OAI212 \u_inFIFO/U380  ( .A(\u_inFIFO/n472 ), .B(n1203), .C(n1209), .Q(
        \u_inFIFO/n471 ) );
  OAI212 \u_inFIFO/U377  ( .A(\u_inFIFO/n470 ), .B(n1203), .C(n1209), .Q(
        \u_inFIFO/n469 ) );
  OAI212 \u_inFIFO/U375  ( .A(\u_inFIFO/n468 ), .B(n1206), .C(n1209), .Q(
        \u_inFIFO/n467 ) );
  OAI212 \u_inFIFO/U373  ( .A(\u_inFIFO/n466 ), .B(n1205), .C(n1209), .Q(
        \u_inFIFO/n465 ) );
  OAI212 \u_inFIFO/U371  ( .A(\u_inFIFO/n464 ), .B(n1204), .C(n1209), .Q(
        \u_inFIFO/n463 ) );
  OAI212 \u_inFIFO/U369  ( .A(\u_inFIFO/n462 ), .B(n1208), .C(n1209), .Q(
        \u_inFIFO/n461 ) );
  OAI212 \u_inFIFO/U367  ( .A(\u_inFIFO/n460 ), .B(n1208), .C(n1209), .Q(
        \u_inFIFO/n459 ) );
  OAI212 \u_inFIFO/U365  ( .A(\u_inFIFO/n458 ), .B(n1208), .C(n1209), .Q(
        \u_inFIFO/n457 ) );
  OAI212 \u_inFIFO/U363  ( .A(\u_inFIFO/n456 ), .B(n1208), .C(n1209), .Q(
        \u_inFIFO/n455 ) );
  OAI212 \u_inFIFO/U361  ( .A(\u_inFIFO/n454 ), .B(n1208), .C(n1210), .Q(
        \u_inFIFO/n453 ) );
  OAI212 \u_inFIFO/U359  ( .A(\u_inFIFO/n452 ), .B(n1208), .C(\u_inFIFO/n225 ), 
        .Q(\u_inFIFO/n451 ) );
  OAI212 \u_inFIFO/U357  ( .A(\u_inFIFO/n450 ), .B(n1208), .C(n1210), .Q(
        \u_inFIFO/n449 ) );
  OAI212 \u_inFIFO/U355  ( .A(\u_inFIFO/n448 ), .B(n1208), .C(n1210), .Q(
        \u_inFIFO/n447 ) );
  OAI212 \u_inFIFO/U353  ( .A(\u_inFIFO/n446 ), .B(n1208), .C(\u_inFIFO/n225 ), 
        .Q(\u_inFIFO/n445 ) );
  OAI212 \u_inFIFO/U351  ( .A(\u_inFIFO/n444 ), .B(n1208), .C(\u_inFIFO/n225 ), 
        .Q(\u_inFIFO/n443 ) );
  OAI212 \u_inFIFO/U349  ( .A(\u_inFIFO/n442 ), .B(n1208), .C(n1210), .Q(
        \u_inFIFO/n441 ) );
  OAI212 \u_inFIFO/U347  ( .A(\u_inFIFO/n439 ), .B(n1208), .C(\u_inFIFO/n225 ), 
        .Q(\u_inFIFO/n438 ) );
  OAI212 \u_inFIFO/U344  ( .A(\u_inFIFO/n437 ), .B(n1208), .C(n1210), .Q(
        \u_inFIFO/n436 ) );
  OAI212 \u_inFIFO/U342  ( .A(\u_inFIFO/n435 ), .B(n1208), .C(n1210), .Q(
        \u_inFIFO/n434 ) );
  OAI212 \u_inFIFO/U340  ( .A(\u_inFIFO/n433 ), .B(n1208), .C(\u_inFIFO/n225 ), 
        .Q(\u_inFIFO/n432 ) );
  OAI212 \u_inFIFO/U338  ( .A(\u_inFIFO/n431 ), .B(n1204), .C(\u_inFIFO/n225 ), 
        .Q(\u_inFIFO/n430 ) );
  OAI212 \u_inFIFO/U336  ( .A(\u_inFIFO/n429 ), .B(n1204), .C(n1210), .Q(
        \u_inFIFO/n428 ) );
  OAI212 \u_inFIFO/U334  ( .A(\u_inFIFO/n427 ), .B(n1204), .C(\u_inFIFO/n225 ), 
        .Q(\u_inFIFO/n426 ) );
  OAI212 \u_inFIFO/U332  ( .A(\u_inFIFO/n425 ), .B(n1204), .C(n1210), .Q(
        \u_inFIFO/n424 ) );
  OAI212 \u_inFIFO/U330  ( .A(\u_inFIFO/n423 ), .B(n1204), .C(n1210), .Q(
        \u_inFIFO/n422 ) );
  OAI212 \u_inFIFO/U328  ( .A(\u_inFIFO/n421 ), .B(n1204), .C(\u_inFIFO/n225 ), 
        .Q(\u_inFIFO/n420 ) );
  OAI212 \u_inFIFO/U326  ( .A(\u_inFIFO/n419 ), .B(n1204), .C(\u_inFIFO/n225 ), 
        .Q(\u_inFIFO/n418 ) );
  OAI212 \u_inFIFO/U324  ( .A(\u_inFIFO/n417 ), .B(n1204), .C(n1210), .Q(
        \u_inFIFO/n416 ) );
  OAI212 \u_inFIFO/U322  ( .A(\u_inFIFO/n415 ), .B(n1204), .C(\u_inFIFO/n225 ), 
        .Q(\u_inFIFO/n414 ) );
  OAI212 \u_inFIFO/U320  ( .A(\u_inFIFO/n413 ), .B(n1204), .C(n1210), .Q(
        \u_inFIFO/n412 ) );
  OAI212 \u_inFIFO/U318  ( .A(\u_inFIFO/n411 ), .B(n1204), .C(n1210), .Q(
        \u_inFIFO/n410 ) );
  OAI212 \u_inFIFO/U316  ( .A(\u_inFIFO/n409 ), .B(n1204), .C(\u_inFIFO/n225 ), 
        .Q(\u_inFIFO/n408 ) );
  OAI212 \u_inFIFO/U314  ( .A(\u_inFIFO/n406 ), .B(n1204), .C(n1209), .Q(
        \u_inFIFO/n405 ) );
  OAI212 \u_inFIFO/U311  ( .A(\u_inFIFO/n404 ), .B(n1204), .C(n1210), .Q(
        \u_inFIFO/n403 ) );
  OAI212 \u_inFIFO/U309  ( .A(\u_inFIFO/n402 ), .B(n1204), .C(\u_inFIFO/n225 ), 
        .Q(\u_inFIFO/n401 ) );
  OAI212 \u_inFIFO/U307  ( .A(\u_inFIFO/n400 ), .B(n1204), .C(n1210), .Q(
        \u_inFIFO/n399 ) );
  OAI212 \u_inFIFO/U305  ( .A(\u_inFIFO/n398 ), .B(n1204), .C(n1209), .Q(
        \u_inFIFO/n397 ) );
  OAI212 \u_inFIFO/U303  ( .A(\u_inFIFO/n396 ), .B(n1204), .C(n1209), .Q(
        \u_inFIFO/n395 ) );
  OAI212 \u_inFIFO/U301  ( .A(\u_inFIFO/n394 ), .B(n1205), .C(n1209), .Q(
        \u_inFIFO/n393 ) );
  OAI212 \u_inFIFO/U299  ( .A(\u_inFIFO/n392 ), .B(n1205), .C(n1209), .Q(
        \u_inFIFO/n391 ) );
  OAI212 \u_inFIFO/U297  ( .A(\u_inFIFO/n390 ), .B(n1205), .C(n1209), .Q(
        \u_inFIFO/n389 ) );
  OAI212 \u_inFIFO/U295  ( .A(\u_inFIFO/n388 ), .B(n1205), .C(n1209), .Q(
        \u_inFIFO/n387 ) );
  OAI212 \u_inFIFO/U293  ( .A(\u_inFIFO/n386 ), .B(n1205), .C(n1209), .Q(
        \u_inFIFO/n385 ) );
  OAI212 \u_inFIFO/U291  ( .A(\u_inFIFO/n384 ), .B(n1205), .C(n1209), .Q(
        \u_inFIFO/n383 ) );
  OAI212 \u_inFIFO/U289  ( .A(\u_inFIFO/n382 ), .B(n1205), .C(n1209), .Q(
        \u_inFIFO/n381 ) );
  OAI212 \u_inFIFO/U287  ( .A(\u_inFIFO/n380 ), .B(n1205), .C(n1209), .Q(
        \u_inFIFO/n379 ) );
  OAI212 \u_inFIFO/U285  ( .A(\u_inFIFO/n378 ), .B(n1205), .C(n1209), .Q(
        \u_inFIFO/n377 ) );
  OAI212 \u_inFIFO/U283  ( .A(\u_inFIFO/n376 ), .B(n1205), .C(n1209), .Q(
        \u_inFIFO/n375 ) );
  OAI212 \u_inFIFO/U281  ( .A(\u_inFIFO/n373 ), .B(n1205), .C(n1209), .Q(
        \u_inFIFO/n372 ) );
  OAI212 \u_inFIFO/U278  ( .A(\u_inFIFO/n371 ), .B(n1205), .C(n1209), .Q(
        \u_inFIFO/n370 ) );
  OAI212 \u_inFIFO/U276  ( .A(\u_inFIFO/n369 ), .B(n1205), .C(n1209), .Q(
        \u_inFIFO/n368 ) );
  OAI212 \u_inFIFO/U274  ( .A(\u_inFIFO/n367 ), .B(n1205), .C(n1209), .Q(
        \u_inFIFO/n366 ) );
  OAI212 \u_inFIFO/U272  ( .A(\u_inFIFO/n365 ), .B(n1205), .C(n1209), .Q(
        \u_inFIFO/n364 ) );
  OAI212 \u_inFIFO/U270  ( .A(\u_inFIFO/n363 ), .B(n1205), .C(n1209), .Q(
        \u_inFIFO/n362 ) );
  OAI212 \u_inFIFO/U268  ( .A(\u_inFIFO/n361 ), .B(n1205), .C(n1209), .Q(
        \u_inFIFO/n360 ) );
  OAI212 \u_inFIFO/U266  ( .A(\u_inFIFO/n359 ), .B(n1205), .C(n1209), .Q(
        \u_inFIFO/n358 ) );
  OAI212 \u_inFIFO/U264  ( .A(\u_inFIFO/n357 ), .B(n1206), .C(n1209), .Q(
        \u_inFIFO/n356 ) );
  OAI212 \u_inFIFO/U262  ( .A(\u_inFIFO/n355 ), .B(n1206), .C(n1209), .Q(
        \u_inFIFO/n354 ) );
  OAI212 \u_inFIFO/U260  ( .A(\u_inFIFO/n353 ), .B(n1206), .C(\u_inFIFO/n225 ), 
        .Q(\u_inFIFO/n352 ) );
  OAI212 \u_inFIFO/U258  ( .A(\u_inFIFO/n351 ), .B(n1206), .C(\u_inFIFO/n225 ), 
        .Q(\u_inFIFO/n350 ) );
  OAI212 \u_inFIFO/U256  ( .A(\u_inFIFO/n349 ), .B(n1206), .C(\u_inFIFO/n225 ), 
        .Q(\u_inFIFO/n348 ) );
  OAI212 \u_inFIFO/U254  ( .A(\u_inFIFO/n347 ), .B(n1206), .C(n1210), .Q(
        \u_inFIFO/n346 ) );
  OAI212 \u_inFIFO/U252  ( .A(\u_inFIFO/n345 ), .B(n1206), .C(n1210), .Q(
        \u_inFIFO/n344 ) );
  OAI212 \u_inFIFO/U250  ( .A(\u_inFIFO/n343 ), .B(n1206), .C(n1210), .Q(
        \u_inFIFO/n342 ) );
  OAI212 \u_inFIFO/U248  ( .A(\u_inFIFO/n340 ), .B(n1206), .C(n1210), .Q(
        \u_inFIFO/n339 ) );
  OAI212 \u_inFIFO/U245  ( .A(\u_inFIFO/n338 ), .B(n1206), .C(n1210), .Q(
        \u_inFIFO/n337 ) );
  OAI212 \u_inFIFO/U243  ( .A(\u_inFIFO/n336 ), .B(n1206), .C(n1210), .Q(
        \u_inFIFO/n335 ) );
  OAI212 \u_inFIFO/U241  ( .A(\u_inFIFO/n334 ), .B(n1206), .C(n1210), .Q(
        \u_inFIFO/n333 ) );
  OAI212 \u_inFIFO/U239  ( .A(\u_inFIFO/n332 ), .B(n1206), .C(n1210), .Q(
        \u_inFIFO/n331 ) );
  OAI212 \u_inFIFO/U237  ( .A(\u_inFIFO/n330 ), .B(n1206), .C(n1210), .Q(
        \u_inFIFO/n329 ) );
  OAI212 \u_inFIFO/U235  ( .A(\u_inFIFO/n328 ), .B(n1206), .C(n1210), .Q(
        \u_inFIFO/n327 ) );
  OAI212 \u_inFIFO/U233  ( .A(\u_inFIFO/n326 ), .B(n1206), .C(n1210), .Q(
        \u_inFIFO/n325 ) );
  OAI212 \u_inFIFO/U231  ( .A(\u_inFIFO/n324 ), .B(n1206), .C(n1210), .Q(
        \u_inFIFO/n323 ) );
  OAI212 \u_inFIFO/U229  ( .A(\u_inFIFO/n322 ), .B(n1206), .C(n1210), .Q(
        \u_inFIFO/n321 ) );
  OAI212 \u_inFIFO/U227  ( .A(\u_inFIFO/n320 ), .B(\u_inFIFO/n224 ), .C(n1210), 
        .Q(\u_inFIFO/n319 ) );
  OAI212 \u_inFIFO/U225  ( .A(\u_inFIFO/n318 ), .B(\u_inFIFO/n224 ), .C(n1210), 
        .Q(\u_inFIFO/n317 ) );
  OAI212 \u_inFIFO/U223  ( .A(\u_inFIFO/n316 ), .B(\u_inFIFO/n224 ), .C(n1210), 
        .Q(\u_inFIFO/n315 ) );
  OAI212 \u_inFIFO/U221  ( .A(\u_inFIFO/n314 ), .B(\u_inFIFO/n224 ), .C(n1210), 
        .Q(\u_inFIFO/n313 ) );
  OAI212 \u_inFIFO/U219  ( .A(\u_inFIFO/n312 ), .B(\u_inFIFO/n224 ), .C(n1210), 
        .Q(\u_inFIFO/n311 ) );
  OAI212 \u_inFIFO/U217  ( .A(\u_inFIFO/n310 ), .B(\u_inFIFO/n224 ), .C(n1210), 
        .Q(\u_inFIFO/n309 ) );
  OAI212 \u_inFIFO/U215  ( .A(\u_inFIFO/n307 ), .B(\u_inFIFO/n224 ), .C(n1210), 
        .Q(\u_inFIFO/n306 ) );
  OAI212 \u_inFIFO/U212  ( .A(\u_inFIFO/n305 ), .B(\u_inFIFO/n224 ), .C(n1210), 
        .Q(\u_inFIFO/n304 ) );
  OAI212 \u_inFIFO/U210  ( .A(\u_inFIFO/n303 ), .B(\u_inFIFO/n224 ), .C(n1210), 
        .Q(\u_inFIFO/n302 ) );
  OAI212 \u_inFIFO/U208  ( .A(\u_inFIFO/n301 ), .B(\u_inFIFO/n224 ), .C(n1210), 
        .Q(\u_inFIFO/n300 ) );
  OAI212 \u_inFIFO/U206  ( .A(\u_inFIFO/n299 ), .B(n1203), .C(n1210), .Q(
        \u_inFIFO/n298 ) );
  OAI212 \u_inFIFO/U204  ( .A(\u_inFIFO/n297 ), .B(n1206), .C(n1210), .Q(
        \u_inFIFO/n296 ) );
  OAI212 \u_inFIFO/U202  ( .A(\u_inFIFO/n295 ), .B(n1205), .C(n1210), .Q(
        \u_inFIFO/n294 ) );
  OAI212 \u_inFIFO/U200  ( .A(\u_inFIFO/n293 ), .B(n1204), .C(\u_inFIFO/n225 ), 
        .Q(\u_inFIFO/n292 ) );
  OAI212 \u_inFIFO/U198  ( .A(\u_inFIFO/n291 ), .B(n1208), .C(\u_inFIFO/n225 ), 
        .Q(\u_inFIFO/n290 ) );
  OAI212 \u_inFIFO/U196  ( .A(\u_inFIFO/n289 ), .B(n1207), .C(\u_inFIFO/n225 ), 
        .Q(\u_inFIFO/n288 ) );
  OAI212 \u_inFIFO/U194  ( .A(\u_inFIFO/n287 ), .B(n1208), .C(\u_inFIFO/n225 ), 
        .Q(\u_inFIFO/n286 ) );
  OAI212 \u_inFIFO/U192  ( .A(\u_inFIFO/n285 ), .B(n1207), .C(\u_inFIFO/n225 ), 
        .Q(\u_inFIFO/n284 ) );
  OAI212 \u_inFIFO/U190  ( .A(\u_inFIFO/n283 ), .B(n1207), .C(n1209), .Q(
        \u_inFIFO/n282 ) );
  OAI212 \u_inFIFO/U188  ( .A(\u_inFIFO/n281 ), .B(n1207), .C(n1210), .Q(
        \u_inFIFO/n280 ) );
  OAI212 \u_inFIFO/U186  ( .A(\u_inFIFO/n279 ), .B(n1207), .C(\u_inFIFO/n225 ), 
        .Q(\u_inFIFO/n278 ) );
  OAI212 \u_inFIFO/U184  ( .A(\u_inFIFO/n277 ), .B(n1207), .C(n1210), .Q(
        \u_inFIFO/n276 ) );
  OAI212 \u_inFIFO/U182  ( .A(\u_inFIFO/n274 ), .B(n1207), .C(\u_inFIFO/n225 ), 
        .Q(\u_inFIFO/n273 ) );
  OAI212 \u_inFIFO/U179  ( .A(\u_inFIFO/n271 ), .B(n1207), .C(n1210), .Q(
        \u_inFIFO/n270 ) );
  OAI212 \u_inFIFO/U177  ( .A(\u_inFIFO/n268 ), .B(n1207), .C(\u_inFIFO/n225 ), 
        .Q(\u_inFIFO/n267 ) );
  OAI212 \u_inFIFO/U175  ( .A(\u_inFIFO/n265 ), .B(n1207), .C(n1210), .Q(
        \u_inFIFO/n264 ) );
  OAI212 \u_inFIFO/U173  ( .A(\u_inFIFO/n262 ), .B(n1207), .C(\u_inFIFO/n225 ), 
        .Q(\u_inFIFO/n261 ) );
  OAI212 \u_inFIFO/U171  ( .A(\u_inFIFO/n259 ), .B(n1207), .C(n1210), .Q(
        \u_inFIFO/n258 ) );
  OAI212 \u_inFIFO/U169  ( .A(\u_inFIFO/n256 ), .B(n1207), .C(\u_inFIFO/n225 ), 
        .Q(\u_inFIFO/n255 ) );
  OAI212 \u_inFIFO/U167  ( .A(\u_inFIFO/n253 ), .B(n1207), .C(n1210), .Q(
        \u_inFIFO/n252 ) );
  OAI212 \u_inFIFO/U165  ( .A(\u_inFIFO/n250 ), .B(n1207), .C(\u_inFIFO/n225 ), 
        .Q(\u_inFIFO/n249 ) );
  OAI212 \u_inFIFO/U163  ( .A(\u_inFIFO/n247 ), .B(n1207), .C(n1210), .Q(
        \u_inFIFO/n246 ) );
  OAI212 \u_inFIFO/U161  ( .A(\u_inFIFO/n244 ), .B(n1207), .C(\u_inFIFO/n225 ), 
        .Q(\u_inFIFO/n243 ) );
  OAI212 \u_inFIFO/U159  ( .A(\u_inFIFO/n241 ), .B(n1207), .C(n1210), .Q(
        \u_inFIFO/n240 ) );
  OAI212 \u_inFIFO/U157  ( .A(\u_inFIFO/n238 ), .B(n1207), .C(\u_inFIFO/n225 ), 
        .Q(\u_inFIFO/n237 ) );
  OAI212 \u_inFIFO/U155  ( .A(\u_inFIFO/n235 ), .B(n1207), .C(n1210), .Q(
        \u_inFIFO/n234 ) );
  OAI212 \u_inFIFO/U153  ( .A(\u_inFIFO/n232 ), .B(n1208), .C(\u_inFIFO/n225 ), 
        .Q(\u_inFIFO/n231 ) );
  OAI212 \u_inFIFO/U151  ( .A(\u_inFIFO/n229 ), .B(n1208), .C(n1210), .Q(
        \u_inFIFO/n228 ) );
  OAI212 \u_inFIFO/U149  ( .A(\u_inFIFO/n223 ), .B(n1208), .C(\u_inFIFO/n225 ), 
        .Q(\u_inFIFO/n218 ) );
  OAI222 \u_inFIFO/U148  ( .A(n379), .B(\u_inFIFO/n216 ), .C(\u_inFIFO/n200 ), 
        .D(\u_inFIFO/n217 ), .Q(\u_inFIFO/n572 ) );
  OAI212 \u_coder/U199  ( .A(\u_coder/N1149 ), .B(\u_coder/n131 ), .C(
        \u_coder/n313 ), .Q(\u_coder/n356 ) );
  OAI212 \u_coder/U186  ( .A(\u_coder/IorQ ), .B(\u_coder/n307 ), .C(
        \u_coder/n308 ), .Q(\u_coder/n355 ) );
  OAI212 \u_coder/U183  ( .A(\u_coder/N1143 ), .B(\u_coder/n130 ), .C(
        \u_coder/n306 ), .Q(\u_coder/n354 ) );
  OAI212 \u_coder/U132  ( .A(\u_coder/n259 ), .B(\u_coder/n144 ), .C(
        \u_coder/n260 ), .Q(\u_coder/n257 ) );
  OAI222 \u_coder/U130  ( .A(\u_coder/n257 ), .B(\u_coder/n258 ), .C(n2160), 
        .D(n3112), .Q(\u_coder/n353 ) );
  OAI222 \u_coder/U123  ( .A(\u_coder/n126 ), .B(\u_coder/n254 ), .C(n2095), 
        .D(\u_coder/n167 ), .Q(\u_coder/n352 ) );
  OAI222 \u_coder/U122  ( .A(\u_coder/n123 ), .B(\u_coder/n255 ), .C(
        \u_coder/n126 ), .D(\u_coder/n139 ), .Q(\u_coder/n351 ) );
  OAI212 \u_coder/U119  ( .A(\u_coder/n251 ), .B(\u_coder/n246 ), .C(n2168), 
        .Q(\u_coder/n253 ) );
  OAI212 \u_coder/U109  ( .A(\u_coder/n243 ), .B(\u_coder/n144 ), .C(
        \u_coder/n244 ), .Q(\u_coder/n347 ) );
  OAI222 \u_coder/U100  ( .A(\u_coder/n125 ), .B(\u_coder/n239 ), .C(
        \u_coder/n127 ), .D(\u_coder/n182 ), .Q(\u_coder/n345 ) );
  OAI212 \u_coder/U95  ( .A(n2172), .B(n2174), .C(n2185), .Q(\u_coder/n233 )
         );
  OAI212 \u_coder/U85  ( .A(\u_coder/n226 ), .B(\u_coder/n183 ), .C(
        \u_coder/n227 ), .Q(\u_coder/n341 ) );
  OAI222 \u_coder/U78  ( .A(\u_coder/n181 ), .B(n2181), .C(\u_coder/n191 ), 
        .D(n2181), .Q(\u_coder/n219 ) );
  OAI222 \u_coder/U71  ( .A(\u_coder/n184 ), .B(n2181), .C(n2181), .D(
        \u_coder/n216 ), .Q(\u_coder/n214 ) );
  OAI212 \u_coder/U58  ( .A(\u_coder/n200 ), .B(\u_coder/n192 ), .C(
        \u_coder/n202 ), .Q(\u_coder/n198 ) );
  OAI222 \u_coder/U57  ( .A(\u_coder/n200 ), .B(\u_coder/n181 ), .C(
        \u_coder/n201 ), .D(\u_coder/n191 ), .Q(\u_coder/n199 ) );
  OAI212 \u_coder/U51  ( .A(\u_coder/n189 ), .B(\u_coder/n192 ), .C(
        \u_coder/n193 ), .Q(\u_coder/n187 ) );
  OAI222 \u_coder/U50  ( .A(\u_coder/n189 ), .B(\u_coder/n181 ), .C(
        \u_coder/n190 ), .D(\u_coder/n191 ), .Q(\u_coder/n188 ) );
  OAI222 \u_coder/U46  ( .A(\u_coder/n181 ), .B(\u_coder/n182 ), .C(
        \u_coder/n183 ), .D(\u_coder/n184 ), .Q(\u_coder/n180 ) );
  OAI212 \u_coder/U35  ( .A(\u_coder/n148 ), .B(n2155), .C(\u_coder/n158 ), 
        .Q(\u_coder/n138 ) );
  OAI212 \u_coder/U26  ( .A(\u_coder/n105 ), .B(\u_coder/n104 ), .C(
        \u_coder/i [2]), .Q(\u_coder/n160 ) );
  OAI222 \u_coder/U20  ( .A(n2165), .B(\u_coder/n147 ), .C(\u_coder/n148 ), 
        .D(n2155), .Q(\u_coder/n156 ) );
  OAI222 \u_coder/U18  ( .A(\u_coder/n153 ), .B(\u_coder/n139 ), .C(
        \u_coder/n154 ), .D(\u_coder/n144 ), .Q(\u_coder/n152 ) );
  OAI222 \u_coder/U14  ( .A(n2167), .B(\u_coder/n147 ), .C(\u_coder/n148 ), 
        .D(n2155), .Q(\u_coder/n146 ) );
  OAI222 \u_coder/U12  ( .A(\u_coder/n142 ), .B(\u_coder/n139 ), .C(
        \u_coder/n143 ), .D(\u_coder/n144 ), .Q(\u_coder/n141 ) );
  OAI212 \u_coder/U5  ( .A(\u_coder/n135 ), .B(\u_coder/n129 ), .C(
        \u_coder/n136 ), .Q(\u_coder/n335 ) );
  OAI212 \u_cordic/U23  ( .A(\u_cordic/present_state [2]), .B(n2107), .C(
        \u_cordic/n10 ), .Q(\u_cordic/n31 ) );
  OAI212 \u_cordic/U3  ( .A(\u_cordic/n15 ), .B(\u_cordic/n12 ), .C(
        \u_cordic/n16 ), .Q(\u_cordic/n32 ) );
  OAI222 \u_cdr/U35  ( .A(n289), .B(\u_cdr/n44 ), .C(n2210), .D(\u_cdr/n47 ), 
        .Q(\u_cdr/n59 ) );
  OAI222 \u_cdr/U34  ( .A(n20), .B(\u_cdr/n44 ), .C(n371), .D(\u_cdr/n47 ), 
        .Q(\u_cdr/n58 ) );
  OAI222 \u_cdr/U33  ( .A(n290), .B(\u_cdr/n44 ), .C(n372), .D(\u_cdr/n47 ), 
        .Q(\u_cdr/n57 ) );
  OAI222 \u_cdr/U32  ( .A(\u_cdr/n44 ), .B(n50), .C(\u_cdr/n46 ), .D(
        \u_cdr/n47 ), .Q(\u_cdr/n56 ) );
  OAI212 \u_cdr/U25  ( .A(\u_cdr/n43 ), .B(n1238), .C(\u_cdr/n44 ), .Q(
        \u_cdr/n27 ) );
  OAI222 \u_cdr/U23  ( .A(\u_cdr/cnt_d [0]), .B(\u_cdr/n24 ), .C(\u_cdr/n42 ), 
        .D(\u_cdr/n15 ), .Q(\u_cdr/n55 ) );
  OAI222 \u_cdr/U22  ( .A(n1232), .B(\u_cdr/n14 ), .C(\u_cdr/n24 ), .D(
        \u_cdr/n15 ), .Q(\u_cdr/n54 ) );
  OAI212 \u_cdr/U15  ( .A(\u_cdr/cnt [0]), .B(n1806), .C(\u_cdr/n35 ), .Q(
        \u_cdr/n34 ) );
  OAI212 \u_cdr/U12  ( .A(\u_cdr/n36 ), .B(\u_cdr/n16 ), .C(\u_cdr/n37 ), .Q(
        \u_cdr/n52 ) );
  OAI222 \u_cdr/U10  ( .A(n1805), .B(\u_cdr/n17 ), .C(\u_cdr/n18 ), .D(
        \u_cdr/n32 ), .Q(\u_cdr/n51 ) );
  OAI212 \u_cdr/U5  ( .A(\u_cdr/n26 ), .B(\u_cdr/n27 ), .C(\u_cdr/dir ), .Q(
        \u_cdr/n25 ) );
  OAI212 \u_outFIFO/U1095  ( .A(\u_outFIFO/currentState [1]), .B(
        \u_outFIFO/n1127 ), .C(\u_outFIFO/n1153 ), .Q(\u_outFIFO/n1158 ) );
  OAI212 \u_outFIFO/U1094  ( .A(\u_outFIFO/n1157 ), .B(n1240), .C(n1913), .Q(
        \u_outFIFO/N47 ) );
  OAI212 \u_outFIFO/U1088  ( .A(\u_outFIFO/n1152 ), .B(n1241), .C(
        \u_outFIFO/n1153 ), .Q(\u_outFIFO/N48 ) );
  OAI222 \u_outFIFO/U1087  ( .A(\u_outFIFO/N1269 ), .B(n2219), .C(n2224), .D(
        n2220), .Q(\u_outFIFO/n1151 ) );
  OAI212 \u_outFIFO/U1085  ( .A(\u_outFIFO/n1150 ), .B(n1240), .C(n1913), .Q(
        \u_outFIFO/N49 ) );
  OAI222 \u_outFIFO/U1078  ( .A(\u_outFIFO/n280 ), .B(n1796), .C(
        \u_outFIFO/n1143 ), .D(\u_outFIFO/i_FIFO [0]), .Q(\u_outFIFO/n1392 )
         );
  OAI222 \u_outFIFO/U1077  ( .A(\u_outFIFO/n279 ), .B(n1796), .C(
        \u_outFIFO/n1143 ), .D(n2236), .Q(\u_outFIFO/n1391 ) );
  OAI222 \u_outFIFO/U1076  ( .A(\u_outFIFO/n278 ), .B(n1796), .C(
        \u_outFIFO/n1143 ), .D(n2235), .Q(\u_outFIFO/n1390 ) );
  OAI222 \u_outFIFO/U1075  ( .A(\u_outFIFO/n277 ), .B(n1796), .C(
        \u_outFIFO/n1143 ), .D(n2234), .Q(\u_outFIFO/n1389 ) );
  OAI222 \u_outFIFO/U1074  ( .A(\u_outFIFO/n276 ), .B(n1796), .C(
        \u_outFIFO/n1143 ), .D(n2233), .Q(\u_outFIFO/n1388 ) );
  OAI222 \u_outFIFO/U1073  ( .A(\u_outFIFO/n275 ), .B(n1796), .C(
        \u_outFIFO/n1143 ), .D(n2232), .Q(\u_outFIFO/n1387 ) );
  OAI222 \u_outFIFO/U1072  ( .A(\u_outFIFO/n267 ), .B(n1796), .C(
        \u_outFIFO/n1143 ), .D(n376), .Q(\u_outFIFO/n1386 ) );
  OAI212 \u_outFIFO/U1068  ( .A(\u_outFIFO/sigEnableCounter ), .B(
        \u_outFIFO/n1127 ), .C(\u_outFIFO/n1128 ), .Q(\u_outFIFO/n1139 ) );
  OAI212 \u_outFIFO/U1064  ( .A(n1797), .B(\u_outFIFO/n258 ), .C(
        \u_outFIFO/n1138 ), .Q(\u_outFIFO/n1385 ) );
  OAI212 \u_outFIFO/U1062  ( .A(n1797), .B(\u_outFIFO/n266 ), .C(
        \u_outFIFO/n1137 ), .Q(\u_outFIFO/n1384 ) );
  OAI212 \u_outFIFO/U1060  ( .A(n1797), .B(\u_outFIFO/n265 ), .C(
        \u_outFIFO/n1136 ), .Q(\u_outFIFO/n1383 ) );
  OAI212 \u_outFIFO/U1058  ( .A(n1797), .B(\u_outFIFO/n264 ), .C(
        \u_outFIFO/n1135 ), .Q(\u_outFIFO/n1382 ) );
  OAI212 \u_outFIFO/U1056  ( .A(n1797), .B(\u_outFIFO/n263 ), .C(
        \u_outFIFO/n1134 ), .Q(\u_outFIFO/n1381 ) );
  OAI212 \u_outFIFO/U1054  ( .A(n1797), .B(\u_outFIFO/n262 ), .C(
        \u_outFIFO/n1133 ), .Q(\u_outFIFO/n1380 ) );
  OAI212 \u_outFIFO/U1052  ( .A(n1797), .B(\u_outFIFO/n261 ), .C(
        \u_outFIFO/n1132 ), .Q(\u_outFIFO/n1379 ) );
  OAI212 \u_outFIFO/U1050  ( .A(n1797), .B(\u_outFIFO/n260 ), .C(
        \u_outFIFO/n1130 ), .Q(\u_outFIFO/n1378 ) );
  OAI222 \u_outFIFO/U1035  ( .A(\u_outFIFO/n284 ), .B(n1191), .C(
        \u_outFIFO/n1116 ), .D(\u_outFIFO/n1112 ), .Q(\u_outFIFO/n1377 ) );
  OAI222 \u_outFIFO/U1032  ( .A(\u_outFIFO/n1113 ), .B(\u_outFIFO/n301 ), .C(
        \u_outFIFO/n1114 ), .D(n1180), .Q(\u_outFIFO/n1376 ) );
  OAI222 \u_outFIFO/U1031  ( .A(\u_outFIFO/n1113 ), .B(\u_outFIFO/n300 ), .C(
        \u_outFIFO/n1114 ), .D(n2216), .Q(\u_outFIFO/n1375 ) );
  OAI222 \u_outFIFO/U1030  ( .A(\u_outFIFO/n1113 ), .B(\u_outFIFO/n299 ), .C(
        \u_outFIFO/n1114 ), .D(n2215), .Q(\u_outFIFO/n1374 ) );
  OAI222 \u_outFIFO/U1029  ( .A(\u_outFIFO/n1113 ), .B(\u_outFIFO/n298 ), .C(
        \u_outFIFO/n1114 ), .D(n2214), .Q(\u_outFIFO/n1373 ) );
  OAI222 \u_outFIFO/U1028  ( .A(\u_outFIFO/n1113 ), .B(\u_outFIFO/n297 ), .C(
        \u_outFIFO/n1114 ), .D(n2213), .Q(\u_outFIFO/n1372 ) );
  OAI222 \u_outFIFO/U1027  ( .A(\u_outFIFO/n1113 ), .B(\u_outFIFO/n296 ), .C(
        \u_outFIFO/n1114 ), .D(n2212), .Q(\u_outFIFO/n1371 ) );
  OAI222 \u_outFIFO/U1026  ( .A(\u_outFIFO/n1113 ), .B(\u_outFIFO/n295 ), .C(
        \u_outFIFO/n1114 ), .D(n383), .Q(\u_outFIFO/n1370 ) );
  OAI212 \u_outFIFO/U1019  ( .A(\u_outFIFO/n396 ), .B(n885), .C(n927), .Q(
        \u_outFIFO/n1111 ) );
  OAI212 \u_outFIFO/U1016  ( .A(n1793), .B(n1184), .C(\u_outFIFO/FIFO[127][3] ), .Q(\u_outFIFO/n1109 ) );
  OAI212 \u_outFIFO/U1015  ( .A(n1793), .B(n1795), .C(\u_outFIFO/n1109 ), .Q(
        \u_outFIFO/n1369 ) );
  OAI212 \u_outFIFO/U1013  ( .A(\u_outFIFO/n396 ), .B(n882), .C(n951), .Q(
        \u_outFIFO/n1108 ) );
  OAI212 \u_outFIFO/U1012  ( .A(n1792), .B(n1185), .C(\u_outFIFO/FIFO[127][2] ), .Q(\u_outFIFO/n1107 ) );
  OAI212 \u_outFIFO/U1011  ( .A(n1792), .B(n1795), .C(\u_outFIFO/n1107 ), .Q(
        \u_outFIFO/n1368 ) );
  OAI212 \u_outFIFO/U1009  ( .A(\u_outFIFO/n396 ), .B(n880), .C(n951), .Q(
        \u_outFIFO/n1106 ) );
  OAI212 \u_outFIFO/U1008  ( .A(n1791), .B(n1189), .C(\u_outFIFO/FIFO[127][1] ), .Q(\u_outFIFO/n1105 ) );
  OAI212 \u_outFIFO/U1007  ( .A(n1791), .B(n1795), .C(\u_outFIFO/n1105 ), .Q(
        \u_outFIFO/n1367 ) );
  OAI212 \u_outFIFO/U1005  ( .A(\u_outFIFO/n396 ), .B(n878), .C(n951), .Q(
        \u_outFIFO/n1103 ) );
  OAI212 \u_outFIFO/U1004  ( .A(n1790), .B(n1188), .C(\u_outFIFO/FIFO[127][0] ), .Q(\u_outFIFO/n1102 ) );
  OAI212 \u_outFIFO/U1003  ( .A(n1790), .B(n1795), .C(\u_outFIFO/n1102 ), .Q(
        \u_outFIFO/n1366 ) );
  OAI212 \u_outFIFO/U1000  ( .A(\u_outFIFO/n391 ), .B(n885), .C(n951), .Q(
        \u_outFIFO/n1101 ) );
  OAI212 \u_outFIFO/U999  ( .A(n1789), .B(n1186), .C(\u_outFIFO/FIFO[126][3] ), 
        .Q(\u_outFIFO/n1100 ) );
  OAI212 \u_outFIFO/U998  ( .A(n1789), .B(n1795), .C(\u_outFIFO/n1100 ), .Q(
        \u_outFIFO/n1365 ) );
  OAI212 \u_outFIFO/U997  ( .A(\u_outFIFO/n391 ), .B(n882), .C(n951), .Q(
        \u_outFIFO/n1099 ) );
  OAI212 \u_outFIFO/U996  ( .A(n1788), .B(n1185), .C(\u_outFIFO/FIFO[126][2] ), 
        .Q(\u_outFIFO/n1098 ) );
  OAI212 \u_outFIFO/U995  ( .A(n1788), .B(n1795), .C(\u_outFIFO/n1098 ), .Q(
        \u_outFIFO/n1364 ) );
  OAI212 \u_outFIFO/U994  ( .A(\u_outFIFO/n391 ), .B(n880), .C(n951), .Q(
        \u_outFIFO/n1097 ) );
  OAI212 \u_outFIFO/U993  ( .A(n1787), .B(n1185), .C(\u_outFIFO/FIFO[126][1] ), 
        .Q(\u_outFIFO/n1096 ) );
  OAI212 \u_outFIFO/U992  ( .A(n1787), .B(n1795), .C(\u_outFIFO/n1096 ), .Q(
        \u_outFIFO/n1363 ) );
  OAI212 \u_outFIFO/U991  ( .A(\u_outFIFO/n391 ), .B(n878), .C(n951), .Q(
        \u_outFIFO/n1095 ) );
  OAI212 \u_outFIFO/U990  ( .A(n1786), .B(n1187), .C(\u_outFIFO/FIFO[126][0] ), 
        .Q(\u_outFIFO/n1094 ) );
  OAI212 \u_outFIFO/U989  ( .A(n1786), .B(n1795), .C(\u_outFIFO/n1094 ), .Q(
        \u_outFIFO/n1362 ) );
  OAI212 \u_outFIFO/U986  ( .A(\u_outFIFO/n386 ), .B(n885), .C(n951), .Q(
        \u_outFIFO/n1093 ) );
  OAI212 \u_outFIFO/U985  ( .A(n1785), .B(n1187), .C(\u_outFIFO/FIFO[125][3] ), 
        .Q(\u_outFIFO/n1092 ) );
  OAI212 \u_outFIFO/U984  ( .A(n1785), .B(n1795), .C(\u_outFIFO/n1092 ), .Q(
        \u_outFIFO/n1361 ) );
  OAI212 \u_outFIFO/U983  ( .A(\u_outFIFO/n386 ), .B(n882), .C(n950), .Q(
        \u_outFIFO/n1091 ) );
  OAI212 \u_outFIFO/U982  ( .A(n1784), .B(n1189), .C(\u_outFIFO/FIFO[125][2] ), 
        .Q(\u_outFIFO/n1090 ) );
  OAI212 \u_outFIFO/U981  ( .A(n1784), .B(n1795), .C(\u_outFIFO/n1090 ), .Q(
        \u_outFIFO/n1360 ) );
  OAI212 \u_outFIFO/U980  ( .A(\u_outFIFO/n386 ), .B(n880), .C(n950), .Q(
        \u_outFIFO/n1089 ) );
  OAI212 \u_outFIFO/U979  ( .A(n1783), .B(n1190), .C(\u_outFIFO/FIFO[125][1] ), 
        .Q(\u_outFIFO/n1088 ) );
  OAI212 \u_outFIFO/U978  ( .A(n1783), .B(n1795), .C(\u_outFIFO/n1088 ), .Q(
        \u_outFIFO/n1359 ) );
  OAI212 \u_outFIFO/U977  ( .A(\u_outFIFO/n386 ), .B(n878), .C(n950), .Q(
        \u_outFIFO/n1087 ) );
  OAI212 \u_outFIFO/U976  ( .A(n1782), .B(n1188), .C(\u_outFIFO/FIFO[125][0] ), 
        .Q(\u_outFIFO/n1086 ) );
  OAI212 \u_outFIFO/U975  ( .A(n1782), .B(n1795), .C(\u_outFIFO/n1086 ), .Q(
        \u_outFIFO/n1358 ) );
  OAI212 \u_outFIFO/U972  ( .A(n873), .B(n885), .C(n950), .Q(\u_outFIFO/n1084 ) );
  OAI212 \u_outFIFO/U971  ( .A(n1781), .B(n1187), .C(\u_outFIFO/FIFO[124][3] ), 
        .Q(\u_outFIFO/n1083 ) );
  OAI212 \u_outFIFO/U970  ( .A(n1781), .B(n1795), .C(\u_outFIFO/n1083 ), .Q(
        \u_outFIFO/n1357 ) );
  OAI212 \u_outFIFO/U969  ( .A(\u_outFIFO/n381 ), .B(n882), .C(n950), .Q(
        \u_outFIFO/n1082 ) );
  OAI212 \u_outFIFO/U968  ( .A(n1780), .B(n1188), .C(\u_outFIFO/FIFO[124][2] ), 
        .Q(\u_outFIFO/n1081 ) );
  OAI212 \u_outFIFO/U967  ( .A(n1780), .B(n960), .C(\u_outFIFO/n1081 ), .Q(
        \u_outFIFO/n1356 ) );
  OAI212 \u_outFIFO/U966  ( .A(\u_outFIFO/n381 ), .B(n880), .C(n950), .Q(
        \u_outFIFO/n1080 ) );
  OAI212 \u_outFIFO/U965  ( .A(n1779), .B(n1189), .C(\u_outFIFO/FIFO[124][1] ), 
        .Q(\u_outFIFO/n1079 ) );
  OAI212 \u_outFIFO/U964  ( .A(n1779), .B(n952), .C(\u_outFIFO/n1079 ), .Q(
        \u_outFIFO/n1355 ) );
  OAI212 \u_outFIFO/U963  ( .A(\u_outFIFO/n381 ), .B(n878), .C(n950), .Q(
        \u_outFIFO/n1078 ) );
  OAI212 \u_outFIFO/U962  ( .A(n1778), .B(n1190), .C(\u_outFIFO/FIFO[124][0] ), 
        .Q(\u_outFIFO/n1077 ) );
  OAI212 \u_outFIFO/U961  ( .A(n1778), .B(n1795), .C(\u_outFIFO/n1077 ), .Q(
        \u_outFIFO/n1354 ) );
  OAI212 \u_outFIFO/U958  ( .A(n869), .B(n885), .C(n950), .Q(\u_outFIFO/n1076 ) );
  OAI212 \u_outFIFO/U957  ( .A(n1777), .B(n1185), .C(\u_outFIFO/FIFO[123][3] ), 
        .Q(\u_outFIFO/n1075 ) );
  OAI212 \u_outFIFO/U956  ( .A(n1777), .B(n1795), .C(\u_outFIFO/n1075 ), .Q(
        \u_outFIFO/n1353 ) );
  OAI212 \u_outFIFO/U955  ( .A(n869), .B(n882), .C(n949), .Q(\u_outFIFO/n1074 ) );
  OAI212 \u_outFIFO/U954  ( .A(n1776), .B(n1186), .C(\u_outFIFO/FIFO[123][2] ), 
        .Q(\u_outFIFO/n1073 ) );
  OAI212 \u_outFIFO/U953  ( .A(n1776), .B(n1795), .C(\u_outFIFO/n1073 ), .Q(
        \u_outFIFO/n1352 ) );
  OAI212 \u_outFIFO/U952  ( .A(n869), .B(n880), .C(n949), .Q(\u_outFIFO/n1072 ) );
  OAI212 \u_outFIFO/U951  ( .A(n1775), .B(n1190), .C(\u_outFIFO/FIFO[123][1] ), 
        .Q(\u_outFIFO/n1071 ) );
  OAI212 \u_outFIFO/U950  ( .A(n1775), .B(n1795), .C(\u_outFIFO/n1071 ), .Q(
        \u_outFIFO/n1351 ) );
  OAI212 \u_outFIFO/U949  ( .A(n869), .B(n878), .C(n949), .Q(\u_outFIFO/n1070 ) );
  OAI212 \u_outFIFO/U948  ( .A(n1774), .B(n1187), .C(\u_outFIFO/FIFO[123][0] ), 
        .Q(\u_outFIFO/n1069 ) );
  OAI212 \u_outFIFO/U947  ( .A(n1774), .B(n1795), .C(\u_outFIFO/n1069 ), .Q(
        \u_outFIFO/n1350 ) );
  OAI212 \u_outFIFO/U945  ( .A(n866), .B(n885), .C(n949), .Q(\u_outFIFO/n1068 ) );
  OAI212 \u_outFIFO/U944  ( .A(n1773), .B(n1188), .C(\u_outFIFO/FIFO[122][3] ), 
        .Q(\u_outFIFO/n1067 ) );
  OAI212 \u_outFIFO/U943  ( .A(n1773), .B(n1795), .C(\u_outFIFO/n1067 ), .Q(
        \u_outFIFO/n1349 ) );
  OAI212 \u_outFIFO/U942  ( .A(n866), .B(n882), .C(n949), .Q(\u_outFIFO/n1066 ) );
  OAI212 \u_outFIFO/U941  ( .A(n1772), .B(n1189), .C(\u_outFIFO/FIFO[122][2] ), 
        .Q(\u_outFIFO/n1065 ) );
  OAI212 \u_outFIFO/U940  ( .A(n1772), .B(n1795), .C(\u_outFIFO/n1065 ), .Q(
        \u_outFIFO/n1348 ) );
  OAI212 \u_outFIFO/U939  ( .A(n866), .B(n880), .C(n949), .Q(\u_outFIFO/n1064 ) );
  OAI212 \u_outFIFO/U938  ( .A(n1771), .B(n1190), .C(\u_outFIFO/FIFO[122][1] ), 
        .Q(\u_outFIFO/n1063 ) );
  OAI212 \u_outFIFO/U937  ( .A(n1771), .B(n1795), .C(\u_outFIFO/n1063 ), .Q(
        \u_outFIFO/n1347 ) );
  OAI212 \u_outFIFO/U936  ( .A(n866), .B(n878), .C(n949), .Q(\u_outFIFO/n1062 ) );
  OAI212 \u_outFIFO/U935  ( .A(n1770), .B(n1185), .C(\u_outFIFO/FIFO[122][0] ), 
        .Q(\u_outFIFO/n1061 ) );
  OAI212 \u_outFIFO/U934  ( .A(n1770), .B(n1795), .C(\u_outFIFO/n1061 ), .Q(
        \u_outFIFO/n1346 ) );
  OAI212 \u_outFIFO/U932  ( .A(n863), .B(n887), .C(n949), .Q(\u_outFIFO/n1060 ) );
  OAI212 \u_outFIFO/U931  ( .A(n1769), .B(n1186), .C(\u_outFIFO/FIFO[121][3] ), 
        .Q(\u_outFIFO/n1059 ) );
  OAI212 \u_outFIFO/U930  ( .A(n1769), .B(n1795), .C(\u_outFIFO/n1059 ), .Q(
        \u_outFIFO/n1345 ) );
  OAI212 \u_outFIFO/U929  ( .A(n863), .B(n884), .C(n948), .Q(\u_outFIFO/n1058 ) );
  OAI212 \u_outFIFO/U928  ( .A(n1768), .B(n1186), .C(\u_outFIFO/FIFO[121][2] ), 
        .Q(\u_outFIFO/n1057 ) );
  OAI212 \u_outFIFO/U927  ( .A(n1768), .B(n1795), .C(\u_outFIFO/n1057 ), .Q(
        \u_outFIFO/n1344 ) );
  OAI212 \u_outFIFO/U926  ( .A(n863), .B(n880), .C(n948), .Q(\u_outFIFO/n1056 ) );
  OAI212 \u_outFIFO/U925  ( .A(n1767), .B(n1187), .C(\u_outFIFO/FIFO[121][1] ), 
        .Q(\u_outFIFO/n1055 ) );
  OAI212 \u_outFIFO/U924  ( .A(n1767), .B(n953), .C(\u_outFIFO/n1055 ), .Q(
        \u_outFIFO/n1343 ) );
  OAI212 \u_outFIFO/U923  ( .A(n863), .B(n878), .C(n948), .Q(\u_outFIFO/n1054 ) );
  OAI212 \u_outFIFO/U922  ( .A(n1766), .B(n1188), .C(\u_outFIFO/FIFO[121][0] ), 
        .Q(\u_outFIFO/n1053 ) );
  OAI212 \u_outFIFO/U921  ( .A(n1766), .B(n952), .C(\u_outFIFO/n1053 ), .Q(
        \u_outFIFO/n1342 ) );
  OAI212 \u_outFIFO/U919  ( .A(n860), .B(n886), .C(n948), .Q(\u_outFIFO/n1051 ) );
  OAI212 \u_outFIFO/U918  ( .A(n1765), .B(n1189), .C(\u_outFIFO/FIFO[120][3] ), 
        .Q(\u_outFIFO/n1050 ) );
  OAI212 \u_outFIFO/U917  ( .A(n1765), .B(n953), .C(\u_outFIFO/n1050 ), .Q(
        \u_outFIFO/n1341 ) );
  OAI212 \u_outFIFO/U916  ( .A(n860), .B(n883), .C(n948), .Q(\u_outFIFO/n1049 ) );
  OAI212 \u_outFIFO/U915  ( .A(n1764), .B(n1189), .C(\u_outFIFO/FIFO[120][2] ), 
        .Q(\u_outFIFO/n1048 ) );
  OAI212 \u_outFIFO/U914  ( .A(n1764), .B(n961), .C(\u_outFIFO/n1048 ), .Q(
        \u_outFIFO/n1340 ) );
  OAI212 \u_outFIFO/U913  ( .A(n860), .B(n880), .C(n948), .Q(\u_outFIFO/n1047 ) );
  OAI212 \u_outFIFO/U912  ( .A(n1763), .B(n1189), .C(\u_outFIFO/FIFO[120][1] ), 
        .Q(\u_outFIFO/n1046 ) );
  OAI212 \u_outFIFO/U911  ( .A(n1763), .B(n960), .C(\u_outFIFO/n1046 ), .Q(
        \u_outFIFO/n1339 ) );
  OAI212 \u_outFIFO/U910  ( .A(n860), .B(n878), .C(n948), .Q(\u_outFIFO/n1045 ) );
  OAI212 \u_outFIFO/U909  ( .A(n1762), .B(n1189), .C(\u_outFIFO/FIFO[120][0] ), 
        .Q(\u_outFIFO/n1044 ) );
  OAI212 \u_outFIFO/U908  ( .A(n1762), .B(n959), .C(\u_outFIFO/n1044 ), .Q(
        \u_outFIFO/n1338 ) );
  OAI212 \u_outFIFO/U905  ( .A(n857), .B(n887), .C(n948), .Q(\u_outFIFO/n1043 ) );
  OAI212 \u_outFIFO/U904  ( .A(n1761), .B(n1189), .C(\u_outFIFO/FIFO[119][3] ), 
        .Q(\u_outFIFO/n1042 ) );
  OAI212 \u_outFIFO/U903  ( .A(n1761), .B(n958), .C(\u_outFIFO/n1042 ), .Q(
        \u_outFIFO/n1337 ) );
  OAI212 \u_outFIFO/U902  ( .A(n857), .B(n884), .C(n947), .Q(\u_outFIFO/n1041 ) );
  OAI212 \u_outFIFO/U901  ( .A(n1760), .B(n1189), .C(\u_outFIFO/FIFO[119][2] ), 
        .Q(\u_outFIFO/n1040 ) );
  OAI212 \u_outFIFO/U900  ( .A(n1760), .B(n957), .C(\u_outFIFO/n1040 ), .Q(
        \u_outFIFO/n1336 ) );
  OAI212 \u_outFIFO/U899  ( .A(n857), .B(n881), .C(n947), .Q(\u_outFIFO/n1039 ) );
  OAI212 \u_outFIFO/U898  ( .A(n1759), .B(n1189), .C(\u_outFIFO/FIFO[119][1] ), 
        .Q(\u_outFIFO/n1038 ) );
  OAI212 \u_outFIFO/U897  ( .A(n1759), .B(n956), .C(\u_outFIFO/n1038 ), .Q(
        \u_outFIFO/n1335 ) );
  OAI212 \u_outFIFO/U896  ( .A(n857), .B(n879), .C(n947), .Q(\u_outFIFO/n1037 ) );
  OAI212 \u_outFIFO/U895  ( .A(n1758), .B(n1189), .C(\u_outFIFO/FIFO[119][0] ), 
        .Q(\u_outFIFO/n1036 ) );
  OAI212 \u_outFIFO/U894  ( .A(n1758), .B(n955), .C(\u_outFIFO/n1036 ), .Q(
        \u_outFIFO/n1334 ) );
  OAI212 \u_outFIFO/U892  ( .A(n854), .B(n886), .C(n947), .Q(\u_outFIFO/n1035 ) );
  OAI212 \u_outFIFO/U891  ( .A(n1757), .B(n1189), .C(\u_outFIFO/FIFO[118][3] ), 
        .Q(\u_outFIFO/n1034 ) );
  OAI212 \u_outFIFO/U890  ( .A(n1757), .B(n954), .C(\u_outFIFO/n1034 ), .Q(
        \u_outFIFO/n1333 ) );
  OAI212 \u_outFIFO/U889  ( .A(n854), .B(n883), .C(n947), .Q(\u_outFIFO/n1033 ) );
  OAI212 \u_outFIFO/U888  ( .A(n1756), .B(n1189), .C(\u_outFIFO/FIFO[118][2] ), 
        .Q(\u_outFIFO/n1032 ) );
  OAI212 \u_outFIFO/U887  ( .A(n1756), .B(n953), .C(\u_outFIFO/n1032 ), .Q(
        \u_outFIFO/n1332 ) );
  OAI212 \u_outFIFO/U886  ( .A(n854), .B(n881), .C(n947), .Q(\u_outFIFO/n1031 ) );
  OAI212 \u_outFIFO/U885  ( .A(n1755), .B(n1189), .C(\u_outFIFO/FIFO[118][1] ), 
        .Q(\u_outFIFO/n1030 ) );
  OAI212 \u_outFIFO/U884  ( .A(n1755), .B(n952), .C(\u_outFIFO/n1030 ), .Q(
        \u_outFIFO/n1331 ) );
  OAI212 \u_outFIFO/U883  ( .A(n854), .B(n879), .C(n947), .Q(\u_outFIFO/n1029 ) );
  OAI212 \u_outFIFO/U882  ( .A(n1754), .B(n1189), .C(\u_outFIFO/FIFO[118][0] ), 
        .Q(\u_outFIFO/n1028 ) );
  OAI212 \u_outFIFO/U881  ( .A(n1754), .B(n953), .C(\u_outFIFO/n1028 ), .Q(
        \u_outFIFO/n1330 ) );
  OAI212 \u_outFIFO/U879  ( .A(n851), .B(n887), .C(n947), .Q(\u_outFIFO/n1027 ) );
  OAI212 \u_outFIFO/U878  ( .A(n1753), .B(n1189), .C(\u_outFIFO/FIFO[117][3] ), 
        .Q(\u_outFIFO/n1026 ) );
  OAI212 \u_outFIFO/U877  ( .A(n1753), .B(n952), .C(\u_outFIFO/n1026 ), .Q(
        \u_outFIFO/n1329 ) );
  OAI212 \u_outFIFO/U876  ( .A(n851), .B(n884), .C(n946), .Q(\u_outFIFO/n1025 ) );
  OAI212 \u_outFIFO/U875  ( .A(n1752), .B(n1189), .C(\u_outFIFO/FIFO[117][2] ), 
        .Q(\u_outFIFO/n1024 ) );
  OAI212 \u_outFIFO/U874  ( .A(n1752), .B(n959), .C(\u_outFIFO/n1024 ), .Q(
        \u_outFIFO/n1328 ) );
  OAI212 \u_outFIFO/U873  ( .A(n851), .B(n881), .C(n946), .Q(\u_outFIFO/n1023 ) );
  OAI212 \u_outFIFO/U872  ( .A(n1751), .B(n1189), .C(\u_outFIFO/FIFO[117][1] ), 
        .Q(\u_outFIFO/n1022 ) );
  OAI212 \u_outFIFO/U871  ( .A(n1751), .B(n958), .C(\u_outFIFO/n1022 ), .Q(
        \u_outFIFO/n1327 ) );
  OAI212 \u_outFIFO/U870  ( .A(n851), .B(n879), .C(n946), .Q(\u_outFIFO/n1021 ) );
  OAI212 \u_outFIFO/U869  ( .A(n1750), .B(n1189), .C(\u_outFIFO/FIFO[117][0] ), 
        .Q(\u_outFIFO/n1020 ) );
  OAI212 \u_outFIFO/U868  ( .A(n1750), .B(n957), .C(\u_outFIFO/n1020 ), .Q(
        \u_outFIFO/n1326 ) );
  OAI212 \u_outFIFO/U866  ( .A(n848), .B(n886), .C(n946), .Q(\u_outFIFO/n1018 ) );
  OAI212 \u_outFIFO/U865  ( .A(n1749), .B(n1189), .C(\u_outFIFO/FIFO[116][3] ), 
        .Q(\u_outFIFO/n1017 ) );
  OAI212 \u_outFIFO/U864  ( .A(n1749), .B(n956), .C(\u_outFIFO/n1017 ), .Q(
        \u_outFIFO/n1325 ) );
  OAI212 \u_outFIFO/U863  ( .A(n848), .B(n883), .C(n946), .Q(\u_outFIFO/n1016 ) );
  OAI212 \u_outFIFO/U862  ( .A(n1748), .B(n1189), .C(\u_outFIFO/FIFO[116][2] ), 
        .Q(\u_outFIFO/n1015 ) );
  OAI212 \u_outFIFO/U861  ( .A(n1748), .B(n955), .C(\u_outFIFO/n1015 ), .Q(
        \u_outFIFO/n1324 ) );
  OAI212 \u_outFIFO/U860  ( .A(n848), .B(n881), .C(n946), .Q(\u_outFIFO/n1014 ) );
  OAI212 \u_outFIFO/U859  ( .A(n1747), .B(n1185), .C(\u_outFIFO/FIFO[116][1] ), 
        .Q(\u_outFIFO/n1013 ) );
  OAI212 \u_outFIFO/U858  ( .A(n1747), .B(n954), .C(\u_outFIFO/n1013 ), .Q(
        \u_outFIFO/n1323 ) );
  OAI212 \u_outFIFO/U857  ( .A(n848), .B(n879), .C(n946), .Q(\u_outFIFO/n1012 ) );
  OAI212 \u_outFIFO/U856  ( .A(n1746), .B(n1187), .C(\u_outFIFO/FIFO[116][0] ), 
        .Q(\u_outFIFO/n1011 ) );
  OAI212 \u_outFIFO/U855  ( .A(n1746), .B(n961), .C(\u_outFIFO/n1011 ), .Q(
        \u_outFIFO/n1322 ) );
  OAI212 \u_outFIFO/U852  ( .A(n844), .B(n887), .C(n946), .Q(\u_outFIFO/n1009 ) );
  OAI212 \u_outFIFO/U851  ( .A(n1745), .B(n1187), .C(\u_outFIFO/FIFO[115][3] ), 
        .Q(\u_outFIFO/n1008 ) );
  OAI212 \u_outFIFO/U850  ( .A(n1745), .B(n960), .C(\u_outFIFO/n1008 ), .Q(
        \u_outFIFO/n1321 ) );
  OAI212 \u_outFIFO/U849  ( .A(n845), .B(n884), .C(n945), .Q(\u_outFIFO/n1007 ) );
  OAI212 \u_outFIFO/U848  ( .A(n1744), .B(n1188), .C(\u_outFIFO/FIFO[115][2] ), 
        .Q(\u_outFIFO/n1006 ) );
  OAI212 \u_outFIFO/U847  ( .A(n1744), .B(n953), .C(\u_outFIFO/n1006 ), .Q(
        \u_outFIFO/n1320 ) );
  OAI212 \u_outFIFO/U846  ( .A(n846), .B(n881), .C(n945), .Q(\u_outFIFO/n1005 ) );
  OAI212 \u_outFIFO/U845  ( .A(n1743), .B(n1188), .C(\u_outFIFO/FIFO[115][1] ), 
        .Q(\u_outFIFO/n1004 ) );
  OAI212 \u_outFIFO/U844  ( .A(n1743), .B(n952), .C(\u_outFIFO/n1004 ), .Q(
        \u_outFIFO/n1319 ) );
  OAI212 \u_outFIFO/U843  ( .A(n847), .B(n879), .C(n945), .Q(\u_outFIFO/n1003 ) );
  OAI212 \u_outFIFO/U842  ( .A(n1742), .B(n1189), .C(\u_outFIFO/FIFO[115][0] ), 
        .Q(\u_outFIFO/n1002 ) );
  OAI212 \u_outFIFO/U841  ( .A(n1742), .B(n961), .C(\u_outFIFO/n1002 ), .Q(
        \u_outFIFO/n1318 ) );
  OAI212 \u_outFIFO/U839  ( .A(\u_outFIFO/n331 ), .B(n886), .C(n945), .Q(
        \u_outFIFO/n1000 ) );
  OAI212 \u_outFIFO/U838  ( .A(n1741), .B(n1190), .C(\u_outFIFO/FIFO[114][3] ), 
        .Q(\u_outFIFO/n999 ) );
  OAI212 \u_outFIFO/U837  ( .A(n1741), .B(n955), .C(\u_outFIFO/n999 ), .Q(
        \u_outFIFO/n1317 ) );
  OAI212 \u_outFIFO/U836  ( .A(\u_outFIFO/n331 ), .B(n883), .C(n945), .Q(
        \u_outFIFO/n998 ) );
  OAI212 \u_outFIFO/U835  ( .A(n1740), .B(n1186), .C(\u_outFIFO/FIFO[114][2] ), 
        .Q(\u_outFIFO/n997 ) );
  OAI212 \u_outFIFO/U834  ( .A(n1740), .B(n1795), .C(\u_outFIFO/n997 ), .Q(
        \u_outFIFO/n1316 ) );
  OAI212 \u_outFIFO/U833  ( .A(\u_outFIFO/n331 ), .B(n881), .C(n945), .Q(
        \u_outFIFO/n996 ) );
  OAI212 \u_outFIFO/U832  ( .A(n1739), .B(n1188), .C(\u_outFIFO/FIFO[114][1] ), 
        .Q(\u_outFIFO/n995 ) );
  OAI212 \u_outFIFO/U831  ( .A(n1739), .B(n961), .C(\u_outFIFO/n995 ), .Q(
        \u_outFIFO/n1315 ) );
  OAI212 \u_outFIFO/U830  ( .A(n842), .B(n879), .C(n945), .Q(\u_outFIFO/n994 )
         );
  OAI212 \u_outFIFO/U829  ( .A(n1738), .B(n1187), .C(\u_outFIFO/FIFO[114][0] ), 
        .Q(\u_outFIFO/n993 ) );
  OAI212 \u_outFIFO/U828  ( .A(n1738), .B(n960), .C(\u_outFIFO/n993 ), .Q(
        \u_outFIFO/n1314 ) );
  OAI212 \u_outFIFO/U826  ( .A(n838), .B(n887), .C(n945), .Q(\u_outFIFO/n991 )
         );
  OAI212 \u_outFIFO/U825  ( .A(n1737), .B(n1188), .C(\u_outFIFO/FIFO[113][3] ), 
        .Q(\u_outFIFO/n990 ) );
  OAI212 \u_outFIFO/U824  ( .A(n1737), .B(n959), .C(\u_outFIFO/n990 ), .Q(
        \u_outFIFO/n1313 ) );
  OAI212 \u_outFIFO/U823  ( .A(n838), .B(n884), .C(n944), .Q(\u_outFIFO/n989 )
         );
  OAI212 \u_outFIFO/U822  ( .A(n1736), .B(n1189), .C(\u_outFIFO/FIFO[113][2] ), 
        .Q(\u_outFIFO/n988 ) );
  OAI212 \u_outFIFO/U821  ( .A(n1736), .B(n958), .C(\u_outFIFO/n988 ), .Q(
        \u_outFIFO/n1312 ) );
  OAI212 \u_outFIFO/U820  ( .A(n838), .B(n881), .C(n944), .Q(\u_outFIFO/n987 )
         );
  OAI212 \u_outFIFO/U819  ( .A(n1735), .B(n1189), .C(\u_outFIFO/FIFO[113][1] ), 
        .Q(\u_outFIFO/n986 ) );
  OAI212 \u_outFIFO/U818  ( .A(n1735), .B(n957), .C(\u_outFIFO/n986 ), .Q(
        \u_outFIFO/n1311 ) );
  OAI212 \u_outFIFO/U817  ( .A(n838), .B(n879), .C(n944), .Q(\u_outFIFO/n985 )
         );
  OAI212 \u_outFIFO/U816  ( .A(n1734), .B(n1190), .C(\u_outFIFO/FIFO[113][0] ), 
        .Q(\u_outFIFO/n984 ) );
  OAI212 \u_outFIFO/U815  ( .A(n1734), .B(n956), .C(\u_outFIFO/n984 ), .Q(
        \u_outFIFO/n1310 ) );
  OAI212 \u_outFIFO/U813  ( .A(\u_outFIFO/n317 ), .B(n886), .C(n944), .Q(
        \u_outFIFO/n980 ) );
  OAI212 \u_outFIFO/U812  ( .A(n1733), .B(n1189), .C(\u_outFIFO/FIFO[112][3] ), 
        .Q(\u_outFIFO/n979 ) );
  OAI212 \u_outFIFO/U811  ( .A(n1733), .B(n955), .C(\u_outFIFO/n979 ), .Q(
        \u_outFIFO/n1309 ) );
  OAI212 \u_outFIFO/U810  ( .A(\u_outFIFO/n317 ), .B(n883), .C(n944), .Q(
        \u_outFIFO/n977 ) );
  OAI212 \u_outFIFO/U809  ( .A(n1732), .B(n1187), .C(\u_outFIFO/FIFO[112][2] ), 
        .Q(\u_outFIFO/n976 ) );
  OAI212 \u_outFIFO/U808  ( .A(n1732), .B(n954), .C(\u_outFIFO/n976 ), .Q(
        \u_outFIFO/n1308 ) );
  OAI212 \u_outFIFO/U807  ( .A(n837), .B(n881), .C(n944), .Q(\u_outFIFO/n974 )
         );
  OAI212 \u_outFIFO/U806  ( .A(n1731), .B(n1186), .C(\u_outFIFO/FIFO[112][1] ), 
        .Q(\u_outFIFO/n973 ) );
  OAI212 \u_outFIFO/U805  ( .A(n1731), .B(n953), .C(\u_outFIFO/n973 ), .Q(
        \u_outFIFO/n1307 ) );
  OAI212 \u_outFIFO/U804  ( .A(n837), .B(n879), .C(n944), .Q(\u_outFIFO/n971 )
         );
  OAI212 \u_outFIFO/U803  ( .A(n1730), .B(n1189), .C(\u_outFIFO/FIFO[112][0] ), 
        .Q(\u_outFIFO/n970 ) );
  OAI212 \u_outFIFO/U802  ( .A(n1730), .B(n952), .C(\u_outFIFO/n970 ), .Q(
        \u_outFIFO/n1306 ) );
  OAI212 \u_outFIFO/U799  ( .A(n889), .B(n833), .C(n944), .Q(\u_outFIFO/n969 )
         );
  OAI212 \u_outFIFO/U798  ( .A(n1729), .B(n1190), .C(\u_outFIFO/FIFO[111][3] ), 
        .Q(\u_outFIFO/n968 ) );
  OAI212 \u_outFIFO/U797  ( .A(n1729), .B(n954), .C(\u_outFIFO/n968 ), .Q(
        \u_outFIFO/n1305 ) );
  OAI212 \u_outFIFO/U795  ( .A(n889), .B(n830), .C(n943), .Q(\u_outFIFO/n967 )
         );
  OAI212 \u_outFIFO/U794  ( .A(n1728), .B(n1189), .C(\u_outFIFO/FIFO[111][2] ), 
        .Q(\u_outFIFO/n966 ) );
  OAI212 \u_outFIFO/U793  ( .A(n1728), .B(n959), .C(\u_outFIFO/n966 ), .Q(
        \u_outFIFO/n1304 ) );
  OAI212 \u_outFIFO/U791  ( .A(\u_outFIFO/n396 ), .B(n827), .C(n943), .Q(
        \u_outFIFO/n965 ) );
  OAI212 \u_outFIFO/U790  ( .A(n1727), .B(n1187), .C(\u_outFIFO/FIFO[111][1] ), 
        .Q(\u_outFIFO/n964 ) );
  OAI212 \u_outFIFO/U789  ( .A(n1727), .B(n958), .C(\u_outFIFO/n964 ), .Q(
        \u_outFIFO/n1303 ) );
  OAI212 \u_outFIFO/U787  ( .A(\u_outFIFO/n396 ), .B(n825), .C(n943), .Q(
        \u_outFIFO/n962 ) );
  OAI212 \u_outFIFO/U786  ( .A(n1726), .B(n1186), .C(\u_outFIFO/FIFO[111][0] ), 
        .Q(\u_outFIFO/n961 ) );
  OAI212 \u_outFIFO/U785  ( .A(n1726), .B(n957), .C(\u_outFIFO/n961 ), .Q(
        \u_outFIFO/n1302 ) );
  OAI212 \u_outFIFO/U784  ( .A(n877), .B(n833), .C(n943), .Q(\u_outFIFO/n960 )
         );
  OAI212 \u_outFIFO/U783  ( .A(n1725), .B(n1185), .C(\u_outFIFO/FIFO[110][3] ), 
        .Q(\u_outFIFO/n959 ) );
  OAI212 \u_outFIFO/U782  ( .A(n1725), .B(n956), .C(\u_outFIFO/n959 ), .Q(
        \u_outFIFO/n1301 ) );
  OAI212 \u_outFIFO/U781  ( .A(n877), .B(n830), .C(n943), .Q(\u_outFIFO/n958 )
         );
  OAI212 \u_outFIFO/U780  ( .A(n1724), .B(n1190), .C(\u_outFIFO/FIFO[110][2] ), 
        .Q(\u_outFIFO/n957 ) );
  OAI212 \u_outFIFO/U779  ( .A(n1724), .B(n955), .C(\u_outFIFO/n957 ), .Q(
        \u_outFIFO/n1300 ) );
  OAI212 \u_outFIFO/U778  ( .A(\u_outFIFO/n391 ), .B(n827), .C(n943), .Q(
        \u_outFIFO/n956 ) );
  OAI212 \u_outFIFO/U777  ( .A(n1723), .B(n1187), .C(\u_outFIFO/FIFO[110][1] ), 
        .Q(\u_outFIFO/n955 ) );
  OAI212 \u_outFIFO/U776  ( .A(n1723), .B(n954), .C(\u_outFIFO/n955 ), .Q(
        \u_outFIFO/n1299 ) );
  OAI212 \u_outFIFO/U775  ( .A(\u_outFIFO/n391 ), .B(n825), .C(n943), .Q(
        \u_outFIFO/n954 ) );
  OAI212 \u_outFIFO/U774  ( .A(n1722), .B(n1186), .C(\u_outFIFO/FIFO[110][0] ), 
        .Q(\u_outFIFO/n953 ) );
  OAI212 \u_outFIFO/U773  ( .A(n1722), .B(n1795), .C(\u_outFIFO/n953 ), .Q(
        \u_outFIFO/n1298 ) );
  OAI212 \u_outFIFO/U772  ( .A(n875), .B(n833), .C(n943), .Q(\u_outFIFO/n952 )
         );
  OAI212 \u_outFIFO/U771  ( .A(n1721), .B(n1185), .C(\u_outFIFO/FIFO[109][3] ), 
        .Q(\u_outFIFO/n951 ) );
  OAI212 \u_outFIFO/U770  ( .A(n1721), .B(n961), .C(\u_outFIFO/n951 ), .Q(
        \u_outFIFO/n1297 ) );
  OAI212 \u_outFIFO/U769  ( .A(n875), .B(n830), .C(n942), .Q(\u_outFIFO/n950 )
         );
  OAI212 \u_outFIFO/U768  ( .A(n1720), .B(n1186), .C(\u_outFIFO/FIFO[109][2] ), 
        .Q(\u_outFIFO/n949 ) );
  OAI212 \u_outFIFO/U767  ( .A(n1720), .B(n960), .C(\u_outFIFO/n949 ), .Q(
        \u_outFIFO/n1296 ) );
  OAI212 \u_outFIFO/U766  ( .A(\u_outFIFO/n386 ), .B(n827), .C(n942), .Q(
        \u_outFIFO/n948 ) );
  OAI212 \u_outFIFO/U765  ( .A(n1719), .B(n1185), .C(\u_outFIFO/FIFO[109][1] ), 
        .Q(\u_outFIFO/n947 ) );
  OAI212 \u_outFIFO/U764  ( .A(n1719), .B(n959), .C(\u_outFIFO/n947 ), .Q(
        \u_outFIFO/n1295 ) );
  OAI212 \u_outFIFO/U763  ( .A(\u_outFIFO/n386 ), .B(n825), .C(n942), .Q(
        \u_outFIFO/n946 ) );
  OAI212 \u_outFIFO/U762  ( .A(n1718), .B(n1186), .C(\u_outFIFO/FIFO[109][0] ), 
        .Q(\u_outFIFO/n945 ) );
  OAI212 \u_outFIFO/U761  ( .A(n1718), .B(n958), .C(\u_outFIFO/n945 ), .Q(
        \u_outFIFO/n1294 ) );
  OAI212 \u_outFIFO/U760  ( .A(\u_outFIFO/n381 ), .B(n833), .C(n942), .Q(
        \u_outFIFO/n944 ) );
  OAI212 \u_outFIFO/U759  ( .A(n1717), .B(n1185), .C(\u_outFIFO/FIFO[108][3] ), 
        .Q(\u_outFIFO/n943 ) );
  OAI212 \u_outFIFO/U758  ( .A(n1717), .B(n957), .C(\u_outFIFO/n943 ), .Q(
        \u_outFIFO/n1293 ) );
  OAI212 \u_outFIFO/U757  ( .A(\u_outFIFO/n381 ), .B(n830), .C(n942), .Q(
        \u_outFIFO/n942 ) );
  OAI212 \u_outFIFO/U756  ( .A(n1716), .B(n1186), .C(\u_outFIFO/FIFO[108][2] ), 
        .Q(\u_outFIFO/n941 ) );
  OAI212 \u_outFIFO/U755  ( .A(n1716), .B(n956), .C(\u_outFIFO/n941 ), .Q(
        \u_outFIFO/n1292 ) );
  OAI212 \u_outFIFO/U754  ( .A(n873), .B(n827), .C(n942), .Q(\u_outFIFO/n940 )
         );
  OAI212 \u_outFIFO/U753  ( .A(n1715), .B(n1185), .C(\u_outFIFO/FIFO[108][1] ), 
        .Q(\u_outFIFO/n939 ) );
  OAI212 \u_outFIFO/U752  ( .A(n1715), .B(n952), .C(\u_outFIFO/n939 ), .Q(
        \u_outFIFO/n1291 ) );
  OAI212 \u_outFIFO/U751  ( .A(n873), .B(n825), .C(n942), .Q(\u_outFIFO/n938 )
         );
  OAI212 \u_outFIFO/U750  ( .A(n1714), .B(n1190), .C(\u_outFIFO/FIFO[108][0] ), 
        .Q(\u_outFIFO/n937 ) );
  OAI212 \u_outFIFO/U749  ( .A(n1714), .B(n952), .C(\u_outFIFO/n937 ), .Q(
        \u_outFIFO/n1290 ) );
  OAI212 \u_outFIFO/U748  ( .A(n869), .B(n833), .C(n942), .Q(\u_outFIFO/n936 )
         );
  OAI212 \u_outFIFO/U747  ( .A(n1713), .B(n1190), .C(\u_outFIFO/FIFO[107][3] ), 
        .Q(\u_outFIFO/n935 ) );
  OAI212 \u_outFIFO/U746  ( .A(n1713), .B(n952), .C(\u_outFIFO/n935 ), .Q(
        \u_outFIFO/n1289 ) );
  OAI212 \u_outFIFO/U745  ( .A(n869), .B(n830), .C(n941), .Q(\u_outFIFO/n934 )
         );
  OAI212 \u_outFIFO/U744  ( .A(n1712), .B(n1190), .C(\u_outFIFO/FIFO[107][2] ), 
        .Q(\u_outFIFO/n933 ) );
  OAI212 \u_outFIFO/U743  ( .A(n1712), .B(n952), .C(\u_outFIFO/n933 ), .Q(
        \u_outFIFO/n1288 ) );
  OAI212 \u_outFIFO/U742  ( .A(n871), .B(n827), .C(n941), .Q(\u_outFIFO/n932 )
         );
  OAI212 \u_outFIFO/U741  ( .A(n1711), .B(n1190), .C(\u_outFIFO/FIFO[107][1] ), 
        .Q(\u_outFIFO/n931 ) );
  OAI212 \u_outFIFO/U740  ( .A(n1711), .B(n952), .C(\u_outFIFO/n931 ), .Q(
        \u_outFIFO/n1287 ) );
  OAI212 \u_outFIFO/U739  ( .A(n870), .B(n825), .C(n941), .Q(\u_outFIFO/n930 )
         );
  OAI212 \u_outFIFO/U738  ( .A(n1710), .B(n1190), .C(\u_outFIFO/FIFO[107][0] ), 
        .Q(\u_outFIFO/n929 ) );
  OAI212 \u_outFIFO/U737  ( .A(n1710), .B(n952), .C(\u_outFIFO/n929 ), .Q(
        \u_outFIFO/n1286 ) );
  OAI212 \u_outFIFO/U736  ( .A(n866), .B(n833), .C(n941), .Q(\u_outFIFO/n928 )
         );
  OAI212 \u_outFIFO/U735  ( .A(n1709), .B(n1190), .C(\u_outFIFO/FIFO[106][3] ), 
        .Q(\u_outFIFO/n927 ) );
  OAI212 \u_outFIFO/U734  ( .A(n1709), .B(n952), .C(\u_outFIFO/n927 ), .Q(
        \u_outFIFO/n1285 ) );
  OAI212 \u_outFIFO/U733  ( .A(n866), .B(n830), .C(n941), .Q(\u_outFIFO/n926 )
         );
  OAI212 \u_outFIFO/U732  ( .A(n1708), .B(n1190), .C(\u_outFIFO/FIFO[106][2] ), 
        .Q(\u_outFIFO/n925 ) );
  OAI212 \u_outFIFO/U731  ( .A(n1708), .B(n952), .C(\u_outFIFO/n925 ), .Q(
        \u_outFIFO/n1284 ) );
  OAI212 \u_outFIFO/U730  ( .A(n868), .B(n827), .C(n941), .Q(\u_outFIFO/n924 )
         );
  OAI212 \u_outFIFO/U729  ( .A(n1707), .B(n1190), .C(\u_outFIFO/FIFO[106][1] ), 
        .Q(\u_outFIFO/n923 ) );
  OAI212 \u_outFIFO/U728  ( .A(n1707), .B(n952), .C(\u_outFIFO/n923 ), .Q(
        \u_outFIFO/n1283 ) );
  OAI212 \u_outFIFO/U727  ( .A(n867), .B(n825), .C(n941), .Q(\u_outFIFO/n922 )
         );
  OAI212 \u_outFIFO/U726  ( .A(n1706), .B(n1190), .C(\u_outFIFO/FIFO[106][0] ), 
        .Q(\u_outFIFO/n921 ) );
  OAI212 \u_outFIFO/U725  ( .A(n1706), .B(n952), .C(\u_outFIFO/n921 ), .Q(
        \u_outFIFO/n1282 ) );
  OAI212 \u_outFIFO/U724  ( .A(n863), .B(n835), .C(n941), .Q(\u_outFIFO/n920 )
         );
  OAI212 \u_outFIFO/U723  ( .A(n1705), .B(n1190), .C(\u_outFIFO/FIFO[105][3] ), 
        .Q(\u_outFIFO/n919 ) );
  OAI212 \u_outFIFO/U722  ( .A(n1705), .B(n952), .C(\u_outFIFO/n919 ), .Q(
        \u_outFIFO/n1281 ) );
  OAI212 \u_outFIFO/U721  ( .A(n863), .B(n832), .C(n940), .Q(\u_outFIFO/n918 )
         );
  OAI212 \u_outFIFO/U720  ( .A(n1704), .B(n1190), .C(\u_outFIFO/FIFO[105][2] ), 
        .Q(\u_outFIFO/n917 ) );
  OAI212 \u_outFIFO/U719  ( .A(n1704), .B(n952), .C(\u_outFIFO/n917 ), .Q(
        \u_outFIFO/n1280 ) );
  OAI212 \u_outFIFO/U718  ( .A(n865), .B(n829), .C(n940), .Q(\u_outFIFO/n916 )
         );
  OAI212 \u_outFIFO/U717  ( .A(n1703), .B(n1190), .C(\u_outFIFO/FIFO[105][1] ), 
        .Q(\u_outFIFO/n915 ) );
  OAI212 \u_outFIFO/U716  ( .A(n1703), .B(n952), .C(\u_outFIFO/n915 ), .Q(
        \u_outFIFO/n1279 ) );
  OAI212 \u_outFIFO/U715  ( .A(n864), .B(n825), .C(n940), .Q(\u_outFIFO/n914 )
         );
  OAI212 \u_outFIFO/U714  ( .A(n1702), .B(n1190), .C(\u_outFIFO/FIFO[105][0] ), 
        .Q(\u_outFIFO/n913 ) );
  OAI212 \u_outFIFO/U713  ( .A(n1702), .B(n953), .C(\u_outFIFO/n913 ), .Q(
        \u_outFIFO/n1278 ) );
  OAI212 \u_outFIFO/U712  ( .A(n860), .B(n834), .C(n940), .Q(\u_outFIFO/n912 )
         );
  OAI212 \u_outFIFO/U711  ( .A(n1701), .B(n1190), .C(\u_outFIFO/FIFO[104][3] ), 
        .Q(\u_outFIFO/n911 ) );
  OAI212 \u_outFIFO/U710  ( .A(n1701), .B(n953), .C(\u_outFIFO/n911 ), .Q(
        \u_outFIFO/n1277 ) );
  OAI212 \u_outFIFO/U709  ( .A(n860), .B(n831), .C(n940), .Q(\u_outFIFO/n910 )
         );
  OAI212 \u_outFIFO/U708  ( .A(n1700), .B(n1190), .C(\u_outFIFO/FIFO[104][2] ), 
        .Q(\u_outFIFO/n909 ) );
  OAI212 \u_outFIFO/U707  ( .A(n1700), .B(n953), .C(\u_outFIFO/n909 ), .Q(
        \u_outFIFO/n1276 ) );
  OAI212 \u_outFIFO/U706  ( .A(n862), .B(n828), .C(n940), .Q(\u_outFIFO/n908 )
         );
  OAI212 \u_outFIFO/U705  ( .A(n1699), .B(n1190), .C(\u_outFIFO/FIFO[104][1] ), 
        .Q(\u_outFIFO/n907 ) );
  OAI212 \u_outFIFO/U704  ( .A(n1699), .B(n953), .C(\u_outFIFO/n907 ), .Q(
        \u_outFIFO/n1275 ) );
  OAI212 \u_outFIFO/U703  ( .A(n861), .B(n825), .C(n940), .Q(\u_outFIFO/n906 )
         );
  OAI212 \u_outFIFO/U702  ( .A(n1698), .B(n1190), .C(\u_outFIFO/FIFO[104][0] ), 
        .Q(\u_outFIFO/n905 ) );
  OAI212 \u_outFIFO/U701  ( .A(n1698), .B(n953), .C(\u_outFIFO/n905 ), .Q(
        \u_outFIFO/n1274 ) );
  OAI212 \u_outFIFO/U700  ( .A(n857), .B(n835), .C(n940), .Q(\u_outFIFO/n904 )
         );
  OAI212 \u_outFIFO/U699  ( .A(n1697), .B(n1188), .C(\u_outFIFO/FIFO[103][3] ), 
        .Q(\u_outFIFO/n903 ) );
  OAI212 \u_outFIFO/U698  ( .A(n1697), .B(n953), .C(\u_outFIFO/n903 ), .Q(
        \u_outFIFO/n1273 ) );
  OAI212 \u_outFIFO/U697  ( .A(n857), .B(n832), .C(n939), .Q(\u_outFIFO/n902 )
         );
  OAI212 \u_outFIFO/U696  ( .A(n1696), .B(n1188), .C(\u_outFIFO/FIFO[103][2] ), 
        .Q(\u_outFIFO/n901 ) );
  OAI212 \u_outFIFO/U695  ( .A(n1696), .B(n953), .C(\u_outFIFO/n901 ), .Q(
        \u_outFIFO/n1272 ) );
  OAI212 \u_outFIFO/U694  ( .A(n859), .B(n829), .C(n939), .Q(\u_outFIFO/n900 )
         );
  OAI212 \u_outFIFO/U693  ( .A(n1695), .B(n1190), .C(\u_outFIFO/FIFO[103][1] ), 
        .Q(\u_outFIFO/n899 ) );
  OAI212 \u_outFIFO/U692  ( .A(n1695), .B(n953), .C(\u_outFIFO/n899 ), .Q(
        \u_outFIFO/n1271 ) );
  OAI212 \u_outFIFO/U691  ( .A(n858), .B(n826), .C(n939), .Q(\u_outFIFO/n898 )
         );
  OAI212 \u_outFIFO/U690  ( .A(n1694), .B(n1189), .C(\u_outFIFO/FIFO[103][0] ), 
        .Q(\u_outFIFO/n897 ) );
  OAI212 \u_outFIFO/U689  ( .A(n1694), .B(n953), .C(\u_outFIFO/n897 ), .Q(
        \u_outFIFO/n1270 ) );
  OAI212 \u_outFIFO/U688  ( .A(n854), .B(n834), .C(n939), .Q(\u_outFIFO/n896 )
         );
  OAI212 \u_outFIFO/U687  ( .A(n1693), .B(n1188), .C(\u_outFIFO/FIFO[102][3] ), 
        .Q(\u_outFIFO/n895 ) );
  OAI212 \u_outFIFO/U686  ( .A(n1693), .B(n953), .C(\u_outFIFO/n895 ), .Q(
        \u_outFIFO/n1269 ) );
  OAI212 \u_outFIFO/U685  ( .A(n854), .B(n831), .C(n939), .Q(\u_outFIFO/n894 )
         );
  OAI212 \u_outFIFO/U684  ( .A(n1692), .B(n1186), .C(\u_outFIFO/FIFO[102][2] ), 
        .Q(\u_outFIFO/n893 ) );
  OAI212 \u_outFIFO/U683  ( .A(n1692), .B(n953), .C(\u_outFIFO/n893 ), .Q(
        \u_outFIFO/n1268 ) );
  OAI212 \u_outFIFO/U682  ( .A(n856), .B(n828), .C(n939), .Q(\u_outFIFO/n892 )
         );
  OAI212 \u_outFIFO/U681  ( .A(n1691), .B(n1185), .C(\u_outFIFO/FIFO[102][1] ), 
        .Q(\u_outFIFO/n891 ) );
  OAI212 \u_outFIFO/U680  ( .A(n1691), .B(n953), .C(\u_outFIFO/n891 ), .Q(
        \u_outFIFO/n1267 ) );
  OAI212 \u_outFIFO/U679  ( .A(n855), .B(n826), .C(n939), .Q(\u_outFIFO/n890 )
         );
  OAI212 \u_outFIFO/U678  ( .A(n1690), .B(n1190), .C(\u_outFIFO/FIFO[102][0] ), 
        .Q(\u_outFIFO/n889 ) );
  OAI212 \u_outFIFO/U677  ( .A(n1690), .B(n953), .C(\u_outFIFO/n889 ), .Q(
        \u_outFIFO/n1266 ) );
  OAI212 \u_outFIFO/U676  ( .A(n851), .B(n835), .C(n939), .Q(\u_outFIFO/n888 )
         );
  OAI212 \u_outFIFO/U675  ( .A(n1689), .B(n1190), .C(\u_outFIFO/FIFO[101][3] ), 
        .Q(\u_outFIFO/n887 ) );
  OAI212 \u_outFIFO/U674  ( .A(n1689), .B(n954), .C(\u_outFIFO/n887 ), .Q(
        \u_outFIFO/n1265 ) );
  OAI212 \u_outFIFO/U673  ( .A(n851), .B(n832), .C(n938), .Q(\u_outFIFO/n886 )
         );
  OAI212 \u_outFIFO/U672  ( .A(n1688), .B(n1190), .C(\u_outFIFO/FIFO[101][2] ), 
        .Q(\u_outFIFO/n885 ) );
  OAI212 \u_outFIFO/U671  ( .A(n1688), .B(n954), .C(\u_outFIFO/n885 ), .Q(
        \u_outFIFO/n1264 ) );
  OAI212 \u_outFIFO/U670  ( .A(n853), .B(n829), .C(n938), .Q(\u_outFIFO/n884 )
         );
  OAI212 \u_outFIFO/U669  ( .A(n1687), .B(n1187), .C(\u_outFIFO/FIFO[101][1] ), 
        .Q(\u_outFIFO/n883 ) );
  OAI212 \u_outFIFO/U668  ( .A(n1687), .B(n954), .C(\u_outFIFO/n883 ), .Q(
        \u_outFIFO/n1263 ) );
  OAI212 \u_outFIFO/U667  ( .A(n852), .B(n826), .C(n938), .Q(\u_outFIFO/n882 )
         );
  OAI212 \u_outFIFO/U666  ( .A(n1686), .B(n1184), .C(\u_outFIFO/FIFO[101][0] ), 
        .Q(\u_outFIFO/n881 ) );
  OAI212 \u_outFIFO/U665  ( .A(n1686), .B(n954), .C(\u_outFIFO/n881 ), .Q(
        \u_outFIFO/n1262 ) );
  OAI212 \u_outFIFO/U664  ( .A(n848), .B(n834), .C(n938), .Q(\u_outFIFO/n880 )
         );
  OAI212 \u_outFIFO/U663  ( .A(n1685), .B(n1184), .C(\u_outFIFO/FIFO[100][3] ), 
        .Q(\u_outFIFO/n879 ) );
  OAI212 \u_outFIFO/U662  ( .A(n1685), .B(n954), .C(\u_outFIFO/n879 ), .Q(
        \u_outFIFO/n1261 ) );
  OAI212 \u_outFIFO/U661  ( .A(n848), .B(n831), .C(n938), .Q(\u_outFIFO/n878 )
         );
  OAI212 \u_outFIFO/U660  ( .A(n1684), .B(n1184), .C(\u_outFIFO/FIFO[100][2] ), 
        .Q(\u_outFIFO/n877 ) );
  OAI212 \u_outFIFO/U659  ( .A(n1684), .B(n954), .C(\u_outFIFO/n877 ), .Q(
        \u_outFIFO/n1260 ) );
  OAI212 \u_outFIFO/U658  ( .A(n850), .B(n828), .C(n938), .Q(\u_outFIFO/n876 )
         );
  OAI212 \u_outFIFO/U657  ( .A(n1683), .B(n1184), .C(\u_outFIFO/FIFO[100][1] ), 
        .Q(\u_outFIFO/n875 ) );
  OAI212 \u_outFIFO/U656  ( .A(n1683), .B(n954), .C(\u_outFIFO/n875 ), .Q(
        \u_outFIFO/n1259 ) );
  OAI212 \u_outFIFO/U655  ( .A(n849), .B(n826), .C(n938), .Q(\u_outFIFO/n874 )
         );
  OAI212 \u_outFIFO/U654  ( .A(n1682), .B(n1184), .C(\u_outFIFO/FIFO[100][0] ), 
        .Q(\u_outFIFO/n873 ) );
  OAI212 \u_outFIFO/U653  ( .A(n1682), .B(n954), .C(\u_outFIFO/n873 ), .Q(
        \u_outFIFO/n1258 ) );
  OAI212 \u_outFIFO/U652  ( .A(n844), .B(n835), .C(n938), .Q(\u_outFIFO/n872 )
         );
  OAI212 \u_outFIFO/U651  ( .A(n1681), .B(n1184), .C(\u_outFIFO/FIFO[99][3] ), 
        .Q(\u_outFIFO/n871 ) );
  OAI212 \u_outFIFO/U650  ( .A(n1681), .B(n954), .C(\u_outFIFO/n871 ), .Q(
        \u_outFIFO/n1257 ) );
  OAI212 \u_outFIFO/U649  ( .A(n845), .B(n832), .C(n937), .Q(\u_outFIFO/n870 )
         );
  OAI212 \u_outFIFO/U648  ( .A(n1680), .B(n1184), .C(\u_outFIFO/FIFO[99][2] ), 
        .Q(\u_outFIFO/n869 ) );
  OAI212 \u_outFIFO/U647  ( .A(n1680), .B(n954), .C(\u_outFIFO/n869 ), .Q(
        \u_outFIFO/n1256 ) );
  OAI212 \u_outFIFO/U646  ( .A(n846), .B(n829), .C(n937), .Q(\u_outFIFO/n868 )
         );
  OAI212 \u_outFIFO/U645  ( .A(n1679), .B(n1184), .C(\u_outFIFO/FIFO[99][1] ), 
        .Q(\u_outFIFO/n867 ) );
  OAI212 \u_outFIFO/U644  ( .A(n1679), .B(n954), .C(\u_outFIFO/n867 ), .Q(
        \u_outFIFO/n1255 ) );
  OAI212 \u_outFIFO/U643  ( .A(n847), .B(n826), .C(n937), .Q(\u_outFIFO/n866 )
         );
  OAI212 \u_outFIFO/U642  ( .A(n1678), .B(n1184), .C(\u_outFIFO/FIFO[99][0] ), 
        .Q(\u_outFIFO/n865 ) );
  OAI212 \u_outFIFO/U641  ( .A(n1678), .B(n954), .C(\u_outFIFO/n865 ), .Q(
        \u_outFIFO/n1254 ) );
  OAI212 \u_outFIFO/U640  ( .A(\u_outFIFO/n331 ), .B(n834), .C(n937), .Q(
        \u_outFIFO/n864 ) );
  OAI212 \u_outFIFO/U639  ( .A(n1677), .B(n1184), .C(\u_outFIFO/FIFO[98][3] ), 
        .Q(\u_outFIFO/n863 ) );
  OAI212 \u_outFIFO/U638  ( .A(n1677), .B(n954), .C(\u_outFIFO/n863 ), .Q(
        \u_outFIFO/n1253 ) );
  OAI212 \u_outFIFO/U637  ( .A(\u_outFIFO/n331 ), .B(n831), .C(n937), .Q(
        \u_outFIFO/n862 ) );
  OAI212 \u_outFIFO/U636  ( .A(n1676), .B(n1184), .C(\u_outFIFO/FIFO[98][2] ), 
        .Q(\u_outFIFO/n861 ) );
  OAI212 \u_outFIFO/U635  ( .A(n1676), .B(n955), .C(\u_outFIFO/n861 ), .Q(
        \u_outFIFO/n1252 ) );
  OAI212 \u_outFIFO/U634  ( .A(n842), .B(n828), .C(n937), .Q(\u_outFIFO/n860 )
         );
  OAI212 \u_outFIFO/U633  ( .A(n1675), .B(n1185), .C(\u_outFIFO/FIFO[98][1] ), 
        .Q(\u_outFIFO/n859 ) );
  OAI212 \u_outFIFO/U632  ( .A(n1675), .B(n955), .C(\u_outFIFO/n859 ), .Q(
        \u_outFIFO/n1251 ) );
  OAI212 \u_outFIFO/U631  ( .A(\u_outFIFO/n331 ), .B(n826), .C(n937), .Q(
        \u_outFIFO/n858 ) );
  OAI212 \u_outFIFO/U630  ( .A(n1674), .B(n1185), .C(\u_outFIFO/FIFO[98][0] ), 
        .Q(\u_outFIFO/n857 ) );
  OAI212 \u_outFIFO/U629  ( .A(n1674), .B(n955), .C(\u_outFIFO/n857 ), .Q(
        \u_outFIFO/n1250 ) );
  OAI212 \u_outFIFO/U628  ( .A(n838), .B(n835), .C(n937), .Q(\u_outFIFO/n856 )
         );
  OAI212 \u_outFIFO/U627  ( .A(n1673), .B(n1185), .C(\u_outFIFO/FIFO[97][3] ), 
        .Q(\u_outFIFO/n855 ) );
  OAI212 \u_outFIFO/U626  ( .A(n1673), .B(n955), .C(\u_outFIFO/n855 ), .Q(
        \u_outFIFO/n1249 ) );
  OAI212 \u_outFIFO/U625  ( .A(n838), .B(n832), .C(n936), .Q(\u_outFIFO/n854 )
         );
  OAI212 \u_outFIFO/U624  ( .A(n1672), .B(n1185), .C(\u_outFIFO/FIFO[97][2] ), 
        .Q(\u_outFIFO/n853 ) );
  OAI212 \u_outFIFO/U623  ( .A(n1672), .B(n955), .C(\u_outFIFO/n853 ), .Q(
        \u_outFIFO/n1248 ) );
  OAI212 \u_outFIFO/U622  ( .A(n840), .B(n829), .C(n936), .Q(\u_outFIFO/n852 )
         );
  OAI212 \u_outFIFO/U621  ( .A(n1671), .B(n1185), .C(\u_outFIFO/FIFO[97][1] ), 
        .Q(\u_outFIFO/n851 ) );
  OAI212 \u_outFIFO/U620  ( .A(n1671), .B(n955), .C(\u_outFIFO/n851 ), .Q(
        \u_outFIFO/n1247 ) );
  OAI212 \u_outFIFO/U619  ( .A(n839), .B(n826), .C(n936), .Q(\u_outFIFO/n850 )
         );
  OAI212 \u_outFIFO/U618  ( .A(n1670), .B(n1185), .C(\u_outFIFO/FIFO[97][0] ), 
        .Q(\u_outFIFO/n849 ) );
  OAI212 \u_outFIFO/U617  ( .A(n1670), .B(n955), .C(\u_outFIFO/n849 ), .Q(
        \u_outFIFO/n1246 ) );
  OAI212 \u_outFIFO/U616  ( .A(\u_outFIFO/n317 ), .B(n834), .C(n936), .Q(
        \u_outFIFO/n847 ) );
  OAI212 \u_outFIFO/U615  ( .A(n1669), .B(n1185), .C(\u_outFIFO/FIFO[96][3] ), 
        .Q(\u_outFIFO/n846 ) );
  OAI212 \u_outFIFO/U614  ( .A(n1669), .B(n955), .C(\u_outFIFO/n846 ), .Q(
        \u_outFIFO/n1245 ) );
  OAI212 \u_outFIFO/U613  ( .A(\u_outFIFO/n317 ), .B(n831), .C(n936), .Q(
        \u_outFIFO/n844 ) );
  OAI212 \u_outFIFO/U612  ( .A(n1668), .B(n1185), .C(\u_outFIFO/FIFO[96][2] ), 
        .Q(\u_outFIFO/n843 ) );
  OAI212 \u_outFIFO/U611  ( .A(n1668), .B(n955), .C(\u_outFIFO/n843 ), .Q(
        \u_outFIFO/n1244 ) );
  OAI212 \u_outFIFO/U610  ( .A(n837), .B(n828), .C(n936), .Q(\u_outFIFO/n841 )
         );
  OAI212 \u_outFIFO/U609  ( .A(n1667), .B(n1185), .C(\u_outFIFO/FIFO[96][1] ), 
        .Q(\u_outFIFO/n840 ) );
  OAI212 \u_outFIFO/U608  ( .A(n1667), .B(n955), .C(\u_outFIFO/n840 ), .Q(
        \u_outFIFO/n1243 ) );
  OAI212 \u_outFIFO/U607  ( .A(n837), .B(n826), .C(n936), .Q(\u_outFIFO/n838 )
         );
  OAI212 \u_outFIFO/U606  ( .A(n1666), .B(n1185), .C(\u_outFIFO/FIFO[96][0] ), 
        .Q(\u_outFIFO/n837 ) );
  OAI212 \u_outFIFO/U605  ( .A(n1666), .B(n955), .C(\u_outFIFO/n837 ), .Q(
        \u_outFIFO/n1242 ) );
  OAI212 \u_outFIFO/U602  ( .A(\u_outFIFO/n396 ), .B(n822), .C(n936), .Q(
        \u_outFIFO/n836 ) );
  OAI212 \u_outFIFO/U601  ( .A(n1665), .B(n1185), .C(\u_outFIFO/FIFO[95][3] ), 
        .Q(\u_outFIFO/n835 ) );
  OAI212 \u_outFIFO/U600  ( .A(n1665), .B(n955), .C(\u_outFIFO/n835 ), .Q(
        \u_outFIFO/n1241 ) );
  OAI212 \u_outFIFO/U598  ( .A(n889), .B(n819), .C(n935), .Q(\u_outFIFO/n834 )
         );
  OAI212 \u_outFIFO/U597  ( .A(n1664), .B(n1185), .C(\u_outFIFO/FIFO[95][2] ), 
        .Q(\u_outFIFO/n833 ) );
  OAI212 \u_outFIFO/U596  ( .A(n1664), .B(n955), .C(\u_outFIFO/n833 ), .Q(
        \u_outFIFO/n1240 ) );
  OAI212 \u_outFIFO/U594  ( .A(n889), .B(n816), .C(n935), .Q(\u_outFIFO/n832 )
         );
  OAI212 \u_outFIFO/U593  ( .A(n1663), .B(n1185), .C(\u_outFIFO/FIFO[95][1] ), 
        .Q(\u_outFIFO/n831 ) );
  OAI212 \u_outFIFO/U592  ( .A(n1663), .B(n956), .C(\u_outFIFO/n831 ), .Q(
        \u_outFIFO/n1239 ) );
  OAI212 \u_outFIFO/U590  ( .A(n889), .B(n814), .C(n935), .Q(\u_outFIFO/n829 )
         );
  OAI212 \u_outFIFO/U589  ( .A(n1662), .B(n1185), .C(\u_outFIFO/FIFO[95][0] ), 
        .Q(\u_outFIFO/n828 ) );
  OAI212 \u_outFIFO/U588  ( .A(n1662), .B(n956), .C(\u_outFIFO/n828 ), .Q(
        \u_outFIFO/n1238 ) );
  OAI212 \u_outFIFO/U587  ( .A(\u_outFIFO/n391 ), .B(n822), .C(n935), .Q(
        \u_outFIFO/n827 ) );
  OAI212 \u_outFIFO/U586  ( .A(n1661), .B(n1185), .C(\u_outFIFO/FIFO[94][3] ), 
        .Q(\u_outFIFO/n826 ) );
  OAI212 \u_outFIFO/U585  ( .A(n1661), .B(n956), .C(\u_outFIFO/n826 ), .Q(
        \u_outFIFO/n1237 ) );
  OAI212 \u_outFIFO/U584  ( .A(n877), .B(n819), .C(n935), .Q(\u_outFIFO/n825 )
         );
  OAI212 \u_outFIFO/U583  ( .A(n1660), .B(n1185), .C(\u_outFIFO/FIFO[94][2] ), 
        .Q(\u_outFIFO/n824 ) );
  OAI212 \u_outFIFO/U582  ( .A(n1660), .B(n956), .C(\u_outFIFO/n824 ), .Q(
        \u_outFIFO/n1236 ) );
  OAI212 \u_outFIFO/U581  ( .A(n877), .B(n816), .C(n935), .Q(\u_outFIFO/n823 )
         );
  OAI212 \u_outFIFO/U580  ( .A(n1659), .B(n1185), .C(\u_outFIFO/FIFO[94][1] ), 
        .Q(\u_outFIFO/n822 ) );
  OAI212 \u_outFIFO/U579  ( .A(n1659), .B(n956), .C(\u_outFIFO/n822 ), .Q(
        \u_outFIFO/n1235 ) );
  OAI212 \u_outFIFO/U578  ( .A(n877), .B(n814), .C(n935), .Q(\u_outFIFO/n821 )
         );
  OAI212 \u_outFIFO/U577  ( .A(n1658), .B(n1186), .C(\u_outFIFO/FIFO[94][0] ), 
        .Q(\u_outFIFO/n820 ) );
  OAI212 \u_outFIFO/U576  ( .A(n1658), .B(n956), .C(\u_outFIFO/n820 ), .Q(
        \u_outFIFO/n1234 ) );
  OAI212 \u_outFIFO/U575  ( .A(\u_outFIFO/n386 ), .B(n822), .C(n935), .Q(
        \u_outFIFO/n819 ) );
  OAI212 \u_outFIFO/U574  ( .A(n1657), .B(n1186), .C(\u_outFIFO/FIFO[93][3] ), 
        .Q(\u_outFIFO/n818 ) );
  OAI212 \u_outFIFO/U573  ( .A(n1657), .B(n956), .C(\u_outFIFO/n818 ), .Q(
        \u_outFIFO/n1233 ) );
  OAI212 \u_outFIFO/U572  ( .A(n875), .B(n819), .C(n934), .Q(\u_outFIFO/n817 )
         );
  OAI212 \u_outFIFO/U571  ( .A(n1656), .B(n1186), .C(\u_outFIFO/FIFO[93][2] ), 
        .Q(\u_outFIFO/n816 ) );
  OAI212 \u_outFIFO/U570  ( .A(n1656), .B(n956), .C(\u_outFIFO/n816 ), .Q(
        \u_outFIFO/n1232 ) );
  OAI212 \u_outFIFO/U569  ( .A(n875), .B(n816), .C(n934), .Q(\u_outFIFO/n815 )
         );
  OAI212 \u_outFIFO/U568  ( .A(n1655), .B(n1186), .C(\u_outFIFO/FIFO[93][1] ), 
        .Q(\u_outFIFO/n814 ) );
  OAI212 \u_outFIFO/U567  ( .A(n1655), .B(n956), .C(\u_outFIFO/n814 ), .Q(
        \u_outFIFO/n1231 ) );
  OAI212 \u_outFIFO/U566  ( .A(n875), .B(n814), .C(n934), .Q(\u_outFIFO/n813 )
         );
  OAI212 \u_outFIFO/U565  ( .A(n1654), .B(n1186), .C(\u_outFIFO/FIFO[93][0] ), 
        .Q(\u_outFIFO/n812 ) );
  OAI212 \u_outFIFO/U564  ( .A(n1654), .B(n956), .C(\u_outFIFO/n812 ), .Q(
        \u_outFIFO/n1230 ) );
  OAI212 \u_outFIFO/U563  ( .A(\u_outFIFO/n381 ), .B(n822), .C(n934), .Q(
        \u_outFIFO/n811 ) );
  OAI212 \u_outFIFO/U562  ( .A(n1653), .B(n1186), .C(\u_outFIFO/FIFO[92][3] ), 
        .Q(\u_outFIFO/n810 ) );
  OAI212 \u_outFIFO/U561  ( .A(n1653), .B(n956), .C(\u_outFIFO/n810 ), .Q(
        \u_outFIFO/n1229 ) );
  OAI212 \u_outFIFO/U560  ( .A(\u_outFIFO/n381 ), .B(n819), .C(n934), .Q(
        \u_outFIFO/n809 ) );
  OAI212 \u_outFIFO/U559  ( .A(n1652), .B(n1186), .C(\u_outFIFO/FIFO[92][2] ), 
        .Q(\u_outFIFO/n808 ) );
  OAI212 \u_outFIFO/U558  ( .A(n1652), .B(n956), .C(\u_outFIFO/n808 ), .Q(
        \u_outFIFO/n1228 ) );
  OAI212 \u_outFIFO/U557  ( .A(n873), .B(n816), .C(n934), .Q(\u_outFIFO/n807 )
         );
  OAI212 \u_outFIFO/U556  ( .A(n1651), .B(n1186), .C(\u_outFIFO/FIFO[92][1] ), 
        .Q(\u_outFIFO/n806 ) );
  OAI212 \u_outFIFO/U555  ( .A(n1651), .B(n956), .C(\u_outFIFO/n806 ), .Q(
        \u_outFIFO/n1227 ) );
  OAI212 \u_outFIFO/U554  ( .A(\u_outFIFO/n381 ), .B(n814), .C(n934), .Q(
        \u_outFIFO/n805 ) );
  OAI212 \u_outFIFO/U553  ( .A(n1650), .B(n1186), .C(\u_outFIFO/FIFO[92][0] ), 
        .Q(\u_outFIFO/n804 ) );
  OAI212 \u_outFIFO/U552  ( .A(n1650), .B(n957), .C(\u_outFIFO/n804 ), .Q(
        \u_outFIFO/n1226 ) );
  OAI212 \u_outFIFO/U551  ( .A(n871), .B(n822), .C(n934), .Q(\u_outFIFO/n803 )
         );
  OAI212 \u_outFIFO/U550  ( .A(n1649), .B(n1186), .C(\u_outFIFO/FIFO[91][3] ), 
        .Q(\u_outFIFO/n802 ) );
  OAI212 \u_outFIFO/U549  ( .A(n1649), .B(n957), .C(\u_outFIFO/n802 ), .Q(
        \u_outFIFO/n1225 ) );
  OAI212 \u_outFIFO/U548  ( .A(n870), .B(n819), .C(n933), .Q(\u_outFIFO/n801 )
         );
  OAI212 \u_outFIFO/U547  ( .A(n1648), .B(n1186), .C(\u_outFIFO/FIFO[91][2] ), 
        .Q(\u_outFIFO/n800 ) );
  OAI212 \u_outFIFO/U546  ( .A(n1648), .B(n957), .C(\u_outFIFO/n800 ), .Q(
        \u_outFIFO/n1224 ) );
  OAI212 \u_outFIFO/U545  ( .A(n871), .B(n816), .C(n933), .Q(\u_outFIFO/n799 )
         );
  OAI212 \u_outFIFO/U544  ( .A(n1647), .B(n1186), .C(\u_outFIFO/FIFO[91][1] ), 
        .Q(\u_outFIFO/n798 ) );
  OAI212 \u_outFIFO/U543  ( .A(n1647), .B(n957), .C(\u_outFIFO/n798 ), .Q(
        \u_outFIFO/n1223 ) );
  OAI212 \u_outFIFO/U542  ( .A(n870), .B(n814), .C(n933), .Q(\u_outFIFO/n797 )
         );
  OAI212 \u_outFIFO/U541  ( .A(n1646), .B(n1186), .C(\u_outFIFO/FIFO[91][0] ), 
        .Q(\u_outFIFO/n796 ) );
  OAI212 \u_outFIFO/U540  ( .A(n1646), .B(n957), .C(\u_outFIFO/n796 ), .Q(
        \u_outFIFO/n1222 ) );
  OAI212 \u_outFIFO/U539  ( .A(n868), .B(n822), .C(n933), .Q(\u_outFIFO/n795 )
         );
  OAI212 \u_outFIFO/U538  ( .A(n1645), .B(n1186), .C(\u_outFIFO/FIFO[90][3] ), 
        .Q(\u_outFIFO/n794 ) );
  OAI212 \u_outFIFO/U537  ( .A(n1645), .B(n957), .C(\u_outFIFO/n794 ), .Q(
        \u_outFIFO/n1221 ) );
  OAI212 \u_outFIFO/U536  ( .A(n867), .B(n819), .C(n933), .Q(\u_outFIFO/n793 )
         );
  OAI212 \u_outFIFO/U535  ( .A(n1644), .B(n1186), .C(\u_outFIFO/FIFO[90][2] ), 
        .Q(\u_outFIFO/n792 ) );
  OAI212 \u_outFIFO/U534  ( .A(n1644), .B(n957), .C(\u_outFIFO/n792 ), .Q(
        \u_outFIFO/n1220 ) );
  OAI212 \u_outFIFO/U533  ( .A(n868), .B(n816), .C(n933), .Q(\u_outFIFO/n791 )
         );
  OAI212 \u_outFIFO/U532  ( .A(n1643), .B(n1186), .C(\u_outFIFO/FIFO[90][1] ), 
        .Q(\u_outFIFO/n790 ) );
  OAI212 \u_outFIFO/U531  ( .A(n1643), .B(n957), .C(\u_outFIFO/n790 ), .Q(
        \u_outFIFO/n1219 ) );
  OAI212 \u_outFIFO/U530  ( .A(n867), .B(n814), .C(n933), .Q(\u_outFIFO/n789 )
         );
  OAI212 \u_outFIFO/U529  ( .A(n1642), .B(n1186), .C(\u_outFIFO/FIFO[90][0] ), 
        .Q(\u_outFIFO/n788 ) );
  OAI212 \u_outFIFO/U528  ( .A(n1642), .B(n957), .C(\u_outFIFO/n788 ), .Q(
        \u_outFIFO/n1218 ) );
  OAI212 \u_outFIFO/U527  ( .A(n865), .B(n824), .C(n933), .Q(\u_outFIFO/n787 )
         );
  OAI212 \u_outFIFO/U526  ( .A(n1641), .B(n1187), .C(\u_outFIFO/FIFO[89][3] ), 
        .Q(\u_outFIFO/n786 ) );
  OAI212 \u_outFIFO/U525  ( .A(n1641), .B(n957), .C(\u_outFIFO/n786 ), .Q(
        \u_outFIFO/n1217 ) );
  OAI212 \u_outFIFO/U524  ( .A(n864), .B(n821), .C(n932), .Q(\u_outFIFO/n785 )
         );
  OAI212 \u_outFIFO/U523  ( .A(n1640), .B(n1187), .C(\u_outFIFO/FIFO[89][2] ), 
        .Q(\u_outFIFO/n784 ) );
  OAI212 \u_outFIFO/U522  ( .A(n1640), .B(n957), .C(\u_outFIFO/n784 ), .Q(
        \u_outFIFO/n1216 ) );
  OAI212 \u_outFIFO/U521  ( .A(n865), .B(n818), .C(n932), .Q(\u_outFIFO/n783 )
         );
  OAI212 \u_outFIFO/U520  ( .A(n1639), .B(n1187), .C(\u_outFIFO/FIFO[89][1] ), 
        .Q(\u_outFIFO/n782 ) );
  OAI212 \u_outFIFO/U519  ( .A(n1639), .B(n957), .C(\u_outFIFO/n782 ), .Q(
        \u_outFIFO/n1215 ) );
  OAI212 \u_outFIFO/U518  ( .A(n864), .B(n814), .C(n932), .Q(\u_outFIFO/n781 )
         );
  OAI212 \u_outFIFO/U517  ( .A(n1638), .B(n1187), .C(\u_outFIFO/FIFO[89][0] ), 
        .Q(\u_outFIFO/n780 ) );
  OAI212 \u_outFIFO/U516  ( .A(n1638), .B(n957), .C(\u_outFIFO/n780 ), .Q(
        \u_outFIFO/n1214 ) );
  OAI212 \u_outFIFO/U515  ( .A(n862), .B(n823), .C(n932), .Q(\u_outFIFO/n779 )
         );
  OAI212 \u_outFIFO/U514  ( .A(n1637), .B(n1187), .C(\u_outFIFO/FIFO[88][3] ), 
        .Q(\u_outFIFO/n778 ) );
  OAI212 \u_outFIFO/U513  ( .A(n1637), .B(n958), .C(\u_outFIFO/n778 ), .Q(
        \u_outFIFO/n1213 ) );
  OAI212 \u_outFIFO/U512  ( .A(n861), .B(n820), .C(n932), .Q(\u_outFIFO/n777 )
         );
  OAI212 \u_outFIFO/U511  ( .A(n1636), .B(n1187), .C(\u_outFIFO/FIFO[88][2] ), 
        .Q(\u_outFIFO/n776 ) );
  OAI212 \u_outFIFO/U510  ( .A(n1636), .B(n958), .C(\u_outFIFO/n776 ), .Q(
        \u_outFIFO/n1212 ) );
  OAI212 \u_outFIFO/U509  ( .A(n862), .B(n817), .C(n932), .Q(\u_outFIFO/n775 )
         );
  OAI212 \u_outFIFO/U508  ( .A(n1635), .B(n1187), .C(\u_outFIFO/FIFO[88][1] ), 
        .Q(\u_outFIFO/n774 ) );
  OAI212 \u_outFIFO/U507  ( .A(n1635), .B(n958), .C(\u_outFIFO/n774 ), .Q(
        \u_outFIFO/n1211 ) );
  OAI212 \u_outFIFO/U506  ( .A(n861), .B(n814), .C(n932), .Q(\u_outFIFO/n773 )
         );
  OAI212 \u_outFIFO/U505  ( .A(n1634), .B(n1189), .C(\u_outFIFO/FIFO[88][0] ), 
        .Q(\u_outFIFO/n772 ) );
  OAI212 \u_outFIFO/U504  ( .A(n1634), .B(n958), .C(\u_outFIFO/n772 ), .Q(
        \u_outFIFO/n1210 ) );
  OAI212 \u_outFIFO/U503  ( .A(n859), .B(n824), .C(n932), .Q(\u_outFIFO/n771 )
         );
  OAI212 \u_outFIFO/U502  ( .A(n1633), .B(n1187), .C(\u_outFIFO/FIFO[87][3] ), 
        .Q(\u_outFIFO/n770 ) );
  OAI212 \u_outFIFO/U501  ( .A(n1633), .B(n958), .C(\u_outFIFO/n770 ), .Q(
        \u_outFIFO/n1209 ) );
  OAI212 \u_outFIFO/U500  ( .A(n858), .B(n821), .C(n931), .Q(\u_outFIFO/n769 )
         );
  OAI212 \u_outFIFO/U499  ( .A(n1632), .B(n1187), .C(\u_outFIFO/FIFO[87][2] ), 
        .Q(\u_outFIFO/n768 ) );
  OAI212 \u_outFIFO/U498  ( .A(n1632), .B(n958), .C(\u_outFIFO/n768 ), .Q(
        \u_outFIFO/n1208 ) );
  OAI212 \u_outFIFO/U497  ( .A(n859), .B(n818), .C(n931), .Q(\u_outFIFO/n767 )
         );
  OAI212 \u_outFIFO/U496  ( .A(n1631), .B(n1187), .C(\u_outFIFO/FIFO[87][1] ), 
        .Q(\u_outFIFO/n766 ) );
  OAI212 \u_outFIFO/U495  ( .A(n1631), .B(n958), .C(\u_outFIFO/n766 ), .Q(
        \u_outFIFO/n1207 ) );
  OAI212 \u_outFIFO/U494  ( .A(n858), .B(n815), .C(n931), .Q(\u_outFIFO/n765 )
         );
  OAI212 \u_outFIFO/U493  ( .A(n1630), .B(n1187), .C(\u_outFIFO/FIFO[87][0] ), 
        .Q(\u_outFIFO/n764 ) );
  OAI212 \u_outFIFO/U492  ( .A(n1630), .B(n958), .C(\u_outFIFO/n764 ), .Q(
        \u_outFIFO/n1206 ) );
  OAI212 \u_outFIFO/U491  ( .A(n856), .B(n823), .C(n931), .Q(\u_outFIFO/n763 )
         );
  OAI212 \u_outFIFO/U490  ( .A(n1629), .B(n1187), .C(\u_outFIFO/FIFO[86][3] ), 
        .Q(\u_outFIFO/n762 ) );
  OAI212 \u_outFIFO/U489  ( .A(n1629), .B(n958), .C(\u_outFIFO/n762 ), .Q(
        \u_outFIFO/n1205 ) );
  OAI212 \u_outFIFO/U488  ( .A(n855), .B(n820), .C(n931), .Q(\u_outFIFO/n761 )
         );
  OAI212 \u_outFIFO/U487  ( .A(n1628), .B(n1187), .C(\u_outFIFO/FIFO[86][2] ), 
        .Q(\u_outFIFO/n760 ) );
  OAI212 \u_outFIFO/U486  ( .A(n1628), .B(n958), .C(\u_outFIFO/n760 ), .Q(
        \u_outFIFO/n1204 ) );
  OAI212 \u_outFIFO/U485  ( .A(n856), .B(n817), .C(n931), .Q(\u_outFIFO/n759 )
         );
  OAI212 \u_outFIFO/U484  ( .A(n1627), .B(n1187), .C(\u_outFIFO/FIFO[86][1] ), 
        .Q(\u_outFIFO/n758 ) );
  OAI212 \u_outFIFO/U483  ( .A(n1627), .B(n958), .C(\u_outFIFO/n758 ), .Q(
        \u_outFIFO/n1203 ) );
  OAI212 \u_outFIFO/U482  ( .A(n855), .B(n815), .C(n931), .Q(\u_outFIFO/n757 )
         );
  OAI212 \u_outFIFO/U481  ( .A(n1626), .B(n1187), .C(\u_outFIFO/FIFO[86][0] ), 
        .Q(\u_outFIFO/n756 ) );
  OAI212 \u_outFIFO/U480  ( .A(n1626), .B(n958), .C(\u_outFIFO/n756 ), .Q(
        \u_outFIFO/n1202 ) );
  OAI212 \u_outFIFO/U479  ( .A(n853), .B(n824), .C(n931), .Q(\u_outFIFO/n755 )
         );
  OAI212 \u_outFIFO/U478  ( .A(n1625), .B(n1187), .C(\u_outFIFO/FIFO[85][3] ), 
        .Q(\u_outFIFO/n754 ) );
  OAI212 \u_outFIFO/U477  ( .A(n1625), .B(n958), .C(\u_outFIFO/n754 ), .Q(
        \u_outFIFO/n1201 ) );
  OAI212 \u_outFIFO/U476  ( .A(n852), .B(n821), .C(n930), .Q(\u_outFIFO/n753 )
         );
  OAI212 \u_outFIFO/U475  ( .A(n1624), .B(\u_outFIFO/n660 ), .C(
        \u_outFIFO/FIFO[85][2] ), .Q(\u_outFIFO/n752 ) );
  OAI212 \u_outFIFO/U474  ( .A(n1624), .B(n959), .C(\u_outFIFO/n752 ), .Q(
        \u_outFIFO/n1200 ) );
  OAI212 \u_outFIFO/U473  ( .A(n853), .B(n818), .C(n930), .Q(\u_outFIFO/n751 )
         );
  OAI212 \u_outFIFO/U472  ( .A(n1623), .B(\u_outFIFO/n660 ), .C(
        \u_outFIFO/FIFO[85][1] ), .Q(\u_outFIFO/n750 ) );
  OAI212 \u_outFIFO/U471  ( .A(n1623), .B(n959), .C(\u_outFIFO/n750 ), .Q(
        \u_outFIFO/n1199 ) );
  OAI212 \u_outFIFO/U470  ( .A(n852), .B(n815), .C(n930), .Q(\u_outFIFO/n749 )
         );
  OAI212 \u_outFIFO/U469  ( .A(n1622), .B(\u_outFIFO/n660 ), .C(
        \u_outFIFO/FIFO[85][0] ), .Q(\u_outFIFO/n748 ) );
  OAI212 \u_outFIFO/U468  ( .A(n1622), .B(n959), .C(\u_outFIFO/n748 ), .Q(
        \u_outFIFO/n1198 ) );
  OAI212 \u_outFIFO/U467  ( .A(n850), .B(n823), .C(n930), .Q(\u_outFIFO/n747 )
         );
  OAI212 \u_outFIFO/U466  ( .A(n1621), .B(\u_outFIFO/n660 ), .C(
        \u_outFIFO/FIFO[84][3] ), .Q(\u_outFIFO/n746 ) );
  OAI212 \u_outFIFO/U465  ( .A(n1621), .B(n959), .C(\u_outFIFO/n746 ), .Q(
        \u_outFIFO/n1197 ) );
  OAI212 \u_outFIFO/U464  ( .A(n849), .B(n820), .C(n930), .Q(\u_outFIFO/n745 )
         );
  OAI212 \u_outFIFO/U463  ( .A(n1620), .B(\u_outFIFO/n660 ), .C(
        \u_outFIFO/FIFO[84][2] ), .Q(\u_outFIFO/n744 ) );
  OAI212 \u_outFIFO/U462  ( .A(n1620), .B(n959), .C(\u_outFIFO/n744 ), .Q(
        \u_outFIFO/n1196 ) );
  OAI212 \u_outFIFO/U461  ( .A(n850), .B(n817), .C(n930), .Q(\u_outFIFO/n743 )
         );
  OAI212 \u_outFIFO/U460  ( .A(n1619), .B(\u_outFIFO/n660 ), .C(
        \u_outFIFO/FIFO[84][1] ), .Q(\u_outFIFO/n742 ) );
  OAI212 \u_outFIFO/U459  ( .A(n1619), .B(n959), .C(\u_outFIFO/n742 ), .Q(
        \u_outFIFO/n1195 ) );
  OAI212 \u_outFIFO/U458  ( .A(n849), .B(n815), .C(n930), .Q(\u_outFIFO/n741 )
         );
  OAI212 \u_outFIFO/U457  ( .A(n1618), .B(\u_outFIFO/n660 ), .C(
        \u_outFIFO/FIFO[84][0] ), .Q(\u_outFIFO/n740 ) );
  OAI212 \u_outFIFO/U456  ( .A(n1618), .B(n959), .C(\u_outFIFO/n740 ), .Q(
        \u_outFIFO/n1194 ) );
  OAI212 \u_outFIFO/U455  ( .A(n844), .B(n824), .C(n930), .Q(\u_outFIFO/n739 )
         );
  OAI212 \u_outFIFO/U454  ( .A(n1617), .B(\u_outFIFO/n660 ), .C(
        \u_outFIFO/FIFO[83][3] ), .Q(\u_outFIFO/n738 ) );
  OAI212 \u_outFIFO/U453  ( .A(n1617), .B(n959), .C(\u_outFIFO/n738 ), .Q(
        \u_outFIFO/n1193 ) );
  OAI212 \u_outFIFO/U452  ( .A(n845), .B(n821), .C(n929), .Q(\u_outFIFO/n737 )
         );
  OAI212 \u_outFIFO/U451  ( .A(n1616), .B(n1184), .C(\u_outFIFO/FIFO[83][2] ), 
        .Q(\u_outFIFO/n736 ) );
  OAI212 \u_outFIFO/U450  ( .A(n1616), .B(n959), .C(\u_outFIFO/n736 ), .Q(
        \u_outFIFO/n1192 ) );
  OAI212 \u_outFIFO/U449  ( .A(n846), .B(n818), .C(n929), .Q(\u_outFIFO/n735 )
         );
  OAI212 \u_outFIFO/U448  ( .A(n1615), .B(n1184), .C(\u_outFIFO/FIFO[83][1] ), 
        .Q(\u_outFIFO/n734 ) );
  OAI212 \u_outFIFO/U447  ( .A(n1615), .B(n959), .C(\u_outFIFO/n734 ), .Q(
        \u_outFIFO/n1191 ) );
  OAI212 \u_outFIFO/U446  ( .A(n847), .B(n815), .C(n929), .Q(\u_outFIFO/n733 )
         );
  OAI212 \u_outFIFO/U445  ( .A(n1614), .B(n1184), .C(\u_outFIFO/FIFO[83][0] ), 
        .Q(\u_outFIFO/n732 ) );
  OAI212 \u_outFIFO/U444  ( .A(n1614), .B(n959), .C(\u_outFIFO/n732 ), .Q(
        \u_outFIFO/n1190 ) );
  OAI212 \u_outFIFO/U443  ( .A(n842), .B(n823), .C(n929), .Q(\u_outFIFO/n731 )
         );
  OAI212 \u_outFIFO/U442  ( .A(n1613), .B(n1187), .C(\u_outFIFO/FIFO[82][3] ), 
        .Q(\u_outFIFO/n730 ) );
  OAI212 \u_outFIFO/U441  ( .A(n1613), .B(n959), .C(\u_outFIFO/n730 ), .Q(
        \u_outFIFO/n1189 ) );
  OAI212 \u_outFIFO/U440  ( .A(\u_outFIFO/n331 ), .B(n820), .C(n929), .Q(
        \u_outFIFO/n729 ) );
  OAI212 \u_outFIFO/U439  ( .A(n1612), .B(n1188), .C(\u_outFIFO/FIFO[82][2] ), 
        .Q(\u_outFIFO/n728 ) );
  OAI212 \u_outFIFO/U438  ( .A(n1612), .B(n959), .C(\u_outFIFO/n728 ), .Q(
        \u_outFIFO/n1188 ) );
  OAI212 \u_outFIFO/U437  ( .A(n842), .B(n817), .C(n929), .Q(\u_outFIFO/n727 )
         );
  OAI212 \u_outFIFO/U436  ( .A(n1611), .B(n1189), .C(\u_outFIFO/FIFO[82][1] ), 
        .Q(\u_outFIFO/n726 ) );
  OAI212 \u_outFIFO/U435  ( .A(n1611), .B(n960), .C(\u_outFIFO/n726 ), .Q(
        \u_outFIFO/n1187 ) );
  OAI212 \u_outFIFO/U434  ( .A(n842), .B(n815), .C(n929), .Q(\u_outFIFO/n725 )
         );
  OAI212 \u_outFIFO/U433  ( .A(n1610), .B(n1190), .C(\u_outFIFO/FIFO[82][0] ), 
        .Q(\u_outFIFO/n724 ) );
  OAI212 \u_outFIFO/U432  ( .A(n1610), .B(n960), .C(\u_outFIFO/n724 ), .Q(
        \u_outFIFO/n1186 ) );
  OAI212 \u_outFIFO/U431  ( .A(n840), .B(n824), .C(n929), .Q(\u_outFIFO/n723 )
         );
  OAI212 \u_outFIFO/U430  ( .A(n1609), .B(n1187), .C(\u_outFIFO/FIFO[81][3] ), 
        .Q(\u_outFIFO/n722 ) );
  OAI212 \u_outFIFO/U429  ( .A(n1609), .B(n960), .C(\u_outFIFO/n722 ), .Q(
        \u_outFIFO/n1185 ) );
  OAI212 \u_outFIFO/U428  ( .A(n839), .B(n821), .C(n928), .Q(\u_outFIFO/n721 )
         );
  OAI212 \u_outFIFO/U427  ( .A(n1608), .B(n1188), .C(\u_outFIFO/FIFO[81][2] ), 
        .Q(\u_outFIFO/n720 ) );
  OAI212 \u_outFIFO/U426  ( .A(n1608), .B(n960), .C(\u_outFIFO/n720 ), .Q(
        \u_outFIFO/n1184 ) );
  OAI212 \u_outFIFO/U425  ( .A(n840), .B(n818), .C(n928), .Q(\u_outFIFO/n719 )
         );
  OAI212 \u_outFIFO/U424  ( .A(n1607), .B(n1188), .C(\u_outFIFO/FIFO[81][1] ), 
        .Q(\u_outFIFO/n718 ) );
  OAI212 \u_outFIFO/U423  ( .A(n1607), .B(n960), .C(\u_outFIFO/n718 ), .Q(
        \u_outFIFO/n1183 ) );
  OAI212 \u_outFIFO/U422  ( .A(n839), .B(n815), .C(n928), .Q(\u_outFIFO/n717 )
         );
  OAI212 \u_outFIFO/U421  ( .A(n1606), .B(n1188), .C(\u_outFIFO/FIFO[81][0] ), 
        .Q(\u_outFIFO/n716 ) );
  OAI212 \u_outFIFO/U420  ( .A(n1606), .B(n960), .C(\u_outFIFO/n716 ), .Q(
        \u_outFIFO/n1182 ) );
  OAI212 \u_outFIFO/U419  ( .A(\u_outFIFO/n317 ), .B(n823), .C(n928), .Q(
        \u_outFIFO/n714 ) );
  OAI212 \u_outFIFO/U418  ( .A(n1605), .B(n1188), .C(\u_outFIFO/FIFO[80][3] ), 
        .Q(\u_outFIFO/n713 ) );
  OAI212 \u_outFIFO/U417  ( .A(n1605), .B(n960), .C(\u_outFIFO/n713 ), .Q(
        \u_outFIFO/n1181 ) );
  OAI212 \u_outFIFO/U416  ( .A(n837), .B(n820), .C(n928), .Q(\u_outFIFO/n711 )
         );
  OAI212 \u_outFIFO/U415  ( .A(n1604), .B(n1188), .C(\u_outFIFO/FIFO[80][2] ), 
        .Q(\u_outFIFO/n710 ) );
  OAI212 \u_outFIFO/U414  ( .A(n1604), .B(n960), .C(\u_outFIFO/n710 ), .Q(
        \u_outFIFO/n1180 ) );
  OAI212 \u_outFIFO/U413  ( .A(\u_outFIFO/n317 ), .B(n817), .C(n928), .Q(
        \u_outFIFO/n708 ) );
  OAI212 \u_outFIFO/U412  ( .A(n1603), .B(n1188), .C(\u_outFIFO/FIFO[80][1] ), 
        .Q(\u_outFIFO/n707 ) );
  OAI212 \u_outFIFO/U411  ( .A(n1603), .B(n960), .C(\u_outFIFO/n707 ), .Q(
        \u_outFIFO/n1179 ) );
  OAI212 \u_outFIFO/U410  ( .A(\u_outFIFO/n317 ), .B(n815), .C(n928), .Q(
        \u_outFIFO/n705 ) );
  OAI212 \u_outFIFO/U409  ( .A(n1602), .B(n1188), .C(\u_outFIFO/FIFO[80][0] ), 
        .Q(\u_outFIFO/n704 ) );
  OAI212 \u_outFIFO/U408  ( .A(n1602), .B(n960), .C(\u_outFIFO/n704 ), .Q(
        \u_outFIFO/n1178 ) );
  OAI212 \u_outFIFO/U405  ( .A(\u_outFIFO/n396 ), .B(\u_outFIFO/n669 ), .C(
        n928), .Q(\u_outFIFO/n703 ) );
  OAI212 \u_outFIFO/U404  ( .A(n1601), .B(n1188), .C(\u_outFIFO/FIFO[79][3] ), 
        .Q(\u_outFIFO/n702 ) );
  OAI212 \u_outFIFO/U403  ( .A(n1601), .B(n960), .C(\u_outFIFO/n702 ), .Q(
        \u_outFIFO/n1177 ) );
  OAI212 \u_outFIFO/U401  ( .A(n889), .B(\u_outFIFO/n677 ), .C(n927), .Q(
        \u_outFIFO/n701 ) );
  OAI212 \u_outFIFO/U400  ( .A(n1600), .B(n1188), .C(\u_outFIFO/FIFO[79][2] ), 
        .Q(\u_outFIFO/n700 ) );
  OAI212 \u_outFIFO/U399  ( .A(n1600), .B(n960), .C(\u_outFIFO/n700 ), .Q(
        \u_outFIFO/n1176 ) );
  OAI212 \u_outFIFO/U397  ( .A(\u_outFIFO/n396 ), .B(\u_outFIFO/n674 ), .C(
        n927), .Q(\u_outFIFO/n699 ) );
  OAI212 \u_outFIFO/U396  ( .A(n1599), .B(n1188), .C(\u_outFIFO/FIFO[79][1] ), 
        .Q(\u_outFIFO/n698 ) );
  OAI212 \u_outFIFO/U395  ( .A(n1599), .B(n960), .C(\u_outFIFO/n698 ), .Q(
        \u_outFIFO/n1175 ) );
  OAI212 \u_outFIFO/U393  ( .A(n889), .B(n812), .C(n927), .Q(\u_outFIFO/n697 )
         );
  OAI212 \u_outFIFO/U392  ( .A(n1598), .B(n1188), .C(\u_outFIFO/FIFO[79][0] ), 
        .Q(\u_outFIFO/n696 ) );
  OAI212 \u_outFIFO/U391  ( .A(n1598), .B(n961), .C(\u_outFIFO/n696 ), .Q(
        \u_outFIFO/n1174 ) );
  OAI212 \u_outFIFO/U390  ( .A(\u_outFIFO/n391 ), .B(\u_outFIFO/n669 ), .C(
        n927), .Q(\u_outFIFO/n695 ) );
  OAI212 \u_outFIFO/U389  ( .A(n1597), .B(n1188), .C(\u_outFIFO/FIFO[78][3] ), 
        .Q(\u_outFIFO/n694 ) );
  OAI212 \u_outFIFO/U388  ( .A(n1597), .B(n961), .C(\u_outFIFO/n694 ), .Q(
        \u_outFIFO/n1173 ) );
  OAI212 \u_outFIFO/U387  ( .A(n877), .B(\u_outFIFO/n677 ), .C(n927), .Q(
        \u_outFIFO/n693 ) );
  OAI212 \u_outFIFO/U386  ( .A(n1596), .B(n1188), .C(\u_outFIFO/FIFO[78][2] ), 
        .Q(\u_outFIFO/n692 ) );
  OAI212 \u_outFIFO/U385  ( .A(n1596), .B(n961), .C(\u_outFIFO/n692 ), .Q(
        \u_outFIFO/n1172 ) );
  OAI212 \u_outFIFO/U384  ( .A(\u_outFIFO/n391 ), .B(\u_outFIFO/n674 ), .C(
        n927), .Q(\u_outFIFO/n691 ) );
  OAI212 \u_outFIFO/U383  ( .A(n1595), .B(n1188), .C(\u_outFIFO/FIFO[78][1] ), 
        .Q(\u_outFIFO/n690 ) );
  OAI212 \u_outFIFO/U382  ( .A(n1595), .B(n961), .C(\u_outFIFO/n690 ), .Q(
        \u_outFIFO/n1171 ) );
  OAI212 \u_outFIFO/U381  ( .A(n877), .B(n812), .C(n927), .Q(\u_outFIFO/n689 )
         );
  OAI212 \u_outFIFO/U380  ( .A(n1594), .B(n1188), .C(\u_outFIFO/FIFO[78][0] ), 
        .Q(\u_outFIFO/n688 ) );
  OAI212 \u_outFIFO/U379  ( .A(n1594), .B(n961), .C(\u_outFIFO/n688 ), .Q(
        \u_outFIFO/n1170 ) );
  OAI212 \u_outFIFO/U378  ( .A(\u_outFIFO/n386 ), .B(\u_outFIFO/n669 ), .C(
        n927), .Q(\u_outFIFO/n687 ) );
  OAI212 \u_outFIFO/U377  ( .A(n1593), .B(n1188), .C(\u_outFIFO/FIFO[77][3] ), 
        .Q(\u_outFIFO/n686 ) );
  OAI212 \u_outFIFO/U376  ( .A(n1593), .B(n961), .C(\u_outFIFO/n686 ), .Q(
        \u_outFIFO/n1169 ) );
  OAI212 \u_outFIFO/U375  ( .A(n875), .B(\u_outFIFO/n677 ), .C(n926), .Q(
        \u_outFIFO/n685 ) );
  OAI212 \u_outFIFO/U374  ( .A(n1592), .B(n1188), .C(\u_outFIFO/FIFO[77][2] ), 
        .Q(\u_outFIFO/n684 ) );
  OAI212 \u_outFIFO/U373  ( .A(n1592), .B(n961), .C(\u_outFIFO/n684 ), .Q(
        \u_outFIFO/n1168 ) );
  OAI212 \u_outFIFO/U372  ( .A(\u_outFIFO/n386 ), .B(\u_outFIFO/n674 ), .C(
        n926), .Q(\u_outFIFO/n683 ) );
  OAI212 \u_outFIFO/U371  ( .A(n1591), .B(n1188), .C(\u_outFIFO/FIFO[77][1] ), 
        .Q(\u_outFIFO/n682 ) );
  OAI212 \u_outFIFO/U370  ( .A(n1591), .B(n961), .C(\u_outFIFO/n682 ), .Q(
        \u_outFIFO/n1167 ) );
  OAI212 \u_outFIFO/U369  ( .A(n875), .B(n812), .C(n926), .Q(\u_outFIFO/n681 )
         );
  OAI212 \u_outFIFO/U368  ( .A(n1590), .B(n1186), .C(\u_outFIFO/FIFO[77][0] ), 
        .Q(\u_outFIFO/n680 ) );
  OAI212 \u_outFIFO/U367  ( .A(n1590), .B(n961), .C(\u_outFIFO/n680 ), .Q(
        \u_outFIFO/n1166 ) );
  OAI212 \u_outFIFO/U366  ( .A(n873), .B(\u_outFIFO/n669 ), .C(n926), .Q(
        \u_outFIFO/n679 ) );
  OAI212 \u_outFIFO/U365  ( .A(n1589), .B(n1185), .C(\u_outFIFO/FIFO[76][3] ), 
        .Q(\u_outFIFO/n678 ) );
  OAI212 \u_outFIFO/U364  ( .A(n1589), .B(n961), .C(\u_outFIFO/n678 ), .Q(
        \u_outFIFO/n1165 ) );
  OAI212 \u_outFIFO/U363  ( .A(n873), .B(\u_outFIFO/n677 ), .C(n926), .Q(
        \u_outFIFO/n676 ) );
  OAI212 \u_outFIFO/U362  ( .A(n1588), .B(n1190), .C(\u_outFIFO/FIFO[76][2] ), 
        .Q(\u_outFIFO/n675 ) );
  OAI212 \u_outFIFO/U361  ( .A(n1588), .B(n961), .C(\u_outFIFO/n675 ), .Q(
        \u_outFIFO/n1164 ) );
  OAI212 \u_outFIFO/U360  ( .A(n873), .B(\u_outFIFO/n674 ), .C(n926), .Q(
        \u_outFIFO/n673 ) );
  OAI212 \u_outFIFO/U359  ( .A(n1587), .B(n1186), .C(\u_outFIFO/FIFO[76][1] ), 
        .Q(\u_outFIFO/n672 ) );
  OAI212 \u_outFIFO/U358  ( .A(n1587), .B(n961), .C(\u_outFIFO/n672 ), .Q(
        \u_outFIFO/n1163 ) );
  OAI212 \u_outFIFO/U357  ( .A(n873), .B(n812), .C(n926), .Q(\u_outFIFO/n671 )
         );
  OAI212 \u_outFIFO/U356  ( .A(n1586), .B(n1187), .C(\u_outFIFO/FIFO[76][0] ), 
        .Q(\u_outFIFO/n670 ) );
  OAI212 \u_outFIFO/U355  ( .A(n1586), .B(n961), .C(\u_outFIFO/n670 ), .Q(
        \u_outFIFO/n1162 ) );
  OAI212 \u_outFIFO/U354  ( .A(n871), .B(\u_outFIFO/n669 ), .C(n926), .Q(
        \u_outFIFO/n668 ) );
  OAI212 \u_outFIFO/U353  ( .A(n1585), .B(n1185), .C(\u_outFIFO/FIFO[75][3] ), 
        .Q(\u_outFIFO/n667 ) );
  OAI212 \u_outFIFO/U352  ( .A(n1585), .B(n1795), .C(\u_outFIFO/n667 ), .Q(
        \u_outFIFO/n1161 ) );
  OAI212 \u_outFIFO/U349  ( .A(n870), .B(\u_outFIFO/n616 ), .C(n1225), .Q(
        \u_outFIFO/n665 ) );
  OAI212 \u_outFIFO/U346  ( .A(n871), .B(\u_outFIFO/n614 ), .C(n1225), .Q(
        \u_outFIFO/n663 ) );
  OAI212 \u_outFIFO/U345  ( .A(n870), .B(n812), .C(n1225), .Q(\u_outFIFO/n662 ) );
  OAI212 \u_outFIFO/U342  ( .A(n868), .B(\u_outFIFO/n618 ), .C(n1225), .Q(
        \u_outFIFO/n658 ) );
  OAI212 \u_outFIFO/U341  ( .A(n867), .B(\u_outFIFO/n616 ), .C(n1225), .Q(
        \u_outFIFO/n657 ) );
  OAI212 \u_outFIFO/U340  ( .A(n868), .B(\u_outFIFO/n614 ), .C(n1225), .Q(
        \u_outFIFO/n656 ) );
  OAI212 \u_outFIFO/U339  ( .A(n867), .B(n812), .C(n1225), .Q(\u_outFIFO/n655 ) );
  OAI212 \u_outFIFO/U338  ( .A(n865), .B(\u_outFIFO/n618 ), .C(n1225), .Q(
        \u_outFIFO/n654 ) );
  OAI212 \u_outFIFO/U337  ( .A(n864), .B(\u_outFIFO/n616 ), .C(n1225), .Q(
        \u_outFIFO/n653 ) );
  OAI212 \u_outFIFO/U336  ( .A(n865), .B(\u_outFIFO/n614 ), .C(n1225), .Q(
        \u_outFIFO/n652 ) );
  OAI212 \u_outFIFO/U335  ( .A(n864), .B(n812), .C(n1224), .Q(\u_outFIFO/n651 ) );
  OAI212 \u_outFIFO/U334  ( .A(n862), .B(\u_outFIFO/n618 ), .C(n1224), .Q(
        \u_outFIFO/n650 ) );
  OAI212 \u_outFIFO/U333  ( .A(n861), .B(\u_outFIFO/n616 ), .C(n1224), .Q(
        \u_outFIFO/n649 ) );
  OAI212 \u_outFIFO/U332  ( .A(n862), .B(\u_outFIFO/n614 ), .C(n1224), .Q(
        \u_outFIFO/n648 ) );
  OAI212 \u_outFIFO/U331  ( .A(n861), .B(n812), .C(n1224), .Q(\u_outFIFO/n647 ) );
  OAI212 \u_outFIFO/U330  ( .A(n859), .B(\u_outFIFO/n618 ), .C(n1224), .Q(
        \u_outFIFO/n646 ) );
  OAI212 \u_outFIFO/U329  ( .A(n858), .B(\u_outFIFO/n616 ), .C(n1224), .Q(
        \u_outFIFO/n645 ) );
  OAI212 \u_outFIFO/U328  ( .A(n859), .B(\u_outFIFO/n614 ), .C(n1224), .Q(
        \u_outFIFO/n644 ) );
  OAI212 \u_outFIFO/U327  ( .A(n858), .B(n813), .C(n1224), .Q(\u_outFIFO/n643 ) );
  OAI212 \u_outFIFO/U326  ( .A(n856), .B(\u_outFIFO/n618 ), .C(n1224), .Q(
        \u_outFIFO/n642 ) );
  OAI212 \u_outFIFO/U325  ( .A(n855), .B(\u_outFIFO/n616 ), .C(n1224), .Q(
        \u_outFIFO/n641 ) );
  OAI212 \u_outFIFO/U324  ( .A(n856), .B(\u_outFIFO/n614 ), .C(n1224), .Q(
        \u_outFIFO/n640 ) );
  OAI212 \u_outFIFO/U323  ( .A(n855), .B(n813), .C(n1224), .Q(\u_outFIFO/n639 ) );
  OAI212 \u_outFIFO/U322  ( .A(n853), .B(\u_outFIFO/n618 ), .C(n1224), .Q(
        \u_outFIFO/n638 ) );
  OAI212 \u_outFIFO/U321  ( .A(n852), .B(\u_outFIFO/n616 ), .C(n1224), .Q(
        \u_outFIFO/n637 ) );
  OAI212 \u_outFIFO/U320  ( .A(n853), .B(\u_outFIFO/n614 ), .C(n1224), .Q(
        \u_outFIFO/n636 ) );
  OAI212 \u_outFIFO/U319  ( .A(n852), .B(n813), .C(n1224), .Q(\u_outFIFO/n635 ) );
  OAI212 \u_outFIFO/U318  ( .A(n850), .B(\u_outFIFO/n618 ), .C(n1224), .Q(
        \u_outFIFO/n634 ) );
  OAI212 \u_outFIFO/U317  ( .A(n849), .B(\u_outFIFO/n616 ), .C(n1224), .Q(
        \u_outFIFO/n633 ) );
  OAI212 \u_outFIFO/U316  ( .A(n850), .B(\u_outFIFO/n614 ), .C(n1224), .Q(
        \u_outFIFO/n632 ) );
  OAI212 \u_outFIFO/U315  ( .A(n849), .B(n813), .C(n1224), .Q(\u_outFIFO/n631 ) );
  OAI212 \u_outFIFO/U314  ( .A(n844), .B(\u_outFIFO/n618 ), .C(n1224), .Q(
        \u_outFIFO/n630 ) );
  OAI212 \u_outFIFO/U313  ( .A(n845), .B(\u_outFIFO/n616 ), .C(n1224), .Q(
        \u_outFIFO/n629 ) );
  OAI212 \u_outFIFO/U312  ( .A(n846), .B(\u_outFIFO/n614 ), .C(n1224), .Q(
        \u_outFIFO/n628 ) );
  OAI212 \u_outFIFO/U311  ( .A(n847), .B(n813), .C(n1224), .Q(\u_outFIFO/n627 ) );
  OAI212 \u_outFIFO/U310  ( .A(n842), .B(\u_outFIFO/n618 ), .C(n1224), .Q(
        \u_outFIFO/n626 ) );
  OAI212 \u_outFIFO/U309  ( .A(n842), .B(\u_outFIFO/n616 ), .C(n1224), .Q(
        \u_outFIFO/n625 ) );
  OAI212 \u_outFIFO/U308  ( .A(\u_outFIFO/n331 ), .B(\u_outFIFO/n614 ), .C(
        n1223), .Q(\u_outFIFO/n624 ) );
  OAI212 \u_outFIFO/U307  ( .A(\u_outFIFO/n331 ), .B(n813), .C(n1223), .Q(
        \u_outFIFO/n623 ) );
  OAI212 \u_outFIFO/U306  ( .A(n840), .B(\u_outFIFO/n618 ), .C(n1223), .Q(
        \u_outFIFO/n622 ) );
  OAI212 \u_outFIFO/U305  ( .A(n839), .B(\u_outFIFO/n616 ), .C(n1223), .Q(
        \u_outFIFO/n621 ) );
  OAI212 \u_outFIFO/U304  ( .A(n840), .B(\u_outFIFO/n614 ), .C(n1223), .Q(
        \u_outFIFO/n620 ) );
  OAI212 \u_outFIFO/U303  ( .A(n839), .B(n813), .C(n1223), .Q(\u_outFIFO/n619 ) );
  OAI212 \u_outFIFO/U302  ( .A(n837), .B(\u_outFIFO/n618 ), .C(n1223), .Q(
        \u_outFIFO/n617 ) );
  OAI212 \u_outFIFO/U301  ( .A(n837), .B(\u_outFIFO/n616 ), .C(n1223), .Q(
        \u_outFIFO/n615 ) );
  OAI212 \u_outFIFO/U300  ( .A(n837), .B(\u_outFIFO/n614 ), .C(n1223), .Q(
        \u_outFIFO/n613 ) );
  OAI212 \u_outFIFO/U299  ( .A(\u_outFIFO/n317 ), .B(n813), .C(n1223), .Q(
        \u_outFIFO/n611 ) );
  OAI212 \u_outFIFO/U296  ( .A(\u_outFIFO/n396 ), .B(n809), .C(n1223), .Q(
        \u_outFIFO/n610 ) );
  OAI212 \u_outFIFO/U294  ( .A(n889), .B(n806), .C(n1223), .Q(\u_outFIFO/n609 ) );
  OAI212 \u_outFIFO/U292  ( .A(\u_outFIFO/n396 ), .B(n804), .C(n1223), .Q(
        \u_outFIFO/n608 ) );
  OAI212 \u_outFIFO/U290  ( .A(n889), .B(n802), .C(n1223), .Q(\u_outFIFO/n606 ) );
  OAI212 \u_outFIFO/U289  ( .A(\u_outFIFO/n391 ), .B(n809), .C(n1223), .Q(
        \u_outFIFO/n605 ) );
  OAI212 \u_outFIFO/U288  ( .A(n877), .B(n806), .C(n1223), .Q(\u_outFIFO/n604 ) );
  OAI212 \u_outFIFO/U287  ( .A(\u_outFIFO/n391 ), .B(n804), .C(n1223), .Q(
        \u_outFIFO/n603 ) );
  OAI212 \u_outFIFO/U286  ( .A(n877), .B(n802), .C(n1223), .Q(\u_outFIFO/n602 ) );
  OAI212 \u_outFIFO/U285  ( .A(\u_outFIFO/n386 ), .B(n809), .C(n1223), .Q(
        \u_outFIFO/n601 ) );
  OAI212 \u_outFIFO/U284  ( .A(n875), .B(n806), .C(n1223), .Q(\u_outFIFO/n600 ) );
  OAI212 \u_outFIFO/U283  ( .A(\u_outFIFO/n386 ), .B(n804), .C(n1223), .Q(
        \u_outFIFO/n599 ) );
  OAI212 \u_outFIFO/U282  ( .A(n875), .B(n802), .C(n1223), .Q(\u_outFIFO/n598 ) );
  OAI212 \u_outFIFO/U281  ( .A(n873), .B(n809), .C(n1223), .Q(\u_outFIFO/n597 ) );
  OAI212 \u_outFIFO/U280  ( .A(\u_outFIFO/n381 ), .B(n806), .C(n1223), .Q(
        \u_outFIFO/n596 ) );
  OAI212 \u_outFIFO/U279  ( .A(\u_outFIFO/n381 ), .B(n804), .C(n1223), .Q(
        \u_outFIFO/n595 ) );
  OAI212 \u_outFIFO/U278  ( .A(\u_outFIFO/n381 ), .B(n802), .C(n1223), .Q(
        \u_outFIFO/n594 ) );
  OAI212 \u_outFIFO/U277  ( .A(n871), .B(n809), .C(n1223), .Q(\u_outFIFO/n593 ) );
  OAI212 \u_outFIFO/U276  ( .A(n870), .B(n806), .C(n1222), .Q(\u_outFIFO/n592 ) );
  OAI212 \u_outFIFO/U275  ( .A(n871), .B(n804), .C(n1222), .Q(\u_outFIFO/n591 ) );
  OAI212 \u_outFIFO/U274  ( .A(n870), .B(n802), .C(n1222), .Q(\u_outFIFO/n590 ) );
  OAI212 \u_outFIFO/U273  ( .A(n868), .B(n809), .C(n1222), .Q(\u_outFIFO/n589 ) );
  OAI212 \u_outFIFO/U272  ( .A(n867), .B(n806), .C(n1222), .Q(\u_outFIFO/n588 ) );
  OAI212 \u_outFIFO/U271  ( .A(n868), .B(n804), .C(n1222), .Q(\u_outFIFO/n587 ) );
  OAI212 \u_outFIFO/U270  ( .A(n867), .B(n802), .C(n1222), .Q(\u_outFIFO/n586 ) );
  OAI212 \u_outFIFO/U269  ( .A(n865), .B(n811), .C(n1222), .Q(\u_outFIFO/n585 ) );
  OAI212 \u_outFIFO/U268  ( .A(n864), .B(n808), .C(n1222), .Q(\u_outFIFO/n584 ) );
  OAI212 \u_outFIFO/U267  ( .A(n865), .B(n804), .C(n1222), .Q(\u_outFIFO/n583 ) );
  OAI212 \u_outFIFO/U266  ( .A(n864), .B(n802), .C(n1222), .Q(\u_outFIFO/n582 ) );
  OAI212 \u_outFIFO/U265  ( .A(n862), .B(n810), .C(n1222), .Q(\u_outFIFO/n581 ) );
  OAI212 \u_outFIFO/U264  ( .A(n861), .B(n807), .C(n1225), .Q(\u_outFIFO/n580 ) );
  OAI212 \u_outFIFO/U263  ( .A(n862), .B(n804), .C(n1222), .Q(\u_outFIFO/n579 ) );
  OAI212 \u_outFIFO/U262  ( .A(n861), .B(n802), .C(n1222), .Q(\u_outFIFO/n578 ) );
  OAI212 \u_outFIFO/U261  ( .A(n859), .B(n811), .C(n1222), .Q(\u_outFIFO/n577 ) );
  OAI212 \u_outFIFO/U260  ( .A(n858), .B(n808), .C(n1222), .Q(\u_outFIFO/n576 ) );
  OAI212 \u_outFIFO/U259  ( .A(n859), .B(n805), .C(n1222), .Q(\u_outFIFO/n575 ) );
  OAI212 \u_outFIFO/U258  ( .A(n858), .B(n803), .C(n1222), .Q(\u_outFIFO/n574 ) );
  OAI212 \u_outFIFO/U257  ( .A(n856), .B(n810), .C(n1222), .Q(\u_outFIFO/n573 ) );
  OAI212 \u_outFIFO/U256  ( .A(n855), .B(n807), .C(n1222), .Q(\u_outFIFO/n572 ) );
  OAI212 \u_outFIFO/U255  ( .A(n856), .B(n805), .C(n1222), .Q(\u_outFIFO/n571 ) );
  OAI212 \u_outFIFO/U254  ( .A(n855), .B(n803), .C(n1222), .Q(\u_outFIFO/n570 ) );
  OAI212 \u_outFIFO/U253  ( .A(n853), .B(n811), .C(n1222), .Q(\u_outFIFO/n569 ) );
  OAI212 \u_outFIFO/U252  ( .A(n852), .B(n808), .C(n1222), .Q(\u_outFIFO/n568 ) );
  OAI212 \u_outFIFO/U251  ( .A(n853), .B(n805), .C(n1222), .Q(\u_outFIFO/n567 ) );
  OAI212 \u_outFIFO/U250  ( .A(n852), .B(n803), .C(n1221), .Q(\u_outFIFO/n566 ) );
  OAI212 \u_outFIFO/U249  ( .A(n850), .B(n810), .C(n1221), .Q(\u_outFIFO/n565 ) );
  OAI212 \u_outFIFO/U248  ( .A(n849), .B(n807), .C(n1221), .Q(\u_outFIFO/n564 ) );
  OAI212 \u_outFIFO/U247  ( .A(n850), .B(n805), .C(n1221), .Q(\u_outFIFO/n563 ) );
  OAI212 \u_outFIFO/U246  ( .A(n849), .B(n803), .C(n1222), .Q(\u_outFIFO/n562 ) );
  OAI212 \u_outFIFO/U245  ( .A(n844), .B(n811), .C(n1221), .Q(\u_outFIFO/n561 ) );
  OAI212 \u_outFIFO/U244  ( .A(n845), .B(n808), .C(n1221), .Q(\u_outFIFO/n560 ) );
  OAI212 \u_outFIFO/U243  ( .A(n846), .B(n805), .C(n1221), .Q(\u_outFIFO/n559 ) );
  OAI212 \u_outFIFO/U242  ( .A(n847), .B(n803), .C(n1221), .Q(\u_outFIFO/n558 ) );
  OAI212 \u_outFIFO/U241  ( .A(n842), .B(n810), .C(n1221), .Q(\u_outFIFO/n557 ) );
  OAI212 \u_outFIFO/U240  ( .A(\u_outFIFO/n331 ), .B(n807), .C(n1221), .Q(
        \u_outFIFO/n556 ) );
  OAI212 \u_outFIFO/U239  ( .A(\u_outFIFO/n331 ), .B(n805), .C(n1221), .Q(
        \u_outFIFO/n555 ) );
  OAI212 \u_outFIFO/U238  ( .A(\u_outFIFO/n331 ), .B(n803), .C(n1221), .Q(
        \u_outFIFO/n554 ) );
  OAI212 \u_outFIFO/U237  ( .A(n840), .B(n811), .C(n1221), .Q(\u_outFIFO/n553 ) );
  OAI212 \u_outFIFO/U236  ( .A(n839), .B(n808), .C(n1221), .Q(\u_outFIFO/n552 ) );
  OAI212 \u_outFIFO/U235  ( .A(n840), .B(n805), .C(n1221), .Q(\u_outFIFO/n551 ) );
  OAI212 \u_outFIFO/U234  ( .A(n839), .B(n803), .C(n1221), .Q(\u_outFIFO/n550 ) );
  OAI212 \u_outFIFO/U233  ( .A(\u_outFIFO/n317 ), .B(n810), .C(n1221), .Q(
        \u_outFIFO/n548 ) );
  OAI212 \u_outFIFO/U232  ( .A(n837), .B(n807), .C(n1221), .Q(\u_outFIFO/n546 ) );
  OAI212 \u_outFIFO/U231  ( .A(\u_outFIFO/n317 ), .B(n805), .C(n1221), .Q(
        \u_outFIFO/n544 ) );
  OAI212 \u_outFIFO/U230  ( .A(\u_outFIFO/n317 ), .B(n803), .C(n1221), .Q(
        \u_outFIFO/n542 ) );
  OAI212 \u_outFIFO/U227  ( .A(\u_outFIFO/n396 ), .B(n799), .C(n1221), .Q(
        \u_outFIFO/n541 ) );
  OAI212 \u_outFIFO/U225  ( .A(n889), .B(n796), .C(n1221), .Q(\u_outFIFO/n540 ) );
  OAI212 \u_outFIFO/U223  ( .A(\u_outFIFO/n396 ), .B(n793), .C(n1221), .Q(
        \u_outFIFO/n539 ) );
  OAI212 \u_outFIFO/U221  ( .A(n889), .B(n791), .C(n1221), .Q(\u_outFIFO/n537 ) );
  OAI212 \u_outFIFO/U220  ( .A(\u_outFIFO/n391 ), .B(n799), .C(n1221), .Q(
        \u_outFIFO/n536 ) );
  OAI212 \u_outFIFO/U219  ( .A(n877), .B(n796), .C(n1221), .Q(\u_outFIFO/n535 ) );
  OAI212 \u_outFIFO/U218  ( .A(\u_outFIFO/n391 ), .B(n793), .C(n1220), .Q(
        \u_outFIFO/n534 ) );
  OAI212 \u_outFIFO/U217  ( .A(n877), .B(n791), .C(n1221), .Q(\u_outFIFO/n533 ) );
  OAI212 \u_outFIFO/U216  ( .A(\u_outFIFO/n386 ), .B(n799), .C(n1220), .Q(
        \u_outFIFO/n532 ) );
  OAI212 \u_outFIFO/U215  ( .A(n875), .B(n796), .C(n1220), .Q(\u_outFIFO/n531 ) );
  OAI212 \u_outFIFO/U214  ( .A(\u_outFIFO/n386 ), .B(n793), .C(n1220), .Q(
        \u_outFIFO/n530 ) );
  OAI212 \u_outFIFO/U213  ( .A(n875), .B(n791), .C(n1220), .Q(\u_outFIFO/n529 ) );
  OAI212 \u_outFIFO/U212  ( .A(n873), .B(n799), .C(n1220), .Q(\u_outFIFO/n528 ) );
  OAI212 \u_outFIFO/U211  ( .A(\u_outFIFO/n381 ), .B(n796), .C(n1220), .Q(
        \u_outFIFO/n527 ) );
  OAI212 \u_outFIFO/U210  ( .A(\u_outFIFO/n381 ), .B(n793), .C(n1220), .Q(
        \u_outFIFO/n526 ) );
  OAI212 \u_outFIFO/U209  ( .A(\u_outFIFO/n381 ), .B(n791), .C(n1220), .Q(
        \u_outFIFO/n525 ) );
  OAI212 \u_outFIFO/U208  ( .A(n871), .B(n799), .C(n1220), .Q(\u_outFIFO/n524 ) );
  OAI212 \u_outFIFO/U207  ( .A(n870), .B(n796), .C(n1220), .Q(\u_outFIFO/n523 ) );
  OAI212 \u_outFIFO/U206  ( .A(n871), .B(n793), .C(n1220), .Q(\u_outFIFO/n522 ) );
  OAI212 \u_outFIFO/U205  ( .A(n870), .B(n791), .C(n1220), .Q(\u_outFIFO/n521 ) );
  OAI212 \u_outFIFO/U204  ( .A(n868), .B(n799), .C(n1220), .Q(\u_outFIFO/n520 ) );
  OAI212 \u_outFIFO/U203  ( .A(n867), .B(n796), .C(n1220), .Q(\u_outFIFO/n519 ) );
  OAI212 \u_outFIFO/U202  ( .A(n868), .B(n793), .C(n1220), .Q(\u_outFIFO/n518 ) );
  OAI212 \u_outFIFO/U201  ( .A(n867), .B(n791), .C(n1220), .Q(\u_outFIFO/n517 ) );
  OAI212 \u_outFIFO/U200  ( .A(n865), .B(n801), .C(n1220), .Q(\u_outFIFO/n516 ) );
  OAI212 \u_outFIFO/U199  ( .A(n864), .B(n798), .C(n1220), .Q(\u_outFIFO/n515 ) );
  OAI212 \u_outFIFO/U198  ( .A(n865), .B(n795), .C(n1220), .Q(\u_outFIFO/n514 ) );
  OAI212 \u_outFIFO/U197  ( .A(n864), .B(n791), .C(n1220), .Q(\u_outFIFO/n513 ) );
  OAI212 \u_outFIFO/U196  ( .A(n862), .B(n800), .C(n1220), .Q(\u_outFIFO/n512 ) );
  OAI212 \u_outFIFO/U195  ( .A(n861), .B(n797), .C(n1220), .Q(\u_outFIFO/n511 ) );
  OAI212 \u_outFIFO/U194  ( .A(n862), .B(n794), .C(n1220), .Q(\u_outFIFO/n510 ) );
  OAI212 \u_outFIFO/U193  ( .A(n861), .B(n791), .C(n1222), .Q(\u_outFIFO/n509 ) );
  OAI212 \u_outFIFO/U192  ( .A(n859), .B(n801), .C(n1230), .Q(\u_outFIFO/n508 ) );
  OAI212 \u_outFIFO/U191  ( .A(n858), .B(n798), .C(n1231), .Q(\u_outFIFO/n507 ) );
  OAI212 \u_outFIFO/U190  ( .A(n859), .B(n795), .C(n1231), .Q(\u_outFIFO/n506 ) );
  OAI212 \u_outFIFO/U189  ( .A(n858), .B(n792), .C(n1231), .Q(\u_outFIFO/n505 ) );
  OAI212 \u_outFIFO/U188  ( .A(n856), .B(n800), .C(n1231), .Q(\u_outFIFO/n504 ) );
  OAI212 \u_outFIFO/U187  ( .A(n855), .B(n797), .C(n1231), .Q(\u_outFIFO/n503 ) );
  OAI212 \u_outFIFO/U186  ( .A(n856), .B(n794), .C(n1231), .Q(\u_outFIFO/n502 ) );
  OAI212 \u_outFIFO/U185  ( .A(n855), .B(n792), .C(n1231), .Q(\u_outFIFO/n501 ) );
  OAI212 \u_outFIFO/U184  ( .A(n853), .B(n801), .C(n1231), .Q(\u_outFIFO/n500 ) );
  OAI212 \u_outFIFO/U183  ( .A(n852), .B(n798), .C(n1231), .Q(\u_outFIFO/n499 ) );
  OAI212 \u_outFIFO/U182  ( .A(n853), .B(n795), .C(n1231), .Q(\u_outFIFO/n498 ) );
  OAI212 \u_outFIFO/U181  ( .A(n852), .B(n792), .C(n1231), .Q(\u_outFIFO/n497 ) );
  OAI212 \u_outFIFO/U180  ( .A(n850), .B(n800), .C(n1230), .Q(\u_outFIFO/n496 ) );
  OAI212 \u_outFIFO/U179  ( .A(n849), .B(n797), .C(n1230), .Q(\u_outFIFO/n495 ) );
  OAI212 \u_outFIFO/U178  ( .A(n850), .B(n794), .C(n1230), .Q(\u_outFIFO/n494 ) );
  OAI212 \u_outFIFO/U177  ( .A(n849), .B(n792), .C(n1230), .Q(\u_outFIFO/n493 ) );
  OAI212 \u_outFIFO/U176  ( .A(n844), .B(n801), .C(n1230), .Q(\u_outFIFO/n492 ) );
  OAI212 \u_outFIFO/U175  ( .A(n845), .B(n798), .C(n1230), .Q(\u_outFIFO/n491 ) );
  OAI212 \u_outFIFO/U174  ( .A(n846), .B(n795), .C(n1230), .Q(\u_outFIFO/n490 ) );
  OAI212 \u_outFIFO/U173  ( .A(n847), .B(n792), .C(n1230), .Q(\u_outFIFO/n489 ) );
  OAI212 \u_outFIFO/U172  ( .A(n842), .B(n800), .C(n1230), .Q(\u_outFIFO/n488 ) );
  OAI212 \u_outFIFO/U171  ( .A(\u_outFIFO/n331 ), .B(n797), .C(n1230), .Q(
        \u_outFIFO/n487 ) );
  OAI212 \u_outFIFO/U170  ( .A(\u_outFIFO/n331 ), .B(n794), .C(n1230), .Q(
        \u_outFIFO/n486 ) );
  OAI212 \u_outFIFO/U169  ( .A(\u_outFIFO/n331 ), .B(n792), .C(n1230), .Q(
        \u_outFIFO/n485 ) );
  OAI212 \u_outFIFO/U168  ( .A(n840), .B(n801), .C(n1230), .Q(\u_outFIFO/n484 ) );
  OAI212 \u_outFIFO/U167  ( .A(n839), .B(n798), .C(n1230), .Q(\u_outFIFO/n483 ) );
  OAI212 \u_outFIFO/U166  ( .A(n840), .B(n795), .C(n1230), .Q(\u_outFIFO/n482 ) );
  OAI212 \u_outFIFO/U165  ( .A(n839), .B(n792), .C(n1230), .Q(\u_outFIFO/n481 ) );
  OAI212 \u_outFIFO/U164  ( .A(\u_outFIFO/n317 ), .B(n800), .C(n1230), .Q(
        \u_outFIFO/n479 ) );
  OAI212 \u_outFIFO/U163  ( .A(\u_outFIFO/n317 ), .B(n797), .C(n1230), .Q(
        \u_outFIFO/n477 ) );
  OAI212 \u_outFIFO/U162  ( .A(\u_outFIFO/n317 ), .B(n794), .C(n1230), .Q(
        \u_outFIFO/n475 ) );
  OAI212 \u_outFIFO/U161  ( .A(\u_outFIFO/n317 ), .B(n792), .C(n1230), .Q(
        \u_outFIFO/n473 ) );
  OAI212 \u_outFIFO/U158  ( .A(\u_outFIFO/n396 ), .B(n788), .C(n1230), .Q(
        \u_outFIFO/n472 ) );
  OAI212 \u_outFIFO/U156  ( .A(\u_outFIFO/n396 ), .B(n785), .C(n1230), .Q(
        \u_outFIFO/n471 ) );
  OAI212 \u_outFIFO/U154  ( .A(\u_outFIFO/n396 ), .B(n782), .C(n1230), .Q(
        \u_outFIFO/n470 ) );
  OAI212 \u_outFIFO/U152  ( .A(\u_outFIFO/n396 ), .B(n780), .C(n1230), .Q(
        \u_outFIFO/n468 ) );
  OAI212 \u_outFIFO/U151  ( .A(\u_outFIFO/n391 ), .B(n788), .C(n1230), .Q(
        \u_outFIFO/n467 ) );
  OAI212 \u_outFIFO/U150  ( .A(\u_outFIFO/n391 ), .B(n785), .C(n1230), .Q(
        \u_outFIFO/n466 ) );
  OAI212 \u_outFIFO/U149  ( .A(\u_outFIFO/n391 ), .B(n782), .C(n1229), .Q(
        \u_outFIFO/n465 ) );
  OAI212 \u_outFIFO/U148  ( .A(\u_outFIFO/n391 ), .B(n780), .C(n1229), .Q(
        \u_outFIFO/n464 ) );
  OAI212 \u_outFIFO/U147  ( .A(\u_outFIFO/n386 ), .B(n788), .C(n1229), .Q(
        \u_outFIFO/n463 ) );
  OAI212 \u_outFIFO/U146  ( .A(\u_outFIFO/n386 ), .B(n785), .C(n1229), .Q(
        \u_outFIFO/n462 ) );
  OAI212 \u_outFIFO/U145  ( .A(\u_outFIFO/n386 ), .B(n782), .C(n1229), .Q(
        \u_outFIFO/n461 ) );
  OAI212 \u_outFIFO/U144  ( .A(\u_outFIFO/n386 ), .B(n780), .C(n1229), .Q(
        \u_outFIFO/n460 ) );
  OAI212 \u_outFIFO/U143  ( .A(n873), .B(n788), .C(n1229), .Q(\u_outFIFO/n459 ) );
  OAI212 \u_outFIFO/U142  ( .A(\u_outFIFO/n381 ), .B(n785), .C(n1229), .Q(
        \u_outFIFO/n458 ) );
  OAI212 \u_outFIFO/U141  ( .A(\u_outFIFO/n381 ), .B(n782), .C(n1229), .Q(
        \u_outFIFO/n457 ) );
  OAI212 \u_outFIFO/U140  ( .A(\u_outFIFO/n381 ), .B(n780), .C(n1229), .Q(
        \u_outFIFO/n456 ) );
  OAI212 \u_outFIFO/U139  ( .A(n871), .B(n788), .C(n1229), .Q(\u_outFIFO/n455 ) );
  OAI212 \u_outFIFO/U138  ( .A(n870), .B(n785), .C(n1229), .Q(\u_outFIFO/n454 ) );
  OAI212 \u_outFIFO/U137  ( .A(n871), .B(n782), .C(n1229), .Q(\u_outFIFO/n453 ) );
  OAI212 \u_outFIFO/U136  ( .A(n870), .B(n780), .C(n1229), .Q(\u_outFIFO/n452 ) );
  OAI212 \u_outFIFO/U135  ( .A(n868), .B(n788), .C(n1229), .Q(\u_outFIFO/n451 ) );
  OAI212 \u_outFIFO/U134  ( .A(n867), .B(n785), .C(n1229), .Q(\u_outFIFO/n450 ) );
  OAI212 \u_outFIFO/U133  ( .A(n868), .B(n782), .C(n1229), .Q(\u_outFIFO/n449 ) );
  OAI212 \u_outFIFO/U132  ( .A(n867), .B(n780), .C(n1229), .Q(\u_outFIFO/n448 ) );
  OAI212 \u_outFIFO/U131  ( .A(n865), .B(n790), .C(n1229), .Q(\u_outFIFO/n447 ) );
  OAI212 \u_outFIFO/U130  ( .A(n864), .B(n787), .C(n1229), .Q(\u_outFIFO/n446 ) );
  OAI212 \u_outFIFO/U129  ( .A(n865), .B(n784), .C(n1229), .Q(\u_outFIFO/n445 ) );
  OAI212 \u_outFIFO/U128  ( .A(n864), .B(n780), .C(n1229), .Q(\u_outFIFO/n444 ) );
  OAI212 \u_outFIFO/U127  ( .A(n862), .B(n789), .C(n1229), .Q(\u_outFIFO/n443 ) );
  OAI212 \u_outFIFO/U126  ( .A(n861), .B(n786), .C(n1229), .Q(\u_outFIFO/n442 ) );
  OAI212 \u_outFIFO/U125  ( .A(n862), .B(n783), .C(n1229), .Q(\u_outFIFO/n441 ) );
  OAI212 \u_outFIFO/U124  ( .A(n861), .B(n780), .C(n1229), .Q(\u_outFIFO/n440 ) );
  OAI212 \u_outFIFO/U123  ( .A(n859), .B(n790), .C(n1229), .Q(\u_outFIFO/n439 ) );
  OAI212 \u_outFIFO/U122  ( .A(n858), .B(n787), .C(n1228), .Q(\u_outFIFO/n438 ) );
  OAI212 \u_outFIFO/U121  ( .A(n859), .B(n784), .C(n1228), .Q(\u_outFIFO/n437 ) );
  OAI212 \u_outFIFO/U120  ( .A(n858), .B(n781), .C(n1228), .Q(\u_outFIFO/n436 ) );
  OAI212 \u_outFIFO/U119  ( .A(n856), .B(n789), .C(n1228), .Q(\u_outFIFO/n435 ) );
  OAI212 \u_outFIFO/U118  ( .A(n855), .B(n786), .C(n1228), .Q(\u_outFIFO/n434 ) );
  OAI212 \u_outFIFO/U117  ( .A(n856), .B(n783), .C(n1228), .Q(\u_outFIFO/n433 ) );
  OAI212 \u_outFIFO/U116  ( .A(n855), .B(n781), .C(n1228), .Q(\u_outFIFO/n432 ) );
  OAI212 \u_outFIFO/U115  ( .A(n853), .B(n790), .C(n1228), .Q(\u_outFIFO/n431 ) );
  OAI212 \u_outFIFO/U114  ( .A(n852), .B(n787), .C(n1228), .Q(\u_outFIFO/n430 ) );
  OAI212 \u_outFIFO/U113  ( .A(n853), .B(n784), .C(n1228), .Q(\u_outFIFO/n429 ) );
  OAI212 \u_outFIFO/U112  ( .A(n852), .B(n781), .C(n1228), .Q(\u_outFIFO/n428 ) );
  OAI212 \u_outFIFO/U111  ( .A(n850), .B(n789), .C(n1228), .Q(\u_outFIFO/n427 ) );
  OAI212 \u_outFIFO/U110  ( .A(n849), .B(n786), .C(n1228), .Q(\u_outFIFO/n426 ) );
  OAI212 \u_outFIFO/U109  ( .A(n850), .B(n783), .C(n1228), .Q(\u_outFIFO/n425 ) );
  OAI212 \u_outFIFO/U108  ( .A(n849), .B(n781), .C(n1228), .Q(\u_outFIFO/n424 ) );
  OAI212 \u_outFIFO/U107  ( .A(n844), .B(n790), .C(n1228), .Q(\u_outFIFO/n423 ) );
  OAI212 \u_outFIFO/U106  ( .A(n845), .B(n787), .C(n1228), .Q(\u_outFIFO/n422 ) );
  OAI212 \u_outFIFO/U105  ( .A(n846), .B(n784), .C(n1228), .Q(\u_outFIFO/n421 ) );
  OAI212 \u_outFIFO/U104  ( .A(n847), .B(n781), .C(n1228), .Q(\u_outFIFO/n420 ) );
  OAI212 \u_outFIFO/U103  ( .A(n842), .B(n789), .C(n1228), .Q(\u_outFIFO/n419 ) );
  OAI212 \u_outFIFO/U102  ( .A(\u_outFIFO/n331 ), .B(n786), .C(n1228), .Q(
        \u_outFIFO/n418 ) );
  OAI212 \u_outFIFO/U101  ( .A(\u_outFIFO/n331 ), .B(n783), .C(n1228), .Q(
        \u_outFIFO/n417 ) );
  OAI212 \u_outFIFO/U100  ( .A(\u_outFIFO/n331 ), .B(n781), .C(n1228), .Q(
        \u_outFIFO/n416 ) );
  OAI212 \u_outFIFO/U99  ( .A(n840), .B(n790), .C(n1228), .Q(\u_outFIFO/n415 )
         );
  OAI212 \u_outFIFO/U98  ( .A(n839), .B(n787), .C(n1228), .Q(\u_outFIFO/n414 )
         );
  OAI212 \u_outFIFO/U97  ( .A(n840), .B(n784), .C(n1228), .Q(\u_outFIFO/n413 )
         );
  OAI212 \u_outFIFO/U96  ( .A(n839), .B(n781), .C(n1227), .Q(\u_outFIFO/n412 )
         );
  OAI212 \u_outFIFO/U95  ( .A(\u_outFIFO/n317 ), .B(n789), .C(n1227), .Q(
        \u_outFIFO/n410 ) );
  OAI212 \u_outFIFO/U94  ( .A(\u_outFIFO/n317 ), .B(n786), .C(n1227), .Q(
        \u_outFIFO/n408 ) );
  OAI212 \u_outFIFO/U93  ( .A(\u_outFIFO/n317 ), .B(n783), .C(n1227), .Q(
        \u_outFIFO/n406 ) );
  OAI212 \u_outFIFO/U92  ( .A(n837), .B(n781), .C(n1227), .Q(\u_outFIFO/n404 )
         );
  OAI212 \u_outFIFO/U89  ( .A(\u_outFIFO/n324 ), .B(n889), .C(n1227), .Q(
        \u_outFIFO/n402 ) );
  OAI212 \u_outFIFO/U87  ( .A(\u_outFIFO/n322 ), .B(\u_outFIFO/n396 ), .C(
        n1227), .Q(\u_outFIFO/n400 ) );
  OAI212 \u_outFIFO/U85  ( .A(\u_outFIFO/n320 ), .B(\u_outFIFO/n396 ), .C(
        n1227), .Q(\u_outFIFO/n398 ) );
  OAI212 \u_outFIFO/U83  ( .A(\u_outFIFO/n318 ), .B(\u_outFIFO/n396 ), .C(
        n1227), .Q(\u_outFIFO/n395 ) );
  OAI212 \u_outFIFO/U82  ( .A(\u_outFIFO/n324 ), .B(n877), .C(n1227), .Q(
        \u_outFIFO/n394 ) );
  OAI212 \u_outFIFO/U81  ( .A(\u_outFIFO/n322 ), .B(\u_outFIFO/n391 ), .C(
        n1227), .Q(\u_outFIFO/n393 ) );
  OAI212 \u_outFIFO/U80  ( .A(\u_outFIFO/n320 ), .B(\u_outFIFO/n391 ), .C(
        n1227), .Q(\u_outFIFO/n392 ) );
  OAI212 \u_outFIFO/U79  ( .A(\u_outFIFO/n318 ), .B(\u_outFIFO/n391 ), .C(
        n1227), .Q(\u_outFIFO/n390 ) );
  OAI212 \u_outFIFO/U78  ( .A(\u_outFIFO/n324 ), .B(n875), .C(n1227), .Q(
        \u_outFIFO/n389 ) );
  OAI212 \u_outFIFO/U77  ( .A(\u_outFIFO/n322 ), .B(\u_outFIFO/n386 ), .C(
        n1227), .Q(\u_outFIFO/n388 ) );
  OAI212 \u_outFIFO/U76  ( .A(\u_outFIFO/n320 ), .B(\u_outFIFO/n386 ), .C(
        n1227), .Q(\u_outFIFO/n387 ) );
  OAI212 \u_outFIFO/U75  ( .A(\u_outFIFO/n318 ), .B(\u_outFIFO/n386 ), .C(
        n1227), .Q(\u_outFIFO/n385 ) );
  OAI212 \u_outFIFO/U74  ( .A(\u_outFIFO/n324 ), .B(\u_outFIFO/n381 ), .C(
        n1227), .Q(\u_outFIFO/n384 ) );
  OAI212 \u_outFIFO/U73  ( .A(\u_outFIFO/n322 ), .B(\u_outFIFO/n381 ), .C(
        n1227), .Q(\u_outFIFO/n383 ) );
  OAI212 \u_outFIFO/U72  ( .A(\u_outFIFO/n320 ), .B(\u_outFIFO/n381 ), .C(
        n1227), .Q(\u_outFIFO/n382 ) );
  OAI212 \u_outFIFO/U71  ( .A(\u_outFIFO/n318 ), .B(n873), .C(n1227), .Q(
        \u_outFIFO/n380 ) );
  OAI212 \u_outFIFO/U70  ( .A(\u_outFIFO/n324 ), .B(n869), .C(n1227), .Q(
        \u_outFIFO/n379 ) );
  OAI212 \u_outFIFO/U69  ( .A(\u_outFIFO/n322 ), .B(n869), .C(n1227), .Q(
        \u_outFIFO/n378 ) );
  OAI212 \u_outFIFO/U68  ( .A(\u_outFIFO/n320 ), .B(n869), .C(n1227), .Q(
        \u_outFIFO/n377 ) );
  OAI212 \u_outFIFO/U67  ( .A(\u_outFIFO/n318 ), .B(n869), .C(n1227), .Q(
        \u_outFIFO/n375 ) );
  OAI212 \u_outFIFO/U66  ( .A(\u_outFIFO/n324 ), .B(n866), .C(n1227), .Q(
        \u_outFIFO/n374 ) );
  OAI212 \u_outFIFO/U65  ( .A(\u_outFIFO/n322 ), .B(n866), .C(n1227), .Q(
        \u_outFIFO/n373 ) );
  OAI212 \u_outFIFO/U64  ( .A(\u_outFIFO/n320 ), .B(n866), .C(n1226), .Q(
        \u_outFIFO/n372 ) );
  OAI212 \u_outFIFO/U63  ( .A(\u_outFIFO/n318 ), .B(n866), .C(n1226), .Q(
        \u_outFIFO/n370 ) );
  OAI212 \u_outFIFO/U62  ( .A(\u_outFIFO/n324 ), .B(n863), .C(n1226), .Q(
        \u_outFIFO/n369 ) );
  OAI212 \u_outFIFO/U61  ( .A(\u_outFIFO/n322 ), .B(n863), .C(n1226), .Q(
        \u_outFIFO/n368 ) );
  OAI212 \u_outFIFO/U60  ( .A(\u_outFIFO/n320 ), .B(n863), .C(n1226), .Q(
        \u_outFIFO/n367 ) );
  OAI212 \u_outFIFO/U59  ( .A(\u_outFIFO/n318 ), .B(n863), .C(n1226), .Q(
        \u_outFIFO/n365 ) );
  OAI212 \u_outFIFO/U58  ( .A(\u_outFIFO/n324 ), .B(n860), .C(n1226), .Q(
        \u_outFIFO/n364 ) );
  OAI212 \u_outFIFO/U57  ( .A(\u_outFIFO/n322 ), .B(n860), .C(n1226), .Q(
        \u_outFIFO/n363 ) );
  OAI212 \u_outFIFO/U56  ( .A(\u_outFIFO/n320 ), .B(n860), .C(n1226), .Q(
        \u_outFIFO/n362 ) );
  OAI212 \u_outFIFO/U55  ( .A(\u_outFIFO/n318 ), .B(n860), .C(n1226), .Q(
        \u_outFIFO/n360 ) );
  OAI212 \u_outFIFO/U54  ( .A(\u_outFIFO/n324 ), .B(n857), .C(n1226), .Q(
        \u_outFIFO/n359 ) );
  OAI212 \u_outFIFO/U53  ( .A(\u_outFIFO/n322 ), .B(n857), .C(n1226), .Q(
        \u_outFIFO/n358 ) );
  OAI212 \u_outFIFO/U52  ( .A(\u_outFIFO/n320 ), .B(n857), .C(n1226), .Q(
        \u_outFIFO/n357 ) );
  OAI212 \u_outFIFO/U51  ( .A(\u_outFIFO/n318 ), .B(n857), .C(n1226), .Q(
        \u_outFIFO/n355 ) );
  OAI212 \u_outFIFO/U50  ( .A(\u_outFIFO/n324 ), .B(n854), .C(n1228), .Q(
        \u_outFIFO/n354 ) );
  OAI212 \u_outFIFO/U49  ( .A(\u_outFIFO/n322 ), .B(n854), .C(n1226), .Q(
        \u_outFIFO/n353 ) );
  OAI212 \u_outFIFO/U48  ( .A(\u_outFIFO/n320 ), .B(n854), .C(n1226), .Q(
        \u_outFIFO/n352 ) );
  OAI212 \u_outFIFO/U47  ( .A(\u_outFIFO/n318 ), .B(n854), .C(n1226), .Q(
        \u_outFIFO/n350 ) );
  OAI212 \u_outFIFO/U46  ( .A(\u_outFIFO/n324 ), .B(n851), .C(n1226), .Q(
        \u_outFIFO/n349 ) );
  OAI212 \u_outFIFO/U45  ( .A(\u_outFIFO/n322 ), .B(n851), .C(n1226), .Q(
        \u_outFIFO/n348 ) );
  OAI212 \u_outFIFO/U44  ( .A(\u_outFIFO/n320 ), .B(n851), .C(n1226), .Q(
        \u_outFIFO/n347 ) );
  OAI212 \u_outFIFO/U43  ( .A(\u_outFIFO/n318 ), .B(n851), .C(n1226), .Q(
        \u_outFIFO/n345 ) );
  OAI212 \u_outFIFO/U42  ( .A(\u_outFIFO/n324 ), .B(n848), .C(n1226), .Q(
        \u_outFIFO/n344 ) );
  OAI212 \u_outFIFO/U41  ( .A(\u_outFIFO/n322 ), .B(n848), .C(n1226), .Q(
        \u_outFIFO/n343 ) );
  OAI212 \u_outFIFO/U40  ( .A(\u_outFIFO/n320 ), .B(n848), .C(n1226), .Q(
        \u_outFIFO/n342 ) );
  OAI212 \u_outFIFO/U39  ( .A(\u_outFIFO/n318 ), .B(n848), .C(n1226), .Q(
        \u_outFIFO/n340 ) );
  OAI212 \u_outFIFO/U38  ( .A(\u_outFIFO/n324 ), .B(n844), .C(n1226), .Q(
        \u_outFIFO/n339 ) );
  OAI212 \u_outFIFO/U37  ( .A(\u_outFIFO/n322 ), .B(n845), .C(n1226), .Q(
        \u_outFIFO/n338 ) );
  OAI212 \u_outFIFO/U36  ( .A(\u_outFIFO/n320 ), .B(n846), .C(n1225), .Q(
        \u_outFIFO/n337 ) );
  OAI212 \u_outFIFO/U35  ( .A(\u_outFIFO/n318 ), .B(n847), .C(n1225), .Q(
        \u_outFIFO/n335 ) );
  OAI212 \u_outFIFO/U34  ( .A(\u_outFIFO/n324 ), .B(n842), .C(n1225), .Q(
        \u_outFIFO/n334 ) );
  OAI212 \u_outFIFO/U33  ( .A(\u_outFIFO/n322 ), .B(\u_outFIFO/n331 ), .C(
        n1225), .Q(\u_outFIFO/n333 ) );
  OAI212 \u_outFIFO/U32  ( .A(\u_outFIFO/n320 ), .B(\u_outFIFO/n331 ), .C(
        n1225), .Q(\u_outFIFO/n332 ) );
  OAI212 \u_outFIFO/U31  ( .A(\u_outFIFO/n318 ), .B(n842), .C(n1225), .Q(
        \u_outFIFO/n330 ) );
  OAI212 \u_outFIFO/U30  ( .A(\u_outFIFO/n324 ), .B(n838), .C(n1225), .Q(
        \u_outFIFO/n329 ) );
  OAI212 \u_outFIFO/U29  ( .A(\u_outFIFO/n322 ), .B(n838), .C(n1225), .Q(
        \u_outFIFO/n328 ) );
  OAI212 \u_outFIFO/U28  ( .A(\u_outFIFO/n320 ), .B(n838), .C(n1225), .Q(
        \u_outFIFO/n327 ) );
  OAI212 \u_outFIFO/U27  ( .A(\u_outFIFO/n318 ), .B(n838), .C(n1225), .Q(
        \u_outFIFO/n325 ) );
  OAI212 \u_outFIFO/U26  ( .A(n837), .B(\u_outFIFO/n324 ), .C(n1225), .Q(
        \u_outFIFO/n323 ) );
  OAI212 \u_outFIFO/U25  ( .A(\u_outFIFO/n317 ), .B(\u_outFIFO/n322 ), .C(
        n1225), .Q(\u_outFIFO/n321 ) );
  OAI212 \u_outFIFO/U24  ( .A(\u_outFIFO/n317 ), .B(\u_outFIFO/n320 ), .C(
        n1225), .Q(\u_outFIFO/n319 ) );
  OAI212 \u_outFIFO/U23  ( .A(n837), .B(\u_outFIFO/n318 ), .C(n1225), .Q(
        \u_outFIFO/n316 ) );
  OAI222 \u_mux8/U1  ( .A(\u_mux8/n3 ), .B(n2132), .C(in_MUX_inSEL6[1]), .D(
        \u_mux8/n4 ), .Q(sig_MUX_outMUX8) );
  OAI212 \u_decoder/iq_demod/U30  ( .A(\u_decoder/iq_demod/n59 ), .B(
        sig_DEMUX_outDEMUX1[0]), .C(n2398), .Q(\u_decoder/iq_demod/n71 ) );
  OAI212 \u_decoder/fir_filter/U900  ( .A(n1106), .B(n325), .C(
        \u_decoder/fir_filter/n1145 ), .Q(\u_decoder/fir_filter/n1447 ) );
  OAI212 \u_decoder/fir_filter/U898  ( .A(n1129), .B(n339), .C(
        \u_decoder/fir_filter/n1144 ), .Q(\u_decoder/fir_filter/n1446 ) );
  OAI212 \u_decoder/fir_filter/U896  ( .A(n1121), .B(n79), .C(
        \u_decoder/fir_filter/n1143 ), .Q(\u_decoder/fir_filter/n1445 ) );
  OAI212 \u_decoder/fir_filter/U894  ( .A(n1121), .B(n2291), .C(
        \u_decoder/fir_filter/n1142 ), .Q(\u_decoder/fir_filter/n1444 ) );
  OAI212 \u_decoder/fir_filter/U892  ( .A(n1121), .B(n132), .C(
        \u_decoder/fir_filter/n1141 ), .Q(\u_decoder/fir_filter/n1443 ) );
  OAI212 \u_decoder/fir_filter/U890  ( .A(n1121), .B(n343), .C(
        \u_decoder/fir_filter/n1140 ), .Q(\u_decoder/fir_filter/n1442 ) );
  OAI212 \u_decoder/fir_filter/U888  ( .A(n1121), .B(n2890), .C(
        \u_decoder/fir_filter/n1139 ), .Q(\u_decoder/fir_filter/n1441 ) );
  OAI212 \u_decoder/fir_filter/U886  ( .A(n1122), .B(
        \u_decoder/fir_filter/dp_cluster_0/r164/PROD1[4] ), .C(
        \u_decoder/fir_filter/n1138 ), .Q(\u_decoder/fir_filter/n1440 ) );
  OAI212 \u_decoder/fir_filter/U884  ( .A(n1122), .B(n2296), .C(
        \u_decoder/fir_filter/n1137 ), .Q(\u_decoder/fir_filter/n1439 ) );
  OAI212 \u_decoder/fir_filter/U882  ( .A(n1122), .B(n359), .C(
        \u_decoder/fir_filter/n1136 ), .Q(\u_decoder/fir_filter/n1438 ) );
  OAI212 \u_decoder/fir_filter/U880  ( .A(n1122), .B(n74), .C(
        \u_decoder/fir_filter/n1135 ), .Q(\u_decoder/fir_filter/n1437 ) );
  OAI212 \u_decoder/fir_filter/U878  ( .A(n1122), .B(n84), .C(
        \u_decoder/fir_filter/n1134 ), .Q(\u_decoder/fir_filter/n1436 ) );
  OAI212 \u_decoder/fir_filter/U869  ( .A(n1122), .B(n324), .C(
        \u_decoder/fir_filter/n1130 ), .Q(\u_decoder/fir_filter/n1432 ) );
  OAI212 \u_decoder/fir_filter/U867  ( .A(n1122), .B(n330), .C(
        \u_decoder/fir_filter/n1129 ), .Q(\u_decoder/fir_filter/n1431 ) );
  OAI212 \u_decoder/fir_filter/U865  ( .A(n1123), .B(n331), .C(
        \u_decoder/fir_filter/n1128 ), .Q(\u_decoder/fir_filter/n1430 ) );
  OAI212 \u_decoder/fir_filter/U863  ( .A(n1123), .B(n332), .C(
        \u_decoder/fir_filter/n1127 ), .Q(\u_decoder/fir_filter/n1429 ) );
  OAI212 \u_decoder/fir_filter/U861  ( .A(n1123), .B(n128), .C(
        \u_decoder/fir_filter/n1126 ), .Q(\u_decoder/fir_filter/n1428 ) );
  OAI212 \u_decoder/fir_filter/U859  ( .A(n1123), .B(n351), .C(
        \u_decoder/fir_filter/n1125 ), .Q(\u_decoder/fir_filter/n1427 ) );
  OAI212 \u_decoder/fir_filter/U857  ( .A(n1123), .B(n2904), .C(
        \u_decoder/fir_filter/n1124 ), .Q(\u_decoder/fir_filter/n1426 ) );
  OAI212 \u_decoder/fir_filter/U855  ( .A(n1123), .B(
        \u_decoder/fir_filter/dp_cluster_0/r165/PROD1[5] ), .C(
        \u_decoder/fir_filter/n1123 ), .Q(\u_decoder/fir_filter/n1425 ) );
  OAI212 \u_decoder/fir_filter/U853  ( .A(n1123), .B(n2244), .C(
        \u_decoder/fir_filter/n1122 ), .Q(\u_decoder/fir_filter/n1424 ) );
  OAI212 \u_decoder/fir_filter/U851  ( .A(n1124), .B(n355), .C(
        \u_decoder/fir_filter/n1121 ), .Q(\u_decoder/fir_filter/n1423 ) );
  OAI212 \u_decoder/fir_filter/U849  ( .A(n1124), .B(n89), .C(
        \u_decoder/fir_filter/n1120 ), .Q(\u_decoder/fir_filter/n1422 ) );
  OAI212 \u_decoder/fir_filter/U847  ( .A(n1124), .B(n74), .C(
        \u_decoder/fir_filter/n1119 ), .Q(\u_decoder/fir_filter/n1421 ) );
  OAI212 \u_decoder/fir_filter/U845  ( .A(n1124), .B(n84), .C(
        \u_decoder/fir_filter/n1118 ), .Q(\u_decoder/fir_filter/n1420 ) );
  OAI212 \u_decoder/fir_filter/U836  ( .A(n1124), .B(n361), .C(
        \u_decoder/fir_filter/n1114 ), .Q(\u_decoder/fir_filter/n1416 ) );
  OAI212 \u_decoder/fir_filter/U834  ( .A(n1124), .B(n323), .C(
        \u_decoder/fir_filter/n1113 ), .Q(\u_decoder/fir_filter/n1415 ) );
  OAI212 \u_decoder/fir_filter/U832  ( .A(n1124), .B(n329), .C(
        \u_decoder/fir_filter/n1112 ), .Q(\u_decoder/fir_filter/n1414 ) );
  OAI212 \u_decoder/fir_filter/U830  ( .A(n1125), .B(n337), .C(
        \u_decoder/fir_filter/n1111 ), .Q(\u_decoder/fir_filter/n1413 ) );
  OAI212 \u_decoder/fir_filter/U828  ( .A(n1125), .B(n2250), .C(
        \u_decoder/fir_filter/n1110 ), .Q(\u_decoder/fir_filter/n1412 ) );
  OAI212 \u_decoder/fir_filter/U826  ( .A(n1125), .B(n367), .C(
        \u_decoder/fir_filter/n1109 ), .Q(\u_decoder/fir_filter/n1411 ) );
  OAI212 \u_decoder/fir_filter/U824  ( .A(n1125), .B(n2252), .C(
        \u_decoder/fir_filter/n1108 ), .Q(\u_decoder/fir_filter/n1410 ) );
  OAI212 \u_decoder/fir_filter/U822  ( .A(n1125), .B(n2253), .C(
        \u_decoder/fir_filter/n1107 ), .Q(\u_decoder/fir_filter/n1409 ) );
  OAI212 \u_decoder/fir_filter/U820  ( .A(n1125), .B(n2254), .C(
        \u_decoder/fir_filter/n1106 ), .Q(\u_decoder/fir_filter/n1408 ) );
  OAI212 \u_decoder/fir_filter/U818  ( .A(n1125), .B(n353), .C(
        \u_decoder/fir_filter/n1105 ), .Q(\u_decoder/fir_filter/n1407 ) );
  OAI212 \u_decoder/fir_filter/U816  ( .A(n1126), .B(n74), .C(
        \u_decoder/fir_filter/n1104 ), .Q(\u_decoder/fir_filter/n1406 ) );
  OAI212 \u_decoder/fir_filter/U814  ( .A(n1126), .B(n84), .C(
        \u_decoder/fir_filter/n1103 ), .Q(\u_decoder/fir_filter/n1405 ) );
  OAI212 \u_decoder/fir_filter/U808  ( .A(n1126), .B(n68), .C(
        \u_decoder/fir_filter/n1100 ), .Q(\u_decoder/fir_filter/n1402 ) );
  OAI212 \u_decoder/fir_filter/U806  ( .A(n1126), .B(n345), .C(
        \u_decoder/fir_filter/n1099 ), .Q(\u_decoder/fir_filter/n1401 ) );
  OAI212 \u_decoder/fir_filter/U804  ( .A(n1126), .B(n70), .C(
        \u_decoder/fir_filter/n1098 ), .Q(\u_decoder/fir_filter/n1400 ) );
  OAI212 \u_decoder/fir_filter/U802  ( .A(n1126), .B(n77), .C(
        \u_decoder/fir_filter/n1097 ), .Q(\u_decoder/fir_filter/n1399 ) );
  OAI212 \u_decoder/fir_filter/U800  ( .A(n1126), .B(n2281), .C(
        \u_decoder/fir_filter/n1096 ), .Q(\u_decoder/fir_filter/n1398 ) );
  OAI212 \u_decoder/fir_filter/U798  ( .A(n1127), .B(n341), .C(
        \u_decoder/fir_filter/n1095 ), .Q(\u_decoder/fir_filter/n1397 ) );
  OAI212 \u_decoder/fir_filter/U796  ( .A(n1127), .B(n2283), .C(
        \u_decoder/fir_filter/n1094 ), .Q(\u_decoder/fir_filter/n1396 ) );
  OAI212 \u_decoder/fir_filter/U794  ( .A(n1127), .B(n369), .C(
        \u_decoder/fir_filter/n1093 ), .Q(\u_decoder/fir_filter/n1395 ) );
  OAI212 \u_decoder/fir_filter/U792  ( .A(n1127), .B(n2284), .C(
        \u_decoder/fir_filter/n1092 ), .Q(\u_decoder/fir_filter/n1394 ) );
  OAI212 \u_decoder/fir_filter/U790  ( .A(n1127), .B(n2285), .C(
        \u_decoder/fir_filter/n1091 ), .Q(\u_decoder/fir_filter/n1393 ) );
  OAI212 \u_decoder/fir_filter/U788  ( .A(n1127), .B(n2286), .C(
        \u_decoder/fir_filter/n1090 ), .Q(\u_decoder/fir_filter/n1392 ) );
  OAI212 \u_decoder/fir_filter/U786  ( .A(n1127), .B(n2287), .C(
        \u_decoder/fir_filter/n1089 ), .Q(\u_decoder/fir_filter/n1391 ) );
  OAI212 \u_decoder/fir_filter/U784  ( .A(n1128), .B(n2288), .C(
        \u_decoder/fir_filter/n1088 ), .Q(\u_decoder/fir_filter/n1390 ) );
  OAI212 \u_decoder/fir_filter/U782  ( .A(n1128), .B(n357), .C(
        \u_decoder/fir_filter/n1087 ), .Q(\u_decoder/fir_filter/n1389 ) );
  OAI212 \u_decoder/fir_filter/U780  ( .A(n1128), .B(n84), .C(
        \u_decoder/fir_filter/n1086 ), .Q(\u_decoder/fir_filter/n1388 ) );
  OAI212 \u_decoder/fir_filter/U760  ( .A(n1128), .B(n68), .C(
        \u_decoder/fir_filter/n1068 ), .Q(\u_decoder/fir_filter/n1386 ) );
  OAI212 \u_decoder/fir_filter/U758  ( .A(n1128), .B(n345), .C(
        \u_decoder/fir_filter/n1067 ), .Q(\u_decoder/fir_filter/n1385 ) );
  OAI212 \u_decoder/fir_filter/U756  ( .A(n1128), .B(n70), .C(
        \u_decoder/fir_filter/n1066 ), .Q(\u_decoder/fir_filter/n1384 ) );
  OAI212 \u_decoder/fir_filter/U754  ( .A(n1128), .B(n77), .C(
        \u_decoder/fir_filter/n1065 ), .Q(\u_decoder/fir_filter/n1383 ) );
  OAI212 \u_decoder/fir_filter/U752  ( .A(n1129), .B(n2281), .C(
        \u_decoder/fir_filter/n1064 ), .Q(\u_decoder/fir_filter/n1382 ) );
  OAI212 \u_decoder/fir_filter/U750  ( .A(n1129), .B(n341), .C(
        \u_decoder/fir_filter/n1063 ), .Q(\u_decoder/fir_filter/n1381 ) );
  OAI212 \u_decoder/fir_filter/U748  ( .A(n1129), .B(n2283), .C(
        \u_decoder/fir_filter/n1062 ), .Q(\u_decoder/fir_filter/n1380 ) );
  OAI212 \u_decoder/fir_filter/U746  ( .A(n1129), .B(n369), .C(
        \u_decoder/fir_filter/n1061 ), .Q(\u_decoder/fir_filter/n1379 ) );
  OAI212 \u_decoder/fir_filter/U744  ( .A(n1129), .B(n2284), .C(
        \u_decoder/fir_filter/n1060 ), .Q(\u_decoder/fir_filter/n1378 ) );
  OAI212 \u_decoder/fir_filter/U742  ( .A(n1129), .B(n2285), .C(
        \u_decoder/fir_filter/n1059 ), .Q(\u_decoder/fir_filter/n1377 ) );
  OAI212 \u_decoder/fir_filter/U740  ( .A(n1130), .B(n2286), .C(
        \u_decoder/fir_filter/n1058 ), .Q(\u_decoder/fir_filter/n1376 ) );
  OAI212 \u_decoder/fir_filter/U738  ( .A(n1130), .B(n2287), .C(
        \u_decoder/fir_filter/n1057 ), .Q(\u_decoder/fir_filter/n1375 ) );
  OAI212 \u_decoder/fir_filter/U736  ( .A(n1130), .B(n2288), .C(
        \u_decoder/fir_filter/n1056 ), .Q(\u_decoder/fir_filter/n1374 ) );
  OAI212 \u_decoder/fir_filter/U734  ( .A(n1130), .B(n357), .C(
        \u_decoder/fir_filter/n1055 ), .Q(\u_decoder/fir_filter/n1373 ) );
  OAI212 \u_decoder/fir_filter/U732  ( .A(n1130), .B(n84), .C(
        \u_decoder/fir_filter/n1054 ), .Q(\u_decoder/fir_filter/n1372 ) );
  OAI212 \u_decoder/fir_filter/U724  ( .A(n1130), .B(n361), .C(
        \u_decoder/fir_filter/n1049 ), .Q(\u_decoder/fir_filter/n1368 ) );
  OAI212 \u_decoder/fir_filter/U722  ( .A(n1130), .B(n323), .C(
        \u_decoder/fir_filter/n1048 ), .Q(\u_decoder/fir_filter/n1367 ) );
  OAI212 \u_decoder/fir_filter/U720  ( .A(n1131), .B(n329), .C(
        \u_decoder/fir_filter/n1047 ), .Q(\u_decoder/fir_filter/n1366 ) );
  OAI212 \u_decoder/fir_filter/U718  ( .A(n1131), .B(n337), .C(
        \u_decoder/fir_filter/n1046 ), .Q(\u_decoder/fir_filter/n1365 ) );
  OAI212 \u_decoder/fir_filter/U716  ( .A(n1131), .B(n2250), .C(
        \u_decoder/fir_filter/n1045 ), .Q(\u_decoder/fir_filter/n1364 ) );
  OAI212 \u_decoder/fir_filter/U714  ( .A(n1131), .B(n367), .C(
        \u_decoder/fir_filter/n1044 ), .Q(\u_decoder/fir_filter/n1363 ) );
  OAI212 \u_decoder/fir_filter/U712  ( .A(n1131), .B(n2252), .C(
        \u_decoder/fir_filter/n1043 ), .Q(\u_decoder/fir_filter/n1362 ) );
  OAI212 \u_decoder/fir_filter/U710  ( .A(n1131), .B(n2253), .C(
        \u_decoder/fir_filter/n1042 ), .Q(\u_decoder/fir_filter/n1361 ) );
  OAI212 \u_decoder/fir_filter/U708  ( .A(n1131), .B(n2254), .C(
        \u_decoder/fir_filter/n1041 ), .Q(\u_decoder/fir_filter/n1360 ) );
  OAI212 \u_decoder/fir_filter/U706  ( .A(n1132), .B(n353), .C(
        \u_decoder/fir_filter/n1040 ), .Q(\u_decoder/fir_filter/n1359 ) );
  OAI212 \u_decoder/fir_filter/U704  ( .A(n1132), .B(n74), .C(
        \u_decoder/fir_filter/n1039 ), .Q(\u_decoder/fir_filter/n1358 ) );
  OAI212 \u_decoder/fir_filter/U702  ( .A(n1132), .B(n84), .C(
        \u_decoder/fir_filter/n1038 ), .Q(\u_decoder/fir_filter/n1357 ) );
  OAI212 \u_decoder/fir_filter/U692  ( .A(n1132), .B(n324), .C(
        \u_decoder/fir_filter/n1032 ), .Q(\u_decoder/fir_filter/n1352 ) );
  OAI212 \u_decoder/fir_filter/U690  ( .A(n1132), .B(n330), .C(
        \u_decoder/fir_filter/n1031 ), .Q(\u_decoder/fir_filter/n1351 ) );
  OAI212 \u_decoder/fir_filter/U688  ( .A(n1132), .B(n331), .C(
        \u_decoder/fir_filter/n1030 ), .Q(\u_decoder/fir_filter/n1350 ) );
  OAI212 \u_decoder/fir_filter/U686  ( .A(n1132), .B(n332), .C(
        \u_decoder/fir_filter/n1029 ), .Q(\u_decoder/fir_filter/n1349 ) );
  OAI212 \u_decoder/fir_filter/U684  ( .A(n1133), .B(n128), .C(
        \u_decoder/fir_filter/n1028 ), .Q(\u_decoder/fir_filter/n1348 ) );
  OAI212 \u_decoder/fir_filter/U682  ( .A(n1133), .B(n351), .C(
        \u_decoder/fir_filter/n1027 ), .Q(\u_decoder/fir_filter/n1347 ) );
  OAI212 \u_decoder/fir_filter/U680  ( .A(n1133), .B(n2904), .C(
        \u_decoder/fir_filter/n1026 ), .Q(\u_decoder/fir_filter/n1346 ) );
  OAI212 \u_decoder/fir_filter/U678  ( .A(n1133), .B(
        \u_decoder/fir_filter/dp_cluster_0/r165/PROD1[5] ), .C(
        \u_decoder/fir_filter/n1025 ), .Q(\u_decoder/fir_filter/n1345 ) );
  OAI212 \u_decoder/fir_filter/U676  ( .A(n1133), .B(n2244), .C(
        \u_decoder/fir_filter/n1024 ), .Q(\u_decoder/fir_filter/n1344 ) );
  OAI212 \u_decoder/fir_filter/U674  ( .A(n1133), .B(n355), .C(
        \u_decoder/fir_filter/n1023 ), .Q(\u_decoder/fir_filter/n1343 ) );
  OAI212 \u_decoder/fir_filter/U672  ( .A(n1133), .B(n89), .C(
        \u_decoder/fir_filter/n1022 ), .Q(\u_decoder/fir_filter/n1342 ) );
  OAI212 \u_decoder/fir_filter/U670  ( .A(n1134), .B(n74), .C(
        \u_decoder/fir_filter/n1021 ), .Q(\u_decoder/fir_filter/n1341 ) );
  OAI212 \u_decoder/fir_filter/U668  ( .A(n1134), .B(n84), .C(
        \u_decoder/fir_filter/n1020 ), .Q(\u_decoder/fir_filter/n1340 ) );
  OAI212 \u_decoder/fir_filter/U666  ( .A(n1172), .B(
        \u_decoder/fir_filter/n412 ), .C(\u_decoder/fir_filter/n1019 ), .Q(
        \u_decoder/fir_filter/n1338 ) );
  OAI212 \u_decoder/fir_filter/U665  ( .A(n1172), .B(
        \u_decoder/fir_filter/n413 ), .C(\u_decoder/fir_filter/n1019 ), .Q(
        \u_decoder/fir_filter/n1337 ) );
  OAI212 \u_decoder/fir_filter/U664  ( .A(n1172), .B(
        \u_decoder/fir_filter/n414 ), .C(\u_decoder/fir_filter/n1019 ), .Q(
        \u_decoder/fir_filter/n1336 ) );
  OAI222 \u_decoder/fir_filter/U663  ( .A(n1173), .B(
        \u_decoder/fir_filter/n415 ), .C(n1106), .D(n325), .Q(
        \u_decoder/fir_filter/n1335 ) );
  OAI222 \u_decoder/fir_filter/U662  ( .A(n1173), .B(
        \u_decoder/fir_filter/n416 ), .C(n1105), .D(n339), .Q(
        \u_decoder/fir_filter/n1334 ) );
  OAI222 \u_decoder/fir_filter/U661  ( .A(n1173), .B(
        \u_decoder/fir_filter/n417 ), .C(n1106), .D(n79), .Q(
        \u_decoder/fir_filter/n1333 ) );
  OAI222 \u_decoder/fir_filter/U660  ( .A(n1173), .B(
        \u_decoder/fir_filter/n418 ), .C(n1106), .D(n2291), .Q(
        \u_decoder/fir_filter/n1332 ) );
  OAI222 \u_decoder/fir_filter/U659  ( .A(n1173), .B(
        \u_decoder/fir_filter/n419 ), .C(n1104), .D(n132), .Q(
        \u_decoder/fir_filter/n1331 ) );
  OAI222 \u_decoder/fir_filter/U658  ( .A(n1173), .B(
        \u_decoder/fir_filter/n420 ), .C(n1104), .D(n343), .Q(
        \u_decoder/fir_filter/n1330 ) );
  OAI222 \u_decoder/fir_filter/U657  ( .A(n1174), .B(
        \u_decoder/fir_filter/n421 ), .C(n1106), .D(n2890), .Q(
        \u_decoder/fir_filter/n1329 ) );
  OAI222 \u_decoder/fir_filter/U656  ( .A(n1174), .B(
        \u_decoder/fir_filter/n422 ), .C(n1104), .D(
        \u_decoder/fir_filter/dp_cluster_0/r164/PROD1[4] ), .Q(
        \u_decoder/fir_filter/n1328 ) );
  OAI222 \u_decoder/fir_filter/U655  ( .A(n1174), .B(
        \u_decoder/fir_filter/n423 ), .C(n1106), .D(n2296), .Q(
        \u_decoder/fir_filter/n1327 ) );
  OAI222 \u_decoder/fir_filter/U654  ( .A(n1174), .B(
        \u_decoder/fir_filter/n424 ), .C(n1103), .D(n359), .Q(
        \u_decoder/fir_filter/n1326 ) );
  OAI222 \u_decoder/fir_filter/U653  ( .A(n1174), .B(
        \u_decoder/fir_filter/n425 ), .C(n1104), .D(n74), .Q(
        \u_decoder/fir_filter/n1325 ) );
  OAI222 \u_decoder/fir_filter/U652  ( .A(n1174), .B(
        \u_decoder/fir_filter/n426 ), .C(n1105), .D(n84), .Q(
        \u_decoder/fir_filter/n1324 ) );
  OAI212 \u_decoder/fir_filter/U637  ( .A(n1134), .B(
        \u_decoder/fir_filter/n412 ), .C(\u_decoder/fir_filter/n1011 ), .Q(
        \u_decoder/fir_filter/n1317 ) );
  OAI212 \u_decoder/fir_filter/U635  ( .A(n1134), .B(
        \u_decoder/fir_filter/n413 ), .C(\u_decoder/fir_filter/n1010 ), .Q(
        \u_decoder/fir_filter/n1316 ) );
  OAI212 \u_decoder/fir_filter/U633  ( .A(n1134), .B(
        \u_decoder/fir_filter/n414 ), .C(\u_decoder/fir_filter/n1009 ), .Q(
        \u_decoder/fir_filter/n1315 ) );
  OAI212 \u_decoder/fir_filter/U631  ( .A(n1134), .B(
        \u_decoder/fir_filter/n415 ), .C(\u_decoder/fir_filter/n1008 ), .Q(
        \u_decoder/fir_filter/n1314 ) );
  OAI212 \u_decoder/fir_filter/U629  ( .A(n1134), .B(
        \u_decoder/fir_filter/n416 ), .C(\u_decoder/fir_filter/n1007 ), .Q(
        \u_decoder/fir_filter/n1313 ) );
  OAI212 \u_decoder/fir_filter/U627  ( .A(n1135), .B(
        \u_decoder/fir_filter/n417 ), .C(\u_decoder/fir_filter/n1006 ), .Q(
        \u_decoder/fir_filter/n1312 ) );
  OAI212 \u_decoder/fir_filter/U625  ( .A(n1135), .B(
        \u_decoder/fir_filter/n418 ), .C(\u_decoder/fir_filter/n1005 ), .Q(
        \u_decoder/fir_filter/n1311 ) );
  OAI212 \u_decoder/fir_filter/U623  ( .A(n1135), .B(
        \u_decoder/fir_filter/n419 ), .C(\u_decoder/fir_filter/n1004 ), .Q(
        \u_decoder/fir_filter/n1310 ) );
  OAI212 \u_decoder/fir_filter/U621  ( .A(n1135), .B(
        \u_decoder/fir_filter/n420 ), .C(\u_decoder/fir_filter/n1003 ), .Q(
        \u_decoder/fir_filter/n1309 ) );
  OAI212 \u_decoder/fir_filter/U619  ( .A(n1135), .B(
        \u_decoder/fir_filter/n421 ), .C(\u_decoder/fir_filter/n1002 ), .Q(
        \u_decoder/fir_filter/n1308 ) );
  OAI212 \u_decoder/fir_filter/U617  ( .A(n1135), .B(
        \u_decoder/fir_filter/n422 ), .C(\u_decoder/fir_filter/n1001 ), .Q(
        \u_decoder/fir_filter/n1307 ) );
  OAI212 \u_decoder/fir_filter/U615  ( .A(n1135), .B(
        \u_decoder/fir_filter/n423 ), .C(\u_decoder/fir_filter/n1000 ), .Q(
        \u_decoder/fir_filter/n1306 ) );
  OAI212 \u_decoder/fir_filter/U613  ( .A(n1136), .B(
        \u_decoder/fir_filter/n424 ), .C(\u_decoder/fir_filter/n999 ), .Q(
        \u_decoder/fir_filter/n1305 ) );
  OAI212 \u_decoder/fir_filter/U611  ( .A(n1136), .B(
        \u_decoder/fir_filter/n425 ), .C(\u_decoder/fir_filter/n998 ), .Q(
        \u_decoder/fir_filter/n1304 ) );
  OAI212 \u_decoder/fir_filter/U609  ( .A(n1136), .B(
        \u_decoder/fir_filter/n426 ), .C(\u_decoder/fir_filter/n997 ), .Q(
        \u_decoder/fir_filter/n1303 ) );
  OAI212 \u_decoder/fir_filter/U455  ( .A(n1136), .B(n328), .C(
        \u_decoder/fir_filter/n848 ), .Q(\u_decoder/fir_filter/n1299 ) );
  OAI212 \u_decoder/fir_filter/U453  ( .A(n1136), .B(n340), .C(
        \u_decoder/fir_filter/n847 ), .Q(\u_decoder/fir_filter/n1298 ) );
  OAI212 \u_decoder/fir_filter/U451  ( .A(n1136), .B(n78), .C(
        \u_decoder/fir_filter/n846 ), .Q(\u_decoder/fir_filter/n1297 ) );
  OAI212 \u_decoder/fir_filter/U449  ( .A(n1136), .B(n2362), .C(
        \u_decoder/fir_filter/n845 ), .Q(\u_decoder/fir_filter/n1296 ) );
  OAI212 \u_decoder/fir_filter/U447  ( .A(n1137), .B(n131), .C(
        \u_decoder/fir_filter/n844 ), .Q(\u_decoder/fir_filter/n1295 ) );
  OAI212 \u_decoder/fir_filter/U445  ( .A(n1137), .B(n344), .C(
        \u_decoder/fir_filter/n843 ), .Q(\u_decoder/fir_filter/n1294 ) );
  OAI212 \u_decoder/fir_filter/U443  ( .A(n1113), .B(n2804), .C(
        \u_decoder/fir_filter/n842 ), .Q(\u_decoder/fir_filter/n1293 ) );
  OAI212 \u_decoder/fir_filter/U441  ( .A(n1107), .B(
        \u_decoder/fir_filter/dp_cluster_0/r177/PROD1[4] ), .C(
        \u_decoder/fir_filter/n841 ), .Q(\u_decoder/fir_filter/n1292 ) );
  OAI212 \u_decoder/fir_filter/U439  ( .A(n1106), .B(n2367), .C(
        \u_decoder/fir_filter/n840 ), .Q(\u_decoder/fir_filter/n1291 ) );
  OAI212 \u_decoder/fir_filter/U437  ( .A(n1109), .B(n360), .C(
        \u_decoder/fir_filter/n839 ), .Q(\u_decoder/fir_filter/n1290 ) );
  OAI212 \u_decoder/fir_filter/U435  ( .A(n1109), .B(n75), .C(
        \u_decoder/fir_filter/n838 ), .Q(\u_decoder/fir_filter/n1289 ) );
  OAI212 \u_decoder/fir_filter/U433  ( .A(n1107), .B(n88), .C(
        \u_decoder/fir_filter/n837 ), .Q(\u_decoder/fir_filter/n1288 ) );
  OAI212 \u_decoder/fir_filter/U424  ( .A(n1107), .B(n327), .C(
        \u_decoder/fir_filter/n833 ), .Q(\u_decoder/fir_filter/n1284 ) );
  OAI212 \u_decoder/fir_filter/U422  ( .A(n1108), .B(n334), .C(
        \u_decoder/fir_filter/n832 ), .Q(\u_decoder/fir_filter/n1283 ) );
  OAI212 \u_decoder/fir_filter/U420  ( .A(n1107), .B(n335), .C(
        \u_decoder/fir_filter/n831 ), .Q(\u_decoder/fir_filter/n1282 ) );
  OAI212 \u_decoder/fir_filter/U418  ( .A(n1107), .B(n336), .C(
        \u_decoder/fir_filter/n830 ), .Q(\u_decoder/fir_filter/n1281 ) );
  OAI212 \u_decoder/fir_filter/U416  ( .A(n1108), .B(n127), .C(
        \u_decoder/fir_filter/n829 ), .Q(\u_decoder/fir_filter/n1280 ) );
  OAI212 \u_decoder/fir_filter/U414  ( .A(n1108), .B(n352), .C(
        \u_decoder/fir_filter/n828 ), .Q(\u_decoder/fir_filter/n1279 ) );
  OAI212 \u_decoder/fir_filter/U412  ( .A(n1107), .B(n2818), .C(
        \u_decoder/fir_filter/n827 ), .Q(\u_decoder/fir_filter/n1278 ) );
  OAI212 \u_decoder/fir_filter/U410  ( .A(n1108), .B(
        \u_decoder/fir_filter/dp_cluster_0/r178/PROD1[5] ), .C(
        \u_decoder/fir_filter/n826 ), .Q(\u_decoder/fir_filter/n1277 ) );
  OAI212 \u_decoder/fir_filter/U408  ( .A(n1107), .B(n2315), .C(
        \u_decoder/fir_filter/n825 ), .Q(\u_decoder/fir_filter/n1276 ) );
  OAI212 \u_decoder/fir_filter/U406  ( .A(n1108), .B(n356), .C(
        \u_decoder/fir_filter/n824 ), .Q(\u_decoder/fir_filter/n1275 ) );
  OAI212 \u_decoder/fir_filter/U404  ( .A(n1109), .B(n90), .C(
        \u_decoder/fir_filter/n823 ), .Q(\u_decoder/fir_filter/n1274 ) );
  OAI212 \u_decoder/fir_filter/U402  ( .A(n1108), .B(n75), .C(
        \u_decoder/fir_filter/n822 ), .Q(\u_decoder/fir_filter/n1273 ) );
  OAI212 \u_decoder/fir_filter/U400  ( .A(n1108), .B(n88), .C(
        \u_decoder/fir_filter/n821 ), .Q(\u_decoder/fir_filter/n1272 ) );
  OAI212 \u_decoder/fir_filter/U391  ( .A(n1109), .B(n362), .C(
        \u_decoder/fir_filter/n817 ), .Q(\u_decoder/fir_filter/n1268 ) );
  OAI212 \u_decoder/fir_filter/U389  ( .A(n1109), .B(n326), .C(
        \u_decoder/fir_filter/n816 ), .Q(\u_decoder/fir_filter/n1267 ) );
  OAI212 \u_decoder/fir_filter/U387  ( .A(n1109), .B(n333), .C(
        \u_decoder/fir_filter/n815 ), .Q(\u_decoder/fir_filter/n1266 ) );
  OAI212 \u_decoder/fir_filter/U385  ( .A(n1109), .B(n338), .C(
        \u_decoder/fir_filter/n814 ), .Q(\u_decoder/fir_filter/n1265 ) );
  OAI212 \u_decoder/fir_filter/U383  ( .A(n1110), .B(n2321), .C(
        \u_decoder/fir_filter/n813 ), .Q(\u_decoder/fir_filter/n1264 ) );
  OAI212 \u_decoder/fir_filter/U381  ( .A(n1110), .B(n368), .C(
        \u_decoder/fir_filter/n812 ), .Q(\u_decoder/fir_filter/n1263 ) );
  OAI212 \u_decoder/fir_filter/U379  ( .A(n1110), .B(n2323), .C(
        \u_decoder/fir_filter/n811 ), .Q(\u_decoder/fir_filter/n1262 ) );
  OAI212 \u_decoder/fir_filter/U377  ( .A(n1110), .B(n2324), .C(
        \u_decoder/fir_filter/n810 ), .Q(\u_decoder/fir_filter/n1261 ) );
  OAI212 \u_decoder/fir_filter/U375  ( .A(n1110), .B(n2325), .C(
        \u_decoder/fir_filter/n809 ), .Q(\u_decoder/fir_filter/n1260 ) );
  OAI212 \u_decoder/fir_filter/U373  ( .A(n1110), .B(n354), .C(
        \u_decoder/fir_filter/n808 ), .Q(\u_decoder/fir_filter/n1259 ) );
  OAI212 \u_decoder/fir_filter/U371  ( .A(n1110), .B(n75), .C(
        \u_decoder/fir_filter/n807 ), .Q(\u_decoder/fir_filter/n1258 ) );
  OAI212 \u_decoder/fir_filter/U369  ( .A(n1111), .B(n88), .C(
        \u_decoder/fir_filter/n806 ), .Q(\u_decoder/fir_filter/n1257 ) );
  OAI212 \u_decoder/fir_filter/U363  ( .A(n1111), .B(n67), .C(
        \u_decoder/fir_filter/n803 ), .Q(\u_decoder/fir_filter/n1254 ) );
  OAI212 \u_decoder/fir_filter/U361  ( .A(n1111), .B(n346), .C(
        \u_decoder/fir_filter/n802 ), .Q(\u_decoder/fir_filter/n1253 ) );
  OAI212 \u_decoder/fir_filter/U359  ( .A(n1111), .B(n69), .C(
        \u_decoder/fir_filter/n801 ), .Q(\u_decoder/fir_filter/n1252 ) );
  OAI212 \u_decoder/fir_filter/U357  ( .A(n1111), .B(n76), .C(
        \u_decoder/fir_filter/n800 ), .Q(\u_decoder/fir_filter/n1251 ) );
  OAI212 \u_decoder/fir_filter/U355  ( .A(n1111), .B(n2352), .C(
        \u_decoder/fir_filter/n799 ), .Q(\u_decoder/fir_filter/n1250 ) );
  OAI212 \u_decoder/fir_filter/U353  ( .A(n1111), .B(n342), .C(
        \u_decoder/fir_filter/n798 ), .Q(\u_decoder/fir_filter/n1249 ) );
  OAI212 \u_decoder/fir_filter/U351  ( .A(n1112), .B(n2354), .C(
        \u_decoder/fir_filter/n797 ), .Q(\u_decoder/fir_filter/n1248 ) );
  OAI212 \u_decoder/fir_filter/U349  ( .A(n1112), .B(n370), .C(
        \u_decoder/fir_filter/n796 ), .Q(\u_decoder/fir_filter/n1247 ) );
  OAI212 \u_decoder/fir_filter/U347  ( .A(n1112), .B(n2355), .C(
        \u_decoder/fir_filter/n795 ), .Q(\u_decoder/fir_filter/n1246 ) );
  OAI212 \u_decoder/fir_filter/U345  ( .A(n1112), .B(n2356), .C(
        \u_decoder/fir_filter/n794 ), .Q(\u_decoder/fir_filter/n1245 ) );
  OAI212 \u_decoder/fir_filter/U343  ( .A(n1112), .B(n2357), .C(
        \u_decoder/fir_filter/n793 ), .Q(\u_decoder/fir_filter/n1244 ) );
  OAI212 \u_decoder/fir_filter/U341  ( .A(n1112), .B(n2358), .C(
        \u_decoder/fir_filter/n792 ), .Q(\u_decoder/fir_filter/n1243 ) );
  OAI212 \u_decoder/fir_filter/U339  ( .A(n1112), .B(n2359), .C(
        \u_decoder/fir_filter/n791 ), .Q(\u_decoder/fir_filter/n1242 ) );
  OAI212 \u_decoder/fir_filter/U337  ( .A(n1113), .B(n358), .C(
        \u_decoder/fir_filter/n790 ), .Q(\u_decoder/fir_filter/n1241 ) );
  OAI212 \u_decoder/fir_filter/U335  ( .A(n1113), .B(n88), .C(
        \u_decoder/fir_filter/n789 ), .Q(\u_decoder/fir_filter/n1240 ) );
  OAI212 \u_decoder/fir_filter/U315  ( .A(n1113), .B(n67), .C(
        \u_decoder/fir_filter/n771 ), .Q(\u_decoder/fir_filter/n1238 ) );
  OAI212 \u_decoder/fir_filter/U313  ( .A(n1113), .B(n346), .C(
        \u_decoder/fir_filter/n770 ), .Q(\u_decoder/fir_filter/n1237 ) );
  OAI212 \u_decoder/fir_filter/U311  ( .A(n1113), .B(n69), .C(
        \u_decoder/fir_filter/n769 ), .Q(\u_decoder/fir_filter/n1236 ) );
  OAI212 \u_decoder/fir_filter/U309  ( .A(n1113), .B(n76), .C(
        \u_decoder/fir_filter/n768 ), .Q(\u_decoder/fir_filter/n1235 ) );
  OAI212 \u_decoder/fir_filter/U307  ( .A(n1114), .B(n2352), .C(
        \u_decoder/fir_filter/n767 ), .Q(\u_decoder/fir_filter/n1234 ) );
  OAI212 \u_decoder/fir_filter/U305  ( .A(n1114), .B(n342), .C(
        \u_decoder/fir_filter/n766 ), .Q(\u_decoder/fir_filter/n1233 ) );
  OAI212 \u_decoder/fir_filter/U303  ( .A(n1114), .B(n2354), .C(
        \u_decoder/fir_filter/n765 ), .Q(\u_decoder/fir_filter/n1232 ) );
  OAI212 \u_decoder/fir_filter/U301  ( .A(n1114), .B(n370), .C(
        \u_decoder/fir_filter/n764 ), .Q(\u_decoder/fir_filter/n1231 ) );
  OAI212 \u_decoder/fir_filter/U299  ( .A(n1114), .B(n2355), .C(
        \u_decoder/fir_filter/n763 ), .Q(\u_decoder/fir_filter/n1230 ) );
  OAI212 \u_decoder/fir_filter/U297  ( .A(n1114), .B(n2356), .C(
        \u_decoder/fir_filter/n762 ), .Q(\u_decoder/fir_filter/n1229 ) );
  OAI212 \u_decoder/fir_filter/U295  ( .A(n1114), .B(n2357), .C(
        \u_decoder/fir_filter/n761 ), .Q(\u_decoder/fir_filter/n1228 ) );
  OAI212 \u_decoder/fir_filter/U293  ( .A(n1115), .B(n2358), .C(
        \u_decoder/fir_filter/n760 ), .Q(\u_decoder/fir_filter/n1227 ) );
  OAI212 \u_decoder/fir_filter/U291  ( .A(n1115), .B(n2359), .C(
        \u_decoder/fir_filter/n759 ), .Q(\u_decoder/fir_filter/n1226 ) );
  OAI212 \u_decoder/fir_filter/U289  ( .A(n1115), .B(n358), .C(
        \u_decoder/fir_filter/n758 ), .Q(\u_decoder/fir_filter/n1225 ) );
  OAI212 \u_decoder/fir_filter/U287  ( .A(n1115), .B(n88), .C(
        \u_decoder/fir_filter/n757 ), .Q(\u_decoder/fir_filter/n1224 ) );
  OAI212 \u_decoder/fir_filter/U279  ( .A(n1115), .B(n362), .C(
        \u_decoder/fir_filter/n752 ), .Q(\u_decoder/fir_filter/n1220 ) );
  OAI212 \u_decoder/fir_filter/U277  ( .A(n1115), .B(n326), .C(
        \u_decoder/fir_filter/n751 ), .Q(\u_decoder/fir_filter/n1219 ) );
  OAI212 \u_decoder/fir_filter/U275  ( .A(n1115), .B(n333), .C(
        \u_decoder/fir_filter/n750 ), .Q(\u_decoder/fir_filter/n1218 ) );
  OAI212 \u_decoder/fir_filter/U273  ( .A(n1116), .B(n338), .C(
        \u_decoder/fir_filter/n749 ), .Q(\u_decoder/fir_filter/n1217 ) );
  OAI212 \u_decoder/fir_filter/U271  ( .A(n1116), .B(n2321), .C(
        \u_decoder/fir_filter/n748 ), .Q(\u_decoder/fir_filter/n1216 ) );
  OAI212 \u_decoder/fir_filter/U269  ( .A(n1116), .B(n368), .C(
        \u_decoder/fir_filter/n747 ), .Q(\u_decoder/fir_filter/n1215 ) );
  OAI212 \u_decoder/fir_filter/U267  ( .A(n1116), .B(n2323), .C(
        \u_decoder/fir_filter/n746 ), .Q(\u_decoder/fir_filter/n1214 ) );
  OAI212 \u_decoder/fir_filter/U265  ( .A(n1116), .B(n2324), .C(
        \u_decoder/fir_filter/n745 ), .Q(\u_decoder/fir_filter/n1213 ) );
  OAI212 \u_decoder/fir_filter/U263  ( .A(n1116), .B(n2325), .C(
        \u_decoder/fir_filter/n744 ), .Q(\u_decoder/fir_filter/n1212 ) );
  OAI212 \u_decoder/fir_filter/U261  ( .A(n1116), .B(n354), .C(
        \u_decoder/fir_filter/n743 ), .Q(\u_decoder/fir_filter/n1211 ) );
  OAI212 \u_decoder/fir_filter/U259  ( .A(n1117), .B(n75), .C(
        \u_decoder/fir_filter/n742 ), .Q(\u_decoder/fir_filter/n1210 ) );
  OAI212 \u_decoder/fir_filter/U257  ( .A(n1117), .B(n88), .C(
        \u_decoder/fir_filter/n741 ), .Q(\u_decoder/fir_filter/n1209 ) );
  OAI212 \u_decoder/fir_filter/U247  ( .A(n1117), .B(n327), .C(
        \u_decoder/fir_filter/n735 ), .Q(\u_decoder/fir_filter/n1204 ) );
  OAI212 \u_decoder/fir_filter/U245  ( .A(n1117), .B(n334), .C(
        \u_decoder/fir_filter/n734 ), .Q(\u_decoder/fir_filter/n1203 ) );
  OAI212 \u_decoder/fir_filter/U243  ( .A(n1117), .B(n335), .C(
        \u_decoder/fir_filter/n733 ), .Q(\u_decoder/fir_filter/n1202 ) );
  OAI212 \u_decoder/fir_filter/U241  ( .A(n1117), .B(n336), .C(
        \u_decoder/fir_filter/n732 ), .Q(\u_decoder/fir_filter/n1201 ) );
  OAI212 \u_decoder/fir_filter/U239  ( .A(n1117), .B(n127), .C(
        \u_decoder/fir_filter/n731 ), .Q(\u_decoder/fir_filter/n1200 ) );
  OAI212 \u_decoder/fir_filter/U237  ( .A(n1118), .B(n352), .C(
        \u_decoder/fir_filter/n730 ), .Q(\u_decoder/fir_filter/n1199 ) );
  OAI212 \u_decoder/fir_filter/U235  ( .A(n1118), .B(n2818), .C(
        \u_decoder/fir_filter/n729 ), .Q(\u_decoder/fir_filter/n1198 ) );
  OAI212 \u_decoder/fir_filter/U233  ( .A(n1118), .B(
        \u_decoder/fir_filter/dp_cluster_0/r178/PROD1[5] ), .C(
        \u_decoder/fir_filter/n728 ), .Q(\u_decoder/fir_filter/n1197 ) );
  OAI212 \u_decoder/fir_filter/U231  ( .A(n1118), .B(n2315), .C(
        \u_decoder/fir_filter/n727 ), .Q(\u_decoder/fir_filter/n1196 ) );
  OAI212 \u_decoder/fir_filter/U229  ( .A(n1118), .B(n356), .C(
        \u_decoder/fir_filter/n726 ), .Q(\u_decoder/fir_filter/n1195 ) );
  OAI212 \u_decoder/fir_filter/U227  ( .A(n1118), .B(n90), .C(
        \u_decoder/fir_filter/n725 ), .Q(\u_decoder/fir_filter/n1194 ) );
  OAI212 \u_decoder/fir_filter/U225  ( .A(n1118), .B(n75), .C(
        \u_decoder/fir_filter/n724 ), .Q(\u_decoder/fir_filter/n1193 ) );
  OAI212 \u_decoder/fir_filter/U223  ( .A(n1119), .B(n88), .C(
        \u_decoder/fir_filter/n723 ), .Q(\u_decoder/fir_filter/n1192 ) );
  OAI212 \u_decoder/fir_filter/U221  ( .A(n1173), .B(
        \u_decoder/fir_filter/n428 ), .C(\u_decoder/fir_filter/n722 ), .Q(
        \u_decoder/fir_filter/n1190 ) );
  OAI212 \u_decoder/fir_filter/U220  ( .A(n1173), .B(
        \u_decoder/fir_filter/n429 ), .C(\u_decoder/fir_filter/n722 ), .Q(
        \u_decoder/fir_filter/n1189 ) );
  OAI212 \u_decoder/fir_filter/U219  ( .A(n1173), .B(
        \u_decoder/fir_filter/n430 ), .C(\u_decoder/fir_filter/n722 ), .Q(
        \u_decoder/fir_filter/n1188 ) );
  OAI222 \u_decoder/fir_filter/U218  ( .A(n1174), .B(
        \u_decoder/fir_filter/n431 ), .C(n1105), .D(n328), .Q(
        \u_decoder/fir_filter/n1187 ) );
  OAI222 \u_decoder/fir_filter/U217  ( .A(n1174), .B(
        \u_decoder/fir_filter/n432 ), .C(n1104), .D(n340), .Q(
        \u_decoder/fir_filter/n1186 ) );
  OAI222 \u_decoder/fir_filter/U216  ( .A(n1174), .B(
        \u_decoder/fir_filter/n433 ), .C(n1105), .D(n78), .Q(
        \u_decoder/fir_filter/n1185 ) );
  OAI222 \u_decoder/fir_filter/U215  ( .A(n1174), .B(
        \u_decoder/fir_filter/n434 ), .C(n1105), .D(n2362), .Q(
        \u_decoder/fir_filter/n1184 ) );
  OAI222 \u_decoder/fir_filter/U214  ( .A(n1175), .B(
        \u_decoder/fir_filter/n435 ), .C(n1103), .D(n131), .Q(
        \u_decoder/fir_filter/n1183 ) );
  OAI222 \u_decoder/fir_filter/U213  ( .A(n1175), .B(
        \u_decoder/fir_filter/n436 ), .C(n1105), .D(n344), .Q(
        \u_decoder/fir_filter/n1182 ) );
  OAI222 \u_decoder/fir_filter/U212  ( .A(n1175), .B(
        \u_decoder/fir_filter/n437 ), .C(n1105), .D(n2804), .Q(
        \u_decoder/fir_filter/n1181 ) );
  OAI222 \u_decoder/fir_filter/U211  ( .A(n1175), .B(
        \u_decoder/fir_filter/n438 ), .C(n1103), .D(
        \u_decoder/fir_filter/dp_cluster_0/r177/PROD1[4] ), .Q(
        \u_decoder/fir_filter/n1180 ) );
  OAI222 \u_decoder/fir_filter/U210  ( .A(n1175), .B(
        \u_decoder/fir_filter/n439 ), .C(n1103), .D(n2367), .Q(
        \u_decoder/fir_filter/n1179 ) );
  OAI222 \u_decoder/fir_filter/U209  ( .A(n1175), .B(
        \u_decoder/fir_filter/n440 ), .C(n1104), .D(n360), .Q(
        \u_decoder/fir_filter/n1178 ) );
  OAI222 \u_decoder/fir_filter/U208  ( .A(n1175), .B(
        \u_decoder/fir_filter/n441 ), .C(n1103), .D(n75), .Q(
        \u_decoder/fir_filter/n1177 ) );
  OAI222 \u_decoder/fir_filter/U207  ( .A(n1175), .B(
        \u_decoder/fir_filter/n442 ), .C(n1104), .D(n88), .Q(
        \u_decoder/fir_filter/n1176 ) );
  OAI212 \u_decoder/fir_filter/U192  ( .A(n1119), .B(
        \u_decoder/fir_filter/n428 ), .C(\u_decoder/fir_filter/n713 ), .Q(
        \u_decoder/fir_filter/n1169 ) );
  OAI212 \u_decoder/fir_filter/U190  ( .A(n1119), .B(
        \u_decoder/fir_filter/n429 ), .C(\u_decoder/fir_filter/n712 ), .Q(
        \u_decoder/fir_filter/n1168 ) );
  OAI212 \u_decoder/fir_filter/U188  ( .A(n1119), .B(
        \u_decoder/fir_filter/n430 ), .C(\u_decoder/fir_filter/n711 ), .Q(
        \u_decoder/fir_filter/n1167 ) );
  OAI212 \u_decoder/fir_filter/U186  ( .A(n1119), .B(
        \u_decoder/fir_filter/n431 ), .C(\u_decoder/fir_filter/n710 ), .Q(
        \u_decoder/fir_filter/n1166 ) );
  OAI212 \u_decoder/fir_filter/U184  ( .A(n1119), .B(
        \u_decoder/fir_filter/n432 ), .C(\u_decoder/fir_filter/n709 ), .Q(
        \u_decoder/fir_filter/n1165 ) );
  OAI212 \u_decoder/fir_filter/U182  ( .A(n1119), .B(
        \u_decoder/fir_filter/n433 ), .C(\u_decoder/fir_filter/n708 ), .Q(
        \u_decoder/fir_filter/n1164 ) );
  OAI212 \u_decoder/fir_filter/U180  ( .A(n1120), .B(
        \u_decoder/fir_filter/n434 ), .C(\u_decoder/fir_filter/n707 ), .Q(
        \u_decoder/fir_filter/n1163 ) );
  OAI212 \u_decoder/fir_filter/U178  ( .A(n1120), .B(
        \u_decoder/fir_filter/n435 ), .C(\u_decoder/fir_filter/n706 ), .Q(
        \u_decoder/fir_filter/n1162 ) );
  OAI212 \u_decoder/fir_filter/U176  ( .A(n1120), .B(
        \u_decoder/fir_filter/n436 ), .C(\u_decoder/fir_filter/n705 ), .Q(
        \u_decoder/fir_filter/n1161 ) );
  OAI212 \u_decoder/fir_filter/U174  ( .A(n1120), .B(
        \u_decoder/fir_filter/n437 ), .C(\u_decoder/fir_filter/n704 ), .Q(
        \u_decoder/fir_filter/n1160 ) );
  OAI212 \u_decoder/fir_filter/U172  ( .A(n1120), .B(
        \u_decoder/fir_filter/n438 ), .C(\u_decoder/fir_filter/n703 ), .Q(
        \u_decoder/fir_filter/n1159 ) );
  OAI212 \u_decoder/fir_filter/U170  ( .A(n1120), .B(
        \u_decoder/fir_filter/n439 ), .C(\u_decoder/fir_filter/n702 ), .Q(
        \u_decoder/fir_filter/n1158 ) );
  OAI212 \u_decoder/fir_filter/U168  ( .A(n1120), .B(
        \u_decoder/fir_filter/n440 ), .C(\u_decoder/fir_filter/n701 ), .Q(
        \u_decoder/fir_filter/n1157 ) );
  OAI212 \u_decoder/fir_filter/U166  ( .A(n1121), .B(
        \u_decoder/fir_filter/n441 ), .C(\u_decoder/fir_filter/n700 ), .Q(
        \u_decoder/fir_filter/n1156 ) );
  OAI212 \u_decoder/fir_filter/U164  ( .A(n1121), .B(
        \u_decoder/fir_filter/n442 ), .C(\u_decoder/fir_filter/n699 ), .Q(
        \u_decoder/fir_filter/n1155 ) );
  OAI212 \u_cdr/phd1/U11  ( .A(\u_cdr/phd1/n19 ), .B(\u_cdr/phd1/n17 ), .C(
        \u_cdr/phd1/n20 ), .Q(\u_cdr/phd1/n23 ) );
  OAI212 \u_cdr/phd1/U8  ( .A(\u_cdr/phd1/n16 ), .B(\u_cdr/phd1/n17 ), .C(
        \u_cdr/phd1/n18 ), .Q(\u_cdr/phd1/n22 ) );
  OAI222 \u_cdr/dec1/U9  ( .A(n306), .B(\u_cdr/dir ), .C(\u_cdr/dec1/n20 ), 
        .D(\u_cdr/dec1/w_en_dec ), .Q(\u_cdr/dec1/n25 ) );
  OAI212 \u_decoder/iq_demod/cossin_dig/U31  ( .A(
        \u_decoder/iq_demod/cossin_dig/n47 ), .B(
        \u_decoder/iq_demod/cossin_dig/N20 ), .C(
        \u_decoder/iq_demod/cossin_dig/counter [2]), .Q(
        \u_decoder/iq_demod/cossin_dig/n46 ) );
  OAI222 \u_decoder/iq_demod/cossin_dig/U20  ( .A(
        \u_decoder/iq_demod/cossin_dig/n21 ), .B(
        \u_decoder/iq_demod/cossin_dig/n41 ), .C(
        \u_decoder/iq_demod/cossin_dig/N55 ), .D(
        \u_decoder/iq_demod/cossin_dig/n40 ), .Q(
        \u_decoder/iq_demod/cossin_dig/n53 ) );
  OAI222 \u_decoder/iq_demod/cossin_dig/U18  ( .A(
        \u_decoder/iq_demod/cossin_dig/n19 ), .B(n1845), .C(
        \u_decoder/iq_demod/cossin_dig/n21 ), .D(
        \u_decoder/iq_demod/cossin_dig/n40 ), .Q(
        \u_decoder/iq_demod/cossin_dig/n52 ) );
  OAI212 \u_decoder/iq_demod/cossin_dig/U10  ( .A(
        \u_decoder/iq_demod/cossin_dig/N55 ), .B(
        \u_decoder/iq_demod/cossin_dig/n31 ), .C(
        \u_decoder/iq_demod/cossin_dig/n32 ), .Q(
        \u_decoder/iq_demod/cossin_dig/n51 ) );
  OAI222 \u_mux7/mux3/U1  ( .A(n3110), .B(n2132), .C(in_MUX_inSEL6[1]), .D(
        n3111), .Q(sig_MUX_outMUX7[3]) );
  OAI222 \u_mux7/mux2/U1  ( .A(n3108), .B(n2132), .C(in_MUX_inSEL6[1]), .D(
        n3109), .Q(sig_MUX_outMUX7[2]) );
  OAI222 \u_mux7/mux1/U1  ( .A(n3106), .B(n2132), .C(in_MUX_inSEL6[1]), .D(
        n3107), .Q(sig_MUX_outMUX7[1]) );
  OAI222 \u_mux7/mux0/U1  ( .A(n3104), .B(n2132), .C(in_MUX_inSEL6[1]), .D(
        n3105), .Q(sig_MUX_outMUX7[0]) );
  OAI222 \u_mux6/mux3/U1  ( .A(n3102), .B(n2132), .C(in_MUX_inSEL6[1]), .D(
        n3103), .Q(sig_MUX_outMUX6[3]) );
  OAI222 \u_mux6/mux2/U1  ( .A(n3100), .B(n2132), .C(in_MUX_inSEL6[1]), .D(
        n3101), .Q(sig_MUX_outMUX6[2]) );
  OAI222 \u_mux6/mux1/U1  ( .A(n3098), .B(n2132), .C(in_MUX_inSEL6[1]), .D(
        n3099), .Q(sig_MUX_outMUX6[1]) );
  OAI222 \u_mux6/mux0/U1  ( .A(n3096), .B(n2132), .C(in_MUX_inSEL6[1]), .D(
        n3097), .Q(sig_MUX_outMUX6[0]) );
  OAI222 \u_mux10/mux3/U1  ( .A(n3094), .B(n2134), .C(in_MUX_inSEL9[1]), .D(
        n3095), .Q(out_MUX_outMUX10[3]) );
  OAI222 \u_mux10/mux2/U1  ( .A(n3092), .B(n2134), .C(in_MUX_inSEL9[1]), .D(
        n3093), .Q(out_MUX_outMUX10[2]) );
  OAI222 \u_mux10/mux1/U1  ( .A(n3090), .B(n2134), .C(in_MUX_inSEL9[1]), .D(
        n3091), .Q(out_MUX_outMUX10[1]) );
  OAI222 \u_mux10/mux0/U1  ( .A(n3088), .B(n2134), .C(in_MUX_inSEL9[1]), .D(
        n3089), .Q(out_MUX_outMUX10[0]) );
  OAI222 \u_mux9/mux3/U1  ( .A(n3086), .B(n2134), .C(in_MUX_inSEL9[1]), .D(
        n3087), .Q(out_MUX_outMUX9[3]) );
  OAI222 \u_mux9/mux2/U1  ( .A(n3084), .B(n2134), .C(in_MUX_inSEL9[1]), .D(
        n3085), .Q(out_MUX_outMUX9[2]) );
  OAI222 \u_mux9/mux1/U1  ( .A(n3082), .B(n2134), .C(in_MUX_inSEL9[1]), .D(
        n3083), .Q(out_MUX_outMUX9[1]) );
  OAI222 \u_mux9/mux0/U1  ( .A(n3080), .B(n2134), .C(in_MUX_inSEL9[1]), .D(
        n3081), .Q(out_MUX_outMUX9[0]) );
  OAI222 \u_mux16/U1  ( .A(n3078), .B(n2138), .C(in_MUX_inSEL15[1]), .D(n3079), 
        .Q(out_MUX_outMUX16) );
  OAI222 \u_mux15/U1  ( .A(n3076), .B(n2138), .C(in_MUX_inSEL15[1]), .D(n3077), 
        .Q(out_MUX_outMUX15) );
  ADD22 \u_cdr/phd1/cnt_phd/add_58/U1_1_1  ( .A(\u_cdr/phd1/cnt_phd/cnt [1]), 
        .B(\u_cdr/phd1/cnt_phd/cnt [0]), .CO(
        \u_cdr/phd1/cnt_phd/add_58/carry [2]), .S(\u_cdr/phd1/cnt_phd/N72 ) );
  ADD22 \u_cdr/phd1/cnt_phd/add_58/U1_1_2  ( .A(\u_cdr/phd1/cnt_phd/cnt [2]), 
        .B(\u_cdr/phd1/cnt_phd/add_58/carry [2]), .CO(
        \u_cdr/phd1/cnt_phd/add_58/carry [3]), .S(\u_cdr/phd1/cnt_phd/N73 ) );
  ADD22 \u_cdr/phd1/cnt_phd/add_58/U1_1_3  ( .A(\u_cdr/phd1/cnt_phd/cnt [3]), 
        .B(\u_cdr/phd1/cnt_phd/add_58/carry [3]), .CO(
        \u_cdr/phd1/cnt_phd/add_58/carry [4]), .S(\u_cdr/phd1/cnt_phd/N74 ) );
  ADD22 \u_cdr/phd1/cnt_phd/add_58/U1_1_4  ( .A(\u_cdr/phd1/cnt_phd/cnt [4]), 
        .B(\u_cdr/phd1/cnt_phd/add_58/carry [4]), .CO(
        \u_cdr/phd1/cnt_phd/add_58/carry [5]), .S(\u_cdr/phd1/cnt_phd/N75 ) );
  ADD22 \u_cdr/dec1/cnt_dec/add_20/U1_1_1  ( .A(
        \u_cdr/dec1/cnt_dec/cnt_dec [1]), .B(\u_cdr/dec1/cnt_dec/cnt_dec [0]), 
        .CO(\u_cdr/dec1/cnt_dec/add_20/carry [2]), .S(\u_cdr/dec1/cnt_dec/N5 )
         );
  ADD22 \u_cdr/dec1/cnt_dec/add_20/U1_1_2  ( .A(
        \u_cdr/dec1/cnt_dec/cnt_dec [2]), .B(
        \u_cdr/dec1/cnt_dec/add_20/carry [2]), .CO(
        \u_cdr/dec1/cnt_dec/add_20/carry [3]), .S(\u_cdr/dec1/cnt_dec/N6 ) );
  ADD22 \u_cdr/dec1/cnt_dec/add_20/U1_1_3  ( .A(
        \u_cdr/dec1/cnt_dec/cnt_dec [3]), .B(
        \u_cdr/dec1/cnt_dec/add_20/carry [3]), .CO(
        \u_cdr/dec1/cnt_dec/add_20/carry [4]), .S(\u_cdr/dec1/cnt_dec/N7 ) );
  ADD22 \u_cdr/dec1/cnt_dec/add_20/U1_1_4  ( .A(
        \u_cdr/dec1/cnt_dec/cnt_dec [4]), .B(
        \u_cdr/dec1/cnt_dec/add_20/carry [4]), .CO(
        \u_cdr/dec1/cnt_dec/add_20/carry [5]), .S(\u_cdr/dec1/cnt_dec/N8 ) );
  ADD22 \u_cdr/div1/cnt_div/add_58/U1_1_1  ( .A(\u_cdr/div1/cnt_div/cnt [1]), 
        .B(\u_cdr/div1/cnt_div/cnt [0]), .CO(
        \u_cdr/div1/cnt_div/add_58/carry [2]), .S(\u_cdr/div1/cnt_div/N72 ) );
  ADD22 \u_cdr/div1/cnt_div/add_58/U1_1_2  ( .A(\u_cdr/div1/cnt_div/cnt [2]), 
        .B(\u_cdr/div1/cnt_div/add_58/carry [2]), .CO(
        \u_cdr/div1/cnt_div/add_58/carry [3]), .S(\u_cdr/div1/cnt_div/N73 ) );
  ADD22 \u_cdr/div1/cnt_div/add_58/U1_1_3  ( .A(\u_cdr/div1/cnt_div/cnt [3]), 
        .B(\u_cdr/div1/cnt_div/add_58/carry [3]), .CO(
        \u_cdr/div1/cnt_div/add_58/carry [4]), .S(\u_cdr/div1/cnt_div/N74 ) );
  ADD22 \u_cdr/div1/cnt_div/add_58/U1_1_4  ( .A(\u_cdr/div1/cnt_div/cnt [4]), 
        .B(\u_cdr/div1/cnt_div/add_58/carry [4]), .CO(
        \u_cdr/div1/cnt_div/add_58/carry [5]), .S(\u_cdr/div1/cnt_div/N75 ) );
  ADD22 \u_cdr/dec1/add_40/U1_1_1  ( .A(\u_cdr/dec1/cnt_r [1]), .B(
        \u_cdr/dec1/cnt_r [0]), .CO(\u_cdr/dec1/add_40/carry [2]), .S(
        \u_cdr/dec1/N61 ) );
  ADD22 \u_cdr/dec1/add_40/U1_1_2  ( .A(\u_cdr/dec1/cnt_r [2]), .B(
        \u_cdr/dec1/add_40/carry [2]), .CO(\u_cdr/dec1/add_40/carry [3]), .S(
        \u_cdr/dec1/N62 ) );
  ADD22 \u_cdr/dec1/add_40/U1_1_3  ( .A(\u_cdr/dec1/cnt_r [3]), .B(
        \u_cdr/dec1/add_40/carry [3]), .CO(\u_cdr/dec1/add_40/carry [4]), .S(
        \u_cdr/dec1/N63 ) );
  ADD22 \u_cdr/dec1/add_40/U1_1_4  ( .A(\u_cdr/dec1/cnt_r [4]), .B(
        \u_cdr/dec1/add_40/carry [4]), .CO(\u_cdr/dec1/add_40/carry [5]), .S(
        \u_cdr/dec1/N64 ) );
  ADD32 \u_cordic/my_rotation/sub_35/U2_1  ( .A(
        \u_cordic/my_rotation/present_angle[0][1] ), .B(n64), .CI(
        \u_cordic/my_rotation/sub_35/carry [1]), .CO(
        \u_cordic/my_rotation/sub_35/carry [2]), .S(
        \u_cordic/my_rotation/delta [1]) );
  ADD32 \u_cordic/my_rotation/sub_35/U2_2  ( .A(
        \u_cordic/my_rotation/present_angle[0][2] ), .B(n63), .CI(
        \u_cordic/my_rotation/sub_35/carry [2]), .CO(
        \u_cordic/my_rotation/sub_35/carry [3]), .S(
        \u_cordic/my_rotation/delta [2]) );
  ADD32 \u_cordic/my_rotation/sub_35/U2_3  ( .A(
        \u_cordic/my_rotation/present_angle[0][3] ), .B(n21), .CI(
        \u_cordic/my_rotation/sub_35/carry [3]), .CO(
        \u_cordic/my_rotation/sub_35/carry [4]), .S(
        \u_cordic/my_rotation/delta [3]) );
  ADD32 \u_cordic/my_rotation/sub_35/U2_4  ( .A(
        \u_cordic/my_rotation/present_angle[0][4] ), .B(n66), .CI(
        \u_cordic/my_rotation/sub_35/carry [4]), .CO(
        \u_cordic/my_rotation/sub_35/carry [5]), .S(
        \u_cordic/my_rotation/delta [4]) );
  ADD32 \u_cordic/my_rotation/sub_35/U2_5  ( .A(
        \u_cordic/my_rotation/present_angle[0][5] ), .B(n73), .CI(
        \u_cordic/my_rotation/sub_35/carry [5]), .CO(
        \u_cordic/my_rotation/sub_35/carry [6]), .S(
        \u_cordic/my_rotation/delta [5]) );
  ADD32 \u_cordic/my_rotation/sub_35/U2_6  ( .A(
        \u_cordic/my_rotation/present_angle[0][6] ), .B(n72), .CI(
        \u_cordic/my_rotation/sub_35/carry [6]), .CO(
        \u_cordic/my_rotation/sub_35/carry [7]), .S(
        \u_cordic/my_rotation/delta [6]) );
  ADD32 \u_cordic/my_rotation/sub_35/U2_7  ( .A(
        \u_cordic/my_rotation/present_angle[0][7] ), .B(n71), .CI(
        \u_cordic/my_rotation/sub_35/carry [7]), .CO(
        \u_cordic/my_rotation/sub_35/carry [8]), .S(
        \u_cordic/my_rotation/delta [7]) );
  ADD32 \u_cordic/my_rotation/sub_35/U2_8  ( .A(
        \u_cordic/my_rotation/present_angle[0][8] ), .B(n87), .CI(
        \u_cordic/my_rotation/sub_35/carry [8]), .CO(
        \u_cordic/my_rotation/sub_35/carry [9]), .S(
        \u_cordic/my_rotation/delta [8]) );
  ADD32 \u_cordic/my_rotation/sub_35/U2_9  ( .A(
        \u_cordic/my_rotation/present_angle[0][9] ), .B(n86), .CI(
        \u_cordic/my_rotation/sub_35/carry [9]), .CO(
        \u_cordic/my_rotation/sub_35/carry [10]), .S(
        \u_cordic/my_rotation/delta [9]) );
  ADD32 \u_cordic/my_rotation/sub_35/U2_10  ( .A(
        \u_cordic/my_rotation/present_angle[0][10] ), .B(n85), .CI(
        \u_cordic/my_rotation/sub_35/carry [10]), .CO(
        \u_cordic/my_rotation/sub_35/carry [11]), .S(
        \u_cordic/my_rotation/delta [10]) );
  ADD32 \u_cordic/my_rotation/sub_35/U2_11  ( .A(
        \u_cordic/my_rotation/present_angle[0][11] ), .B(n134), .CI(
        \u_cordic/my_rotation/sub_35/carry [11]), .CO(
        \u_cordic/my_rotation/sub_35/carry [12]), .S(
        \u_cordic/my_rotation/delta [11]) );
  ADD32 \u_cordic/my_rotation/sub_35/U2_12  ( .A(
        \u_cordic/my_rotation/present_angle[0][12] ), .B(n133), .CI(
        \u_cordic/my_rotation/sub_35/carry [12]), .CO(
        \u_cordic/my_rotation/sub_35/carry [13]), .S(
        \u_cordic/my_rotation/delta [12]) );
  ADD32 \u_cordic/my_rotation/sub_35/U2_13  ( .A(
        \u_cordic/my_rotation/present_angle[0][13] ), .B(n172), .CI(
        \u_cordic/my_rotation/sub_35/carry [13]), .CO(
        \u_cordic/my_rotation/sub_35/carry [14]), .S(
        \u_cordic/my_rotation/delta [13]) );
  ADD32 \u_cordic/my_rotation/sub_35/U2_14  ( .A(
        \u_cordic/my_rotation/present_angle[0][14] ), .B(n171), .CI(
        \u_cordic/my_rotation/sub_35/carry [14]), .CO(
        \u_cordic/my_rotation/sub_35/carry [15]), .S(
        \u_cordic/my_rotation/delta [14]) );
  ADD32 \u_cordic/mycordic/r144/U1_4  ( .A(
        \u_cordic/mycordic/present_I_table[1][4] ), .B(
        \u_cordic/mycordic/present_Q_table[1][4] ), .CI(
        \u_cordic/mycordic/r144/carry [4]), .CO(
        \u_cordic/mycordic/r144/carry [5]), .S(\u_cordic/mycordic/N256 ) );
  ADD32 \u_cordic/mycordic/r144/U1_5  ( .A(
        \u_cordic/mycordic/present_I_table[1][5] ), .B(
        \u_cordic/mycordic/present_Q_table[1][5] ), .CI(
        \u_cordic/mycordic/r144/carry [5]), .CO(
        \u_cordic/mycordic/r144/carry [6]), .S(\u_cordic/mycordic/N257 ) );
  ADD32 \u_cordic/mycordic/r144/U1_6  ( .A(
        \u_cordic/mycordic/present_I_table[1][6] ), .B(
        \u_cordic/mycordic/present_Q_table[1][6] ), .CI(
        \u_cordic/mycordic/r144/carry [6]), .CO(
        \u_cordic/mycordic/r144/carry [7]), .S(\u_cordic/mycordic/N258 ) );
  ADD32 \u_cordic/mycordic/r144/U1_7  ( .A(
        \u_cordic/mycordic/present_I_table[1][7] ), .B(
        \u_cordic/mycordic/present_Q_table[1][7] ), .CI(
        \u_cordic/mycordic/r144/carry [7]), .S(\u_cordic/mycordic/N259 ) );
  ADD32 \u_cordic/mycordic/sub_178/U2_4  ( .A(
        \u_cordic/mycordic/present_Q_table[1][4] ), .B(n257), .CI(
        \u_cordic/mycordic/sub_178/carry [4]), .CO(
        \u_cordic/mycordic/sub_178/carry [5]), .S(\u_cordic/mycordic/N264 ) );
  ADD32 \u_cordic/mycordic/sub_178/U2_5  ( .A(
        \u_cordic/mycordic/present_Q_table[1][5] ), .B(n256), .CI(
        \u_cordic/mycordic/sub_178/carry [5]), .CO(
        \u_cordic/mycordic/sub_178/carry [6]), .S(\u_cordic/mycordic/N265 ) );
  ADD32 \u_cordic/mycordic/sub_178/U2_6  ( .A(
        \u_cordic/mycordic/present_Q_table[1][6] ), .B(n291), .CI(
        \u_cordic/mycordic/sub_178/carry [6]), .CO(
        \u_cordic/mycordic/sub_178/carry [7]), .S(\u_cordic/mycordic/N266 ) );
  ADD32 \u_cordic/mycordic/sub_182/U2_4  ( .A(
        \u_cordic/mycordic/present_I_table[1][4] ), .B(n259), .CI(
        \u_cordic/mycordic/sub_182/carry [4]), .CO(
        \u_cordic/mycordic/sub_182/carry [5]), .S(\u_cordic/mycordic/N288 ) );
  ADD32 \u_cordic/mycordic/sub_182/U2_5  ( .A(
        \u_cordic/mycordic/present_I_table[1][5] ), .B(n258), .CI(
        \u_cordic/mycordic/sub_182/carry [5]), .CO(
        \u_cordic/mycordic/sub_182/carry [6]), .S(\u_cordic/mycordic/N289 ) );
  ADD32 \u_cordic/mycordic/sub_182/U2_6  ( .A(
        \u_cordic/mycordic/present_I_table[1][6] ), .B(n292), .CI(
        \u_cordic/mycordic/sub_182/carry [6]), .CO(
        \u_cordic/mycordic/sub_182/carry [7]), .S(\u_cordic/mycordic/N290 ) );
  ADD32 \u_cordic/mycordic/add_189/U1_1  ( .A(
        \u_cordic/mycordic/present_I_table[2][1] ), .B(
        \u_cordic/mycordic/present_Q_table[2][2] ), .CI(
        \u_cordic/mycordic/add_189/carry [1]), .CO(
        \u_cordic/mycordic/add_189/carry [2]), .S(\u_cordic/mycordic/N317 ) );
  ADD32 \u_cordic/mycordic/add_189/U1_2  ( .A(
        \u_cordic/mycordic/present_I_table[2][2] ), .B(
        \u_cordic/mycordic/present_Q_table[2][3] ), .CI(
        \u_cordic/mycordic/add_189/carry [2]), .CO(
        \u_cordic/mycordic/add_189/carry [3]), .S(\u_cordic/mycordic/N318 ) );
  ADD32 \u_cordic/mycordic/add_189/U1_3  ( .A(
        \u_cordic/mycordic/present_I_table[2][3] ), .B(
        \u_cordic/mycordic/present_Q_table[2][4] ), .CI(
        \u_cordic/mycordic/add_189/carry [3]), .CO(
        \u_cordic/mycordic/add_189/carry [4]), .S(\u_cordic/mycordic/N319 ) );
  ADD32 \u_cordic/mycordic/add_189/U1_4  ( .A(
        \u_cordic/mycordic/present_I_table[2][4] ), .B(
        \u_cordic/mycordic/present_Q_table[2][5] ), .CI(
        \u_cordic/mycordic/add_189/carry [4]), .CO(
        \u_cordic/mycordic/add_189/carry [5]), .S(\u_cordic/mycordic/N320 ) );
  ADD32 \u_cordic/mycordic/add_189/U1_5  ( .A(
        \u_cordic/mycordic/present_I_table[2][5] ), .B(
        \u_cordic/mycordic/present_Q_table[2][6] ), .CI(
        \u_cordic/mycordic/add_189/carry [5]), .CO(
        \u_cordic/mycordic/add_189/carry [6]), .S(\u_cordic/mycordic/N321 ) );
  ADD32 \u_cordic/mycordic/add_189/U1_6  ( .A(
        \u_cordic/mycordic/present_I_table[2][6] ), .B(
        \u_cordic/mycordic/present_Q_table[2][7] ), .CI(
        \u_cordic/mycordic/add_189/carry [6]), .CO(
        \u_cordic/mycordic/add_189/carry [7]), .S(\u_cordic/mycordic/N322 ) );
  ADD32 \u_cordic/mycordic/sub_190/U2_1  ( .A(
        \u_cordic/mycordic/present_Q_table[2][1] ), .B(n214), .CI(
        \u_cordic/mycordic/sub_190/carry [1]), .CO(
        \u_cordic/mycordic/sub_190/carry [2]), .S(\u_cordic/mycordic/N325 ) );
  ADD32 \u_cordic/mycordic/sub_190/U2_2  ( .A(
        \u_cordic/mycordic/present_Q_table[2][2] ), .B(n213), .CI(
        \u_cordic/mycordic/sub_190/carry [2]), .CO(
        \u_cordic/mycordic/sub_190/carry [3]), .S(\u_cordic/mycordic/N326 ) );
  ADD32 \u_cordic/mycordic/sub_190/U2_3  ( .A(
        \u_cordic/mycordic/present_Q_table[2][3] ), .B(n212), .CI(
        \u_cordic/mycordic/sub_190/carry [3]), .CO(
        \u_cordic/mycordic/sub_190/carry [4]), .S(\u_cordic/mycordic/N327 ) );
  ADD32 \u_cordic/mycordic/sub_190/U2_4  ( .A(
        \u_cordic/mycordic/present_Q_table[2][4] ), .B(n254), .CI(
        \u_cordic/mycordic/sub_190/carry [4]), .CO(
        \u_cordic/mycordic/sub_190/carry [5]), .S(\u_cordic/mycordic/N328 ) );
  ADD32 \u_cordic/mycordic/sub_190/U2_5  ( .A(
        \u_cordic/mycordic/present_Q_table[2][5] ), .B(n253), .CI(
        \u_cordic/mycordic/sub_190/carry [5]), .CO(
        \u_cordic/mycordic/sub_190/carry [6]), .S(\u_cordic/mycordic/N329 ) );
  ADD32 \u_cordic/mycordic/sub_190/U2_6  ( .A(
        \u_cordic/mycordic/present_Q_table[2][6] ), .B(n288), .CI(
        \u_cordic/mycordic/sub_190/carry [6]), .CO(
        \u_cordic/mycordic/sub_190/carry [7]), .S(\u_cordic/mycordic/N330 ) );
  ADD32 \u_cordic/mycordic/sub_194/U2_1  ( .A(
        \u_cordic/mycordic/present_I_table[2][1] ), .B(n211), .CI(
        \u_cordic/mycordic/sub_194/carry [1]), .CO(
        \u_cordic/mycordic/sub_194/carry [2]), .S(\u_cordic/mycordic/N349 ) );
  ADD32 \u_cordic/mycordic/sub_194/U2_2  ( .A(
        \u_cordic/mycordic/present_I_table[2][2] ), .B(n210), .CI(
        \u_cordic/mycordic/sub_194/carry [2]), .CO(
        \u_cordic/mycordic/sub_194/carry [3]), .S(\u_cordic/mycordic/N350 ) );
  ADD32 \u_cordic/mycordic/sub_194/U2_3  ( .A(
        \u_cordic/mycordic/present_I_table[2][3] ), .B(n209), .CI(
        \u_cordic/mycordic/sub_194/carry [3]), .CO(
        \u_cordic/mycordic/sub_194/carry [4]), .S(\u_cordic/mycordic/N351 ) );
  ADD32 \u_cordic/mycordic/sub_194/U2_4  ( .A(
        \u_cordic/mycordic/present_I_table[2][4] ), .B(n252), .CI(
        \u_cordic/mycordic/sub_194/carry [4]), .CO(
        \u_cordic/mycordic/sub_194/carry [5]), .S(\u_cordic/mycordic/N352 ) );
  ADD32 \u_cordic/mycordic/sub_194/U2_5  ( .A(
        \u_cordic/mycordic/present_I_table[2][5] ), .B(n251), .CI(
        \u_cordic/mycordic/sub_194/carry [5]), .CO(
        \u_cordic/mycordic/sub_194/carry [6]), .S(\u_cordic/mycordic/N353 ) );
  ADD32 \u_cordic/mycordic/sub_194/U2_6  ( .A(
        \u_cordic/mycordic/present_I_table[2][6] ), .B(n287), .CI(
        \u_cordic/mycordic/sub_194/carry [6]), .CO(
        \u_cordic/mycordic/sub_194/carry [7]), .S(\u_cordic/mycordic/N354 ) );
  ADD32 \u_cordic/mycordic/add_195/U1_1  ( .A(
        \u_cordic/mycordic/present_Q_table[2][1] ), .B(
        \u_cordic/mycordic/present_I_table[2][2] ), .CI(
        \u_cordic/mycordic/add_195/carry [1]), .CO(
        \u_cordic/mycordic/add_195/carry [2]), .S(\u_cordic/mycordic/N357 ) );
  ADD32 \u_cordic/mycordic/add_195/U1_2  ( .A(
        \u_cordic/mycordic/present_Q_table[2][2] ), .B(
        \u_cordic/mycordic/present_I_table[2][3] ), .CI(
        \u_cordic/mycordic/add_195/carry [2]), .CO(
        \u_cordic/mycordic/add_195/carry [3]), .S(\u_cordic/mycordic/N358 ) );
  ADD32 \u_cordic/mycordic/add_195/U1_3  ( .A(
        \u_cordic/mycordic/present_Q_table[2][3] ), .B(
        \u_cordic/mycordic/present_I_table[2][4] ), .CI(
        \u_cordic/mycordic/add_195/carry [3]), .CO(
        \u_cordic/mycordic/add_195/carry [4]), .S(\u_cordic/mycordic/N359 ) );
  ADD32 \u_cordic/mycordic/add_195/U1_4  ( .A(
        \u_cordic/mycordic/present_Q_table[2][4] ), .B(
        \u_cordic/mycordic/present_I_table[2][5] ), .CI(
        \u_cordic/mycordic/add_195/carry [4]), .CO(
        \u_cordic/mycordic/add_195/carry [5]), .S(\u_cordic/mycordic/N360 ) );
  ADD32 \u_cordic/mycordic/add_195/U1_5  ( .A(
        \u_cordic/mycordic/present_Q_table[2][5] ), .B(
        \u_cordic/mycordic/present_I_table[2][6] ), .CI(
        \u_cordic/mycordic/add_195/carry [5]), .CO(
        \u_cordic/mycordic/add_195/carry [6]), .S(\u_cordic/mycordic/N361 ) );
  ADD32 \u_cordic/mycordic/add_195/U1_6  ( .A(
        \u_cordic/mycordic/present_Q_table[2][6] ), .B(
        \u_cordic/mycordic/present_I_table[2][7] ), .CI(
        \u_cordic/mycordic/add_195/carry [6]), .CO(
        \u_cordic/mycordic/add_195/carry [7]), .S(\u_cordic/mycordic/N362 ) );
  ADD32 \u_cordic/mycordic/add_200/U1_1  ( .A(
        \u_cordic/mycordic/present_I_table[3][1] ), .B(
        \u_cordic/mycordic/present_Q_table[3][3] ), .CI(
        \u_cordic/mycordic/add_200/carry [1]), .CO(
        \u_cordic/mycordic/add_200/carry [2]), .S(\u_cordic/mycordic/N381 ) );
  ADD32 \u_cordic/mycordic/add_200/U1_2  ( .A(
        \u_cordic/mycordic/present_I_table[3][2] ), .B(
        \u_cordic/mycordic/present_Q_table[3][4] ), .CI(
        \u_cordic/mycordic/add_200/carry [2]), .CO(
        \u_cordic/mycordic/add_200/carry [3]), .S(\u_cordic/mycordic/N382 ) );
  ADD32 \u_cordic/mycordic/add_200/U1_3  ( .A(
        \u_cordic/mycordic/present_I_table[3][3] ), .B(
        \u_cordic/mycordic/present_Q_table[3][5] ), .CI(
        \u_cordic/mycordic/add_200/carry [3]), .CO(
        \u_cordic/mycordic/add_200/carry [4]), .S(\u_cordic/mycordic/N383 ) );
  ADD32 \u_cordic/mycordic/add_200/U1_4  ( .A(
        \u_cordic/mycordic/present_I_table[3][4] ), .B(
        \u_cordic/mycordic/present_Q_table[3][6] ), .CI(
        \u_cordic/mycordic/add_200/carry [4]), .CO(
        \u_cordic/mycordic/add_200/carry [5]), .S(\u_cordic/mycordic/N384 ) );
  ADD32 \u_cordic/mycordic/add_200/U1_5  ( .A(
        \u_cordic/mycordic/present_I_table[3][5] ), .B(
        \u_cordic/mycordic/present_Q_table[3][7] ), .CI(
        \u_cordic/mycordic/add_200/carry [5]), .CO(
        \u_cordic/mycordic/add_200/carry [6]), .S(\u_cordic/mycordic/N385 ) );
  ADD32 \u_cordic/mycordic/add_200/U1_6  ( .A(
        \u_cordic/mycordic/present_I_table[3][6] ), .B(
        \u_cordic/mycordic/present_Q_table[3][7] ), .CI(
        \u_cordic/mycordic/add_200/carry [6]), .CO(
        \u_cordic/mycordic/add_200/carry [7]), .S(\u_cordic/mycordic/N386 ) );
  ADD32 \u_cordic/mycordic/sub_201/U2_1  ( .A(
        \u_cordic/mycordic/present_Q_table[3][1] ), .B(n208), .CI(
        \u_cordic/mycordic/sub_201/carry [1]), .CO(
        \u_cordic/mycordic/sub_201/carry [2]), .S(\u_cordic/mycordic/N389 ) );
  ADD32 \u_cordic/mycordic/sub_201/U2_2  ( .A(
        \u_cordic/mycordic/present_Q_table[3][2] ), .B(n207), .CI(
        \u_cordic/mycordic/sub_201/carry [2]), .CO(
        \u_cordic/mycordic/sub_201/carry [3]), .S(\u_cordic/mycordic/N390 ) );
  ADD32 \u_cordic/mycordic/sub_201/U2_3  ( .A(
        \u_cordic/mycordic/present_Q_table[3][3] ), .B(n206), .CI(
        \u_cordic/mycordic/sub_201/carry [3]), .CO(
        \u_cordic/mycordic/sub_201/carry [4]), .S(\u_cordic/mycordic/N391 ) );
  ADD32 \u_cordic/mycordic/sub_201/U2_4  ( .A(
        \u_cordic/mycordic/present_Q_table[3][4] ), .B(n250), .CI(
        \u_cordic/mycordic/sub_201/carry [4]), .CO(
        \u_cordic/mycordic/sub_201/carry [5]), .S(\u_cordic/mycordic/N392 ) );
  ADD32 \u_cordic/mycordic/sub_201/U2_5  ( .A(
        \u_cordic/mycordic/present_Q_table[3][5] ), .B(n246), .CI(
        \u_cordic/mycordic/sub_201/carry [5]), .CO(
        \u_cordic/mycordic/sub_201/carry [6]), .S(\u_cordic/mycordic/N393 ) );
  ADD32 \u_cordic/mycordic/sub_201/U2_6  ( .A(
        \u_cordic/mycordic/present_Q_table[3][6] ), .B(n246), .CI(
        \u_cordic/mycordic/sub_201/carry [6]), .CO(
        \u_cordic/mycordic/sub_201/carry [7]), .S(\u_cordic/mycordic/N394 ) );
  ADD32 \u_cordic/mycordic/sub_205/U2_1  ( .A(
        \u_cordic/mycordic/present_I_table[3][1] ), .B(n205), .CI(
        \u_cordic/mycordic/sub_205/carry [1]), .CO(
        \u_cordic/mycordic/sub_205/carry [2]), .S(\u_cordic/mycordic/N413 ) );
  ADD32 \u_cordic/mycordic/sub_205/U2_2  ( .A(
        \u_cordic/mycordic/present_I_table[3][2] ), .B(n204), .CI(
        \u_cordic/mycordic/sub_205/carry [2]), .CO(
        \u_cordic/mycordic/sub_205/carry [3]), .S(\u_cordic/mycordic/N414 ) );
  ADD32 \u_cordic/mycordic/sub_205/U2_3  ( .A(
        \u_cordic/mycordic/present_I_table[3][3] ), .B(n203), .CI(
        \u_cordic/mycordic/sub_205/carry [3]), .CO(
        \u_cordic/mycordic/sub_205/carry [4]), .S(\u_cordic/mycordic/N415 ) );
  ADD32 \u_cordic/mycordic/sub_205/U2_4  ( .A(
        \u_cordic/mycordic/present_I_table[3][4] ), .B(n249), .CI(
        \u_cordic/mycordic/sub_205/carry [4]), .CO(
        \u_cordic/mycordic/sub_205/carry [5]), .S(\u_cordic/mycordic/N416 ) );
  ADD32 \u_cordic/mycordic/sub_205/U2_5  ( .A(
        \u_cordic/mycordic/present_I_table[3][5] ), .B(n245), .CI(
        \u_cordic/mycordic/sub_205/carry [5]), .CO(
        \u_cordic/mycordic/sub_205/carry [6]), .S(\u_cordic/mycordic/N417 ) );
  ADD32 \u_cordic/mycordic/sub_205/U2_6  ( .A(
        \u_cordic/mycordic/present_I_table[3][6] ), .B(n245), .CI(
        \u_cordic/mycordic/sub_205/carry [6]), .CO(
        \u_cordic/mycordic/sub_205/carry [7]), .S(\u_cordic/mycordic/N418 ) );
  ADD32 \u_cordic/mycordic/add_206/U1_1  ( .A(
        \u_cordic/mycordic/present_Q_table[3][1] ), .B(
        \u_cordic/mycordic/present_I_table[3][3] ), .CI(
        \u_cordic/mycordic/add_206/carry [1]), .CO(
        \u_cordic/mycordic/add_206/carry [2]), .S(\u_cordic/mycordic/N421 ) );
  ADD32 \u_cordic/mycordic/add_206/U1_2  ( .A(
        \u_cordic/mycordic/present_Q_table[3][2] ), .B(
        \u_cordic/mycordic/present_I_table[3][4] ), .CI(
        \u_cordic/mycordic/add_206/carry [2]), .CO(
        \u_cordic/mycordic/add_206/carry [3]), .S(\u_cordic/mycordic/N422 ) );
  ADD32 \u_cordic/mycordic/add_206/U1_3  ( .A(
        \u_cordic/mycordic/present_Q_table[3][3] ), .B(
        \u_cordic/mycordic/present_I_table[3][5] ), .CI(
        \u_cordic/mycordic/add_206/carry [3]), .CO(
        \u_cordic/mycordic/add_206/carry [4]), .S(\u_cordic/mycordic/N423 ) );
  ADD32 \u_cordic/mycordic/add_206/U1_4  ( .A(
        \u_cordic/mycordic/present_Q_table[3][4] ), .B(
        \u_cordic/mycordic/present_I_table[3][6] ), .CI(
        \u_cordic/mycordic/add_206/carry [4]), .CO(
        \u_cordic/mycordic/add_206/carry [5]), .S(\u_cordic/mycordic/N424 ) );
  ADD32 \u_cordic/mycordic/add_206/U1_5  ( .A(
        \u_cordic/mycordic/present_Q_table[3][5] ), .B(
        \u_cordic/mycordic/present_I_table[3][7] ), .CI(
        \u_cordic/mycordic/add_206/carry [5]), .CO(
        \u_cordic/mycordic/add_206/carry [6]), .S(\u_cordic/mycordic/N425 ) );
  ADD32 \u_cordic/mycordic/add_206/U1_6  ( .A(
        \u_cordic/mycordic/present_Q_table[3][6] ), .B(
        \u_cordic/mycordic/present_I_table[3][7] ), .CI(
        \u_cordic/mycordic/add_206/carry [6]), .CO(
        \u_cordic/mycordic/add_206/carry [7]), .S(\u_cordic/mycordic/N426 ) );
  ADD32 \u_cordic/mycordic/add_211/U1_4  ( .A(
        \u_cordic/mycordic/present_I_table[4][4] ), .B(
        \u_cordic/mycordic/present_Q_table[4][7] ), .CI(n2654), .CO(
        \u_cordic/mycordic/add_211/carry [5]), .S(\u_cordic/mycordic/N444 ) );
  ADD32 \u_cordic/mycordic/add_211/U1_5  ( .A(
        \u_cordic/mycordic/present_I_table[4][5] ), .B(
        \u_cordic/mycordic/present_Q_table[4][7] ), .CI(
        \u_cordic/mycordic/add_211/carry [5]), .CO(
        \u_cordic/mycordic/add_211/carry [6]), .S(\u_cordic/mycordic/N445 ) );
  ADD32 \u_cordic/mycordic/add_211/U1_6  ( .A(
        \u_cordic/mycordic/present_I_table[4][6] ), .B(
        \u_cordic/mycordic/present_Q_table[4][7] ), .CI(
        \u_cordic/mycordic/add_211/carry [6]), .CO(
        \u_cordic/mycordic/add_211/carry [7]), .S(\u_cordic/mycordic/N446 ) );
  ADD32 \u_cordic/mycordic/sub_212/U2_1  ( .A(
        \u_cordic/mycordic/present_Q_table[4][1] ), .B(n202), .CI(
        \u_cordic/mycordic/sub_212/carry [1]), .CO(
        \u_cordic/mycordic/sub_212/carry [2]), .S(\u_cordic/mycordic/N449 ) );
  ADD32 \u_cordic/mycordic/sub_212/U2_2  ( .A(
        \u_cordic/mycordic/present_Q_table[4][2] ), .B(n201), .CI(
        \u_cordic/mycordic/sub_212/carry [2]), .CO(
        \u_cordic/mycordic/sub_212/carry [3]), .S(\u_cordic/mycordic/N450 ) );
  ADD32 \u_cordic/mycordic/sub_212/U2_3  ( .A(
        \u_cordic/mycordic/present_Q_table[4][3] ), .B(n200), .CI(
        \u_cordic/mycordic/sub_212/carry [3]), .CO(
        \u_cordic/mycordic/sub_212/carry [4]), .S(\u_cordic/mycordic/N451 ) );
  ADD32 \u_cordic/mycordic/sub_212/U2_4  ( .A(
        \u_cordic/mycordic/present_Q_table[4][4] ), .B(n47), .CI(
        \u_cordic/mycordic/sub_212/carry [4]), .CO(
        \u_cordic/mycordic/sub_212/carry [5]), .S(\u_cordic/mycordic/N452 ) );
  ADD32 \u_cordic/mycordic/sub_212/U2_5  ( .A(
        \u_cordic/mycordic/present_Q_table[4][5] ), .B(n47), .CI(
        \u_cordic/mycordic/sub_212/carry [5]), .CO(
        \u_cordic/mycordic/sub_212/carry [6]), .S(\u_cordic/mycordic/N453 ) );
  ADD32 \u_cordic/mycordic/sub_212/U2_6  ( .A(
        \u_cordic/mycordic/present_Q_table[4][6] ), .B(n47), .CI(
        \u_cordic/mycordic/sub_212/carry [6]), .CO(
        \u_cordic/mycordic/sub_212/carry [7]), .S(\u_cordic/mycordic/N454 ) );
  ADD32 \u_cordic/mycordic/sub_216/U2_4  ( .A(
        \u_cordic/mycordic/present_I_table[4][4] ), .B(n48), .CI(
        \u_cordic/mycordic/sub_216/carry [4]), .CO(
        \u_cordic/mycordic/sub_216/carry [5]), .S(\u_cordic/mycordic/N472 ) );
  ADD32 \u_cordic/mycordic/sub_216/U2_5  ( .A(
        \u_cordic/mycordic/present_I_table[4][5] ), .B(n48), .CI(
        \u_cordic/mycordic/sub_216/carry [5]), .CO(
        \u_cordic/mycordic/sub_216/carry [6]), .S(\u_cordic/mycordic/N473 ) );
  ADD32 \u_cordic/mycordic/sub_216/U2_6  ( .A(
        \u_cordic/mycordic/present_I_table[4][6] ), .B(n48), .CI(
        \u_cordic/mycordic/sub_216/carry [6]), .CO(
        \u_cordic/mycordic/sub_216/carry [7]), .S(\u_cordic/mycordic/N474 ) );
  ADD32 \u_cordic/mycordic/add_217/U1_1  ( .A(
        \u_cordic/mycordic/present_Q_table[4][1] ), .B(
        \u_cordic/mycordic/present_I_table[4][4] ), .CI(
        \u_cordic/mycordic/add_217/carry [1]), .CO(
        \u_cordic/mycordic/add_217/carry [2]), .S(\u_cordic/mycordic/N477 ) );
  ADD32 \u_cordic/mycordic/add_217/U1_2  ( .A(
        \u_cordic/mycordic/present_Q_table[4][2] ), .B(
        \u_cordic/mycordic/present_I_table[4][5] ), .CI(
        \u_cordic/mycordic/add_217/carry [2]), .CO(
        \u_cordic/mycordic/add_217/carry [3]), .S(\u_cordic/mycordic/N478 ) );
  ADD32 \u_cordic/mycordic/add_217/U1_3  ( .A(
        \u_cordic/mycordic/present_Q_table[4][3] ), .B(
        \u_cordic/mycordic/present_I_table[4][6] ), .CI(
        \u_cordic/mycordic/add_217/carry [3]), .CO(
        \u_cordic/mycordic/add_217/carry [4]), .S(\u_cordic/mycordic/N479 ) );
  ADD32 \u_cordic/mycordic/add_217/U1_4  ( .A(
        \u_cordic/mycordic/present_Q_table[4][4] ), .B(
        \u_cordic/mycordic/present_I_table[4][7] ), .CI(
        \u_cordic/mycordic/add_217/carry [4]), .CO(
        \u_cordic/mycordic/add_217/carry [5]), .S(\u_cordic/mycordic/N480 ) );
  ADD32 \u_cordic/mycordic/add_217/U1_5  ( .A(
        \u_cordic/mycordic/present_Q_table[4][5] ), .B(
        \u_cordic/mycordic/present_I_table[4][7] ), .CI(
        \u_cordic/mycordic/add_217/carry [5]), .CO(
        \u_cordic/mycordic/add_217/carry [6]), .S(\u_cordic/mycordic/N481 ) );
  ADD32 \u_cordic/mycordic/add_217/U1_6  ( .A(
        \u_cordic/mycordic/present_Q_table[4][6] ), .B(
        \u_cordic/mycordic/present_I_table[4][7] ), .CI(
        \u_cordic/mycordic/add_217/carry [6]), .CO(
        \u_cordic/mycordic/add_217/carry [7]), .S(\u_cordic/mycordic/N482 ) );
  ADD32 \u_decoder/fir_filter/add_294/U1_11  ( .A(
        \u_decoder/fir_filter/I_data_mult_0_buff [11]), .B(
        \u_decoder/fir_filter/I_data_add_1_buff [11]), .CI(
        \u_decoder/fir_filter/add_294/carry [11]), .CO(
        \u_decoder/fir_filter/add_294/carry [12]), .S(
        \u_decoder/fir_filter/I_data_add_0 [11]) );
  ADD32 \u_decoder/fir_filter/add_294/U1_12  ( .A(
        \u_decoder/fir_filter/I_data_mult_0_buff [12]), .B(
        \u_decoder/fir_filter/I_data_add_1_buff [12]), .CI(
        \u_decoder/fir_filter/add_294/carry [12]), .CO(
        \u_decoder/fir_filter/add_294/carry [13]), .S(
        \u_decoder/fir_filter/I_data_add_0 [12]) );
  ADD32 \u_decoder/fir_filter/add_294/U1_13  ( .A(
        \u_decoder/fir_filter/I_data_mult_0_buff [13]), .B(
        \u_decoder/fir_filter/I_data_add_1_buff [13]), .CI(
        \u_decoder/fir_filter/add_294/carry [13]), .CO(
        \u_decoder/fir_filter/add_294/carry [14]), .S(
        \u_decoder/fir_filter/I_data_add_0 [13]) );
  ADD32 \u_decoder/fir_filter/add_295/U1_1  ( .A(
        \u_decoder/fir_filter/I_data_mult_1_buff [1]), .B(
        \u_decoder/fir_filter/I_data_add_2_buff [1]), .CI(
        \u_decoder/fir_filter/add_295/carry [1]), .CO(
        \u_decoder/fir_filter/add_295/carry [2]), .S(
        \u_decoder/fir_filter/I_data_add_1 [1]) );
  ADD32 \u_decoder/fir_filter/add_295/U1_2  ( .A(
        \u_decoder/fir_filter/I_data_mult_1_buff [2]), .B(
        \u_decoder/fir_filter/I_data_add_2_buff [2]), .CI(
        \u_decoder/fir_filter/add_295/carry [2]), .CO(
        \u_decoder/fir_filter/add_295/carry [3]), .S(
        \u_decoder/fir_filter/I_data_add_1 [2]) );
  ADD32 \u_decoder/fir_filter/add_295/U1_3  ( .A(
        \u_decoder/fir_filter/I_data_mult_1_buff [3]), .B(
        \u_decoder/fir_filter/I_data_add_2_buff [3]), .CI(
        \u_decoder/fir_filter/add_295/carry [3]), .CO(
        \u_decoder/fir_filter/add_295/carry [4]), .S(
        \u_decoder/fir_filter/I_data_add_1 [3]) );
  ADD32 \u_decoder/fir_filter/add_295/U1_4  ( .A(
        \u_decoder/fir_filter/I_data_mult_1_buff [4]), .B(
        \u_decoder/fir_filter/I_data_add_2_buff [4]), .CI(
        \u_decoder/fir_filter/add_295/carry [4]), .CO(
        \u_decoder/fir_filter/add_295/carry [5]), .S(
        \u_decoder/fir_filter/I_data_add_1 [4]) );
  ADD32 \u_decoder/fir_filter/add_295/U1_5  ( .A(
        \u_decoder/fir_filter/I_data_mult_1_buff [5]), .B(
        \u_decoder/fir_filter/I_data_add_2_buff [5]), .CI(
        \u_decoder/fir_filter/add_295/carry [5]), .CO(
        \u_decoder/fir_filter/add_295/carry [6]), .S(
        \u_decoder/fir_filter/I_data_add_1 [5]) );
  ADD32 \u_decoder/fir_filter/add_295/U1_6  ( .A(
        \u_decoder/fir_filter/I_data_mult_1_buff [6]), .B(
        \u_decoder/fir_filter/I_data_add_2_buff [6]), .CI(
        \u_decoder/fir_filter/add_295/carry [6]), .CO(
        \u_decoder/fir_filter/add_295/carry [7]), .S(
        \u_decoder/fir_filter/I_data_add_1 [6]) );
  ADD32 \u_decoder/fir_filter/add_295/U1_7  ( .A(
        \u_decoder/fir_filter/I_data_mult_1_buff [7]), .B(
        \u_decoder/fir_filter/I_data_add_2_buff [7]), .CI(
        \u_decoder/fir_filter/add_295/carry [7]), .CO(
        \u_decoder/fir_filter/add_295/carry [8]), .S(
        \u_decoder/fir_filter/I_data_add_1 [7]) );
  ADD32 \u_decoder/fir_filter/add_295/U1_8  ( .A(
        \u_decoder/fir_filter/I_data_mult_1_buff [8]), .B(
        \u_decoder/fir_filter/I_data_add_2_buff [8]), .CI(
        \u_decoder/fir_filter/add_295/carry [8]), .CO(
        \u_decoder/fir_filter/add_295/carry [9]), .S(
        \u_decoder/fir_filter/I_data_add_1 [8]) );
  ADD32 \u_decoder/fir_filter/add_295/U1_9  ( .A(
        \u_decoder/fir_filter/I_data_mult_1_buff [9]), .B(
        \u_decoder/fir_filter/I_data_add_2_buff [9]), .CI(
        \u_decoder/fir_filter/add_295/carry [9]), .CO(
        \u_decoder/fir_filter/add_295/carry [10]), .S(
        \u_decoder/fir_filter/I_data_add_1 [9]) );
  ADD32 \u_decoder/fir_filter/add_295/U1_10  ( .A(
        \u_decoder/fir_filter/I_data_mult_1_buff [10]), .B(
        \u_decoder/fir_filter/I_data_add_2_buff [10]), .CI(
        \u_decoder/fir_filter/add_295/carry [10]), .CO(
        \u_decoder/fir_filter/add_295/carry [11]), .S(
        \u_decoder/fir_filter/I_data_add_1 [10]) );
  ADD32 \u_decoder/fir_filter/add_295/U1_11  ( .A(
        \u_decoder/fir_filter/I_data_mult_1_buff [11]), .B(
        \u_decoder/fir_filter/I_data_add_2_buff [11]), .CI(
        \u_decoder/fir_filter/add_295/carry [11]), .CO(
        \u_decoder/fir_filter/add_295/carry [12]), .S(
        \u_decoder/fir_filter/I_data_add_1 [11]) );
  ADD32 \u_decoder/fir_filter/add_295/U1_12  ( .A(
        \u_decoder/fir_filter/I_data_mult_1_buff [12]), .B(
        \u_decoder/fir_filter/I_data_add_2_buff [12]), .CI(
        \u_decoder/fir_filter/add_295/carry [12]), .CO(
        \u_decoder/fir_filter/add_295/carry [13]), .S(
        \u_decoder/fir_filter/I_data_add_1 [12]) );
  ADD32 \u_decoder/fir_filter/add_295/U1_13  ( .A(
        \u_decoder/fir_filter/I_data_mult_1_buff [13]), .B(
        \u_decoder/fir_filter/I_data_add_2_buff [13]), .CI(
        \u_decoder/fir_filter/add_295/carry [13]), .CO(
        \u_decoder/fir_filter/add_295/carry [14]), .S(
        \u_decoder/fir_filter/I_data_add_1 [13]) );
  ADD32 \u_decoder/fir_filter/add_296/U1_1  ( .A(
        \u_decoder/fir_filter/I_data_mult_2_buff [1]), .B(
        \u_decoder/fir_filter/I_data_add_3_buff [1]), .CI(
        \u_decoder/fir_filter/add_296/carry [1]), .CO(
        \u_decoder/fir_filter/add_296/carry [2]), .S(
        \u_decoder/fir_filter/I_data_add_2 [1]) );
  ADD32 \u_decoder/fir_filter/add_296/U1_2  ( .A(
        \u_decoder/fir_filter/I_data_mult_2_buff [2]), .B(
        \u_decoder/fir_filter/I_data_add_3_buff [2]), .CI(
        \u_decoder/fir_filter/add_296/carry [2]), .CO(
        \u_decoder/fir_filter/add_296/carry [3]), .S(
        \u_decoder/fir_filter/I_data_add_2 [2]) );
  ADD32 \u_decoder/fir_filter/add_296/U1_3  ( .A(
        \u_decoder/fir_filter/I_data_mult_2_buff [3]), .B(
        \u_decoder/fir_filter/I_data_add_3_buff [3]), .CI(
        \u_decoder/fir_filter/add_296/carry [3]), .CO(
        \u_decoder/fir_filter/add_296/carry [4]), .S(
        \u_decoder/fir_filter/I_data_add_2 [3]) );
  ADD32 \u_decoder/fir_filter/add_296/U1_4  ( .A(
        \u_decoder/fir_filter/I_data_mult_2_buff [4]), .B(
        \u_decoder/fir_filter/I_data_add_3_buff [4]), .CI(
        \u_decoder/fir_filter/add_296/carry [4]), .CO(
        \u_decoder/fir_filter/add_296/carry [5]), .S(
        \u_decoder/fir_filter/I_data_add_2 [4]) );
  ADD32 \u_decoder/fir_filter/add_296/U1_5  ( .A(
        \u_decoder/fir_filter/I_data_mult_2_buff [5]), .B(
        \u_decoder/fir_filter/I_data_add_3_buff [5]), .CI(
        \u_decoder/fir_filter/add_296/carry [5]), .CO(
        \u_decoder/fir_filter/add_296/carry [6]), .S(
        \u_decoder/fir_filter/I_data_add_2 [5]) );
  ADD32 \u_decoder/fir_filter/add_296/U1_6  ( .A(
        \u_decoder/fir_filter/I_data_mult_2_buff [6]), .B(
        \u_decoder/fir_filter/I_data_add_3_buff [6]), .CI(
        \u_decoder/fir_filter/add_296/carry [6]), .CO(
        \u_decoder/fir_filter/add_296/carry [7]), .S(
        \u_decoder/fir_filter/I_data_add_2 [6]) );
  ADD32 \u_decoder/fir_filter/add_296/U1_7  ( .A(
        \u_decoder/fir_filter/I_data_mult_2_buff [7]), .B(
        \u_decoder/fir_filter/I_data_add_3_buff [7]), .CI(
        \u_decoder/fir_filter/add_296/carry [7]), .CO(
        \u_decoder/fir_filter/add_296/carry [8]), .S(
        \u_decoder/fir_filter/I_data_add_2 [7]) );
  ADD32 \u_decoder/fir_filter/add_296/U1_8  ( .A(
        \u_decoder/fir_filter/I_data_mult_2_buff [8]), .B(
        \u_decoder/fir_filter/I_data_add_3_buff [8]), .CI(
        \u_decoder/fir_filter/add_296/carry [8]), .CO(
        \u_decoder/fir_filter/add_296/carry [9]), .S(
        \u_decoder/fir_filter/I_data_add_2 [8]) );
  ADD32 \u_decoder/fir_filter/add_296/U1_9  ( .A(
        \u_decoder/fir_filter/I_data_mult_2_buff [9]), .B(
        \u_decoder/fir_filter/I_data_add_3_buff [9]), .CI(
        \u_decoder/fir_filter/add_296/carry [9]), .CO(
        \u_decoder/fir_filter/add_296/carry [10]), .S(
        \u_decoder/fir_filter/I_data_add_2 [9]) );
  ADD32 \u_decoder/fir_filter/add_296/U1_10  ( .A(
        \u_decoder/fir_filter/I_data_mult_2_buff [10]), .B(
        \u_decoder/fir_filter/I_data_add_3_buff [10]), .CI(
        \u_decoder/fir_filter/add_296/carry [10]), .CO(
        \u_decoder/fir_filter/add_296/carry [11]), .S(
        \u_decoder/fir_filter/I_data_add_2 [10]) );
  ADD32 \u_decoder/fir_filter/add_296/U1_11  ( .A(
        \u_decoder/fir_filter/I_data_mult_2_buff [11]), .B(
        \u_decoder/fir_filter/I_data_add_3_buff [11]), .CI(
        \u_decoder/fir_filter/add_296/carry [11]), .CO(
        \u_decoder/fir_filter/add_296/carry [12]), .S(
        \u_decoder/fir_filter/I_data_add_2 [11]) );
  ADD32 \u_decoder/fir_filter/add_296/U1_12  ( .A(
        \u_decoder/fir_filter/I_data_mult_2_buff [12]), .B(
        \u_decoder/fir_filter/I_data_add_3_buff [12]), .CI(
        \u_decoder/fir_filter/add_296/carry [12]), .CO(
        \u_decoder/fir_filter/add_296/carry [13]), .S(
        \u_decoder/fir_filter/I_data_add_2 [12]) );
  ADD32 \u_decoder/fir_filter/add_296/U1_13  ( .A(
        \u_decoder/fir_filter/I_data_mult_2_buff [13]), .B(
        \u_decoder/fir_filter/I_data_add_3_buff [13]), .CI(
        \u_decoder/fir_filter/add_296/carry [13]), .CO(
        \u_decoder/fir_filter/add_296/carry [14]), .S(
        \u_decoder/fir_filter/I_data_add_2 [13]) );
  ADD32 \u_decoder/fir_filter/add_297/U1_1  ( .A(
        \u_decoder/fir_filter/I_data_mult_3_buff [1]), .B(
        \u_decoder/fir_filter/I_data_add_4_buff [1]), .CI(
        \u_decoder/fir_filter/add_297/carry [1]), .CO(
        \u_decoder/fir_filter/add_297/carry [2]), .S(
        \u_decoder/fir_filter/I_data_add_3 [1]) );
  ADD32 \u_decoder/fir_filter/add_297/U1_2  ( .A(
        \u_decoder/fir_filter/I_data_mult_3_buff [2]), .B(
        \u_decoder/fir_filter/I_data_add_4_buff [2]), .CI(
        \u_decoder/fir_filter/add_297/carry [2]), .CO(
        \u_decoder/fir_filter/add_297/carry [3]), .S(
        \u_decoder/fir_filter/I_data_add_3 [2]) );
  ADD32 \u_decoder/fir_filter/add_297/U1_3  ( .A(
        \u_decoder/fir_filter/I_data_mult_3_buff [3]), .B(
        \u_decoder/fir_filter/I_data_add_4_buff [3]), .CI(
        \u_decoder/fir_filter/add_297/carry [3]), .CO(
        \u_decoder/fir_filter/add_297/carry [4]), .S(
        \u_decoder/fir_filter/I_data_add_3 [3]) );
  ADD32 \u_decoder/fir_filter/add_297/U1_4  ( .A(
        \u_decoder/fir_filter/I_data_mult_3_buff [4]), .B(
        \u_decoder/fir_filter/I_data_add_4_buff [4]), .CI(
        \u_decoder/fir_filter/add_297/carry [4]), .CO(
        \u_decoder/fir_filter/add_297/carry [5]), .S(
        \u_decoder/fir_filter/I_data_add_3 [4]) );
  ADD32 \u_decoder/fir_filter/add_297/U1_5  ( .A(
        \u_decoder/fir_filter/I_data_mult_3_buff [5]), .B(
        \u_decoder/fir_filter/I_data_add_4_buff [5]), .CI(
        \u_decoder/fir_filter/add_297/carry [5]), .CO(
        \u_decoder/fir_filter/add_297/carry [6]), .S(
        \u_decoder/fir_filter/I_data_add_3 [5]) );
  ADD32 \u_decoder/fir_filter/add_297/U1_6  ( .A(
        \u_decoder/fir_filter/I_data_mult_3_buff [6]), .B(
        \u_decoder/fir_filter/I_data_add_4_buff [6]), .CI(
        \u_decoder/fir_filter/add_297/carry [6]), .CO(
        \u_decoder/fir_filter/add_297/carry [7]), .S(
        \u_decoder/fir_filter/I_data_add_3 [6]) );
  ADD32 \u_decoder/fir_filter/add_297/U1_7  ( .A(
        \u_decoder/fir_filter/I_data_mult_3_buff [7]), .B(
        \u_decoder/fir_filter/I_data_add_4_buff [7]), .CI(
        \u_decoder/fir_filter/add_297/carry [7]), .CO(
        \u_decoder/fir_filter/add_297/carry [8]), .S(
        \u_decoder/fir_filter/I_data_add_3 [7]) );
  ADD32 \u_decoder/fir_filter/add_297/U1_8  ( .A(
        \u_decoder/fir_filter/I_data_mult_3_buff [8]), .B(
        \u_decoder/fir_filter/I_data_add_4_buff [8]), .CI(
        \u_decoder/fir_filter/add_297/carry [8]), .CO(
        \u_decoder/fir_filter/add_297/carry [9]), .S(
        \u_decoder/fir_filter/I_data_add_3 [8]) );
  ADD32 \u_decoder/fir_filter/add_297/U1_9  ( .A(
        \u_decoder/fir_filter/I_data_mult_3_buff [9]), .B(
        \u_decoder/fir_filter/I_data_add_4_buff [9]), .CI(
        \u_decoder/fir_filter/add_297/carry [9]), .CO(
        \u_decoder/fir_filter/add_297/carry [10]), .S(
        \u_decoder/fir_filter/I_data_add_3 [9]) );
  ADD32 \u_decoder/fir_filter/add_297/U1_10  ( .A(
        \u_decoder/fir_filter/I_data_mult_3_buff [10]), .B(
        \u_decoder/fir_filter/I_data_add_4_buff [10]), .CI(
        \u_decoder/fir_filter/add_297/carry [10]), .CO(
        \u_decoder/fir_filter/add_297/carry [11]), .S(
        \u_decoder/fir_filter/I_data_add_3 [10]) );
  ADD32 \u_decoder/fir_filter/add_297/U1_11  ( .A(
        \u_decoder/fir_filter/I_data_mult_3_buff [11]), .B(
        \u_decoder/fir_filter/I_data_add_4_buff [11]), .CI(
        \u_decoder/fir_filter/add_297/carry [11]), .CO(
        \u_decoder/fir_filter/add_297/carry [12]), .S(
        \u_decoder/fir_filter/I_data_add_3 [11]) );
  ADD32 \u_decoder/fir_filter/add_297/U1_12  ( .A(
        \u_decoder/fir_filter/I_data_mult_3_buff [12]), .B(
        \u_decoder/fir_filter/I_data_add_4_buff [12]), .CI(
        \u_decoder/fir_filter/add_297/carry [12]), .CO(
        \u_decoder/fir_filter/add_297/carry [13]), .S(
        \u_decoder/fir_filter/I_data_add_3 [12]) );
  ADD32 \u_decoder/fir_filter/add_297/U1_13  ( .A(
        \u_decoder/fir_filter/I_data_mult_3_buff [13]), .B(
        \u_decoder/fir_filter/I_data_add_4_buff [13]), .CI(
        \u_decoder/fir_filter/add_297/carry [13]), .CO(
        \u_decoder/fir_filter/add_297/carry [14]), .S(
        \u_decoder/fir_filter/I_data_add_3 [13]) );
  ADD32 \u_decoder/fir_filter/add_298/U1_1  ( .A(
        \u_decoder/fir_filter/I_data_mult_4_buff [1]), .B(
        \u_decoder/fir_filter/I_data_add_5_buff [1]), .CI(
        \u_decoder/fir_filter/add_298/carry [1]), .CO(
        \u_decoder/fir_filter/add_298/carry [2]), .S(
        \u_decoder/fir_filter/I_data_add_4 [1]) );
  ADD32 \u_decoder/fir_filter/add_298/U1_2  ( .A(
        \u_decoder/fir_filter/I_data_mult_4_buff [2]), .B(
        \u_decoder/fir_filter/I_data_add_5_buff [2]), .CI(
        \u_decoder/fir_filter/add_298/carry [2]), .CO(
        \u_decoder/fir_filter/add_298/carry [3]), .S(
        \u_decoder/fir_filter/I_data_add_4 [2]) );
  ADD32 \u_decoder/fir_filter/add_298/U1_3  ( .A(
        \u_decoder/fir_filter/I_data_mult_4_buff [3]), .B(
        \u_decoder/fir_filter/I_data_add_5_buff [3]), .CI(
        \u_decoder/fir_filter/add_298/carry [3]), .CO(
        \u_decoder/fir_filter/add_298/carry [4]), .S(
        \u_decoder/fir_filter/I_data_add_4 [3]) );
  ADD32 \u_decoder/fir_filter/add_298/U1_4  ( .A(
        \u_decoder/fir_filter/I_data_mult_4_buff [4]), .B(
        \u_decoder/fir_filter/I_data_add_5_buff [4]), .CI(
        \u_decoder/fir_filter/add_298/carry [4]), .CO(
        \u_decoder/fir_filter/add_298/carry [5]), .S(
        \u_decoder/fir_filter/I_data_add_4 [4]) );
  ADD32 \u_decoder/fir_filter/add_298/U1_5  ( .A(
        \u_decoder/fir_filter/I_data_mult_4_buff [5]), .B(
        \u_decoder/fir_filter/I_data_add_5_buff [5]), .CI(
        \u_decoder/fir_filter/add_298/carry [5]), .CO(
        \u_decoder/fir_filter/add_298/carry [6]), .S(
        \u_decoder/fir_filter/I_data_add_4 [5]) );
  ADD32 \u_decoder/fir_filter/add_298/U1_6  ( .A(
        \u_decoder/fir_filter/I_data_mult_4_buff [6]), .B(
        \u_decoder/fir_filter/I_data_add_5_buff [6]), .CI(
        \u_decoder/fir_filter/add_298/carry [6]), .CO(
        \u_decoder/fir_filter/add_298/carry [7]), .S(
        \u_decoder/fir_filter/I_data_add_4 [6]) );
  ADD32 \u_decoder/fir_filter/add_298/U1_7  ( .A(
        \u_decoder/fir_filter/I_data_mult_4_buff [7]), .B(
        \u_decoder/fir_filter/I_data_add_5_buff [7]), .CI(
        \u_decoder/fir_filter/add_298/carry [7]), .CO(
        \u_decoder/fir_filter/add_298/carry [8]), .S(
        \u_decoder/fir_filter/I_data_add_4 [7]) );
  ADD32 \u_decoder/fir_filter/add_298/U1_8  ( .A(
        \u_decoder/fir_filter/I_data_mult_4_buff [8]), .B(
        \u_decoder/fir_filter/I_data_add_5_buff [8]), .CI(
        \u_decoder/fir_filter/add_298/carry [8]), .CO(
        \u_decoder/fir_filter/add_298/carry [9]), .S(
        \u_decoder/fir_filter/I_data_add_4 [8]) );
  ADD32 \u_decoder/fir_filter/add_298/U1_9  ( .A(
        \u_decoder/fir_filter/I_data_mult_4_buff [9]), .B(
        \u_decoder/fir_filter/I_data_add_5_buff [9]), .CI(
        \u_decoder/fir_filter/add_298/carry [9]), .CO(
        \u_decoder/fir_filter/add_298/carry [10]), .S(
        \u_decoder/fir_filter/I_data_add_4 [9]) );
  ADD32 \u_decoder/fir_filter/add_298/U1_10  ( .A(
        \u_decoder/fir_filter/I_data_mult_4_buff [10]), .B(
        \u_decoder/fir_filter/I_data_add_5_buff [10]), .CI(
        \u_decoder/fir_filter/add_298/carry [10]), .CO(
        \u_decoder/fir_filter/add_298/carry [11]), .S(
        \u_decoder/fir_filter/I_data_add_4 [10]) );
  ADD32 \u_decoder/fir_filter/add_298/U1_11  ( .A(
        \u_decoder/fir_filter/I_data_mult_4_buff [11]), .B(
        \u_decoder/fir_filter/I_data_add_5_buff [11]), .CI(
        \u_decoder/fir_filter/add_298/carry [11]), .CO(
        \u_decoder/fir_filter/add_298/carry [12]), .S(
        \u_decoder/fir_filter/I_data_add_4 [11]) );
  ADD32 \u_decoder/fir_filter/add_298/U1_12  ( .A(
        \u_decoder/fir_filter/I_data_mult_4_buff [12]), .B(
        \u_decoder/fir_filter/I_data_add_5_buff [12]), .CI(
        \u_decoder/fir_filter/add_298/carry [12]), .CO(
        \u_decoder/fir_filter/add_298/carry [13]), .S(
        \u_decoder/fir_filter/I_data_add_4 [12]) );
  ADD32 \u_decoder/fir_filter/add_298/U1_13  ( .A(
        \u_decoder/fir_filter/I_data_mult_4_buff [13]), .B(
        \u_decoder/fir_filter/I_data_add_5_buff [13]), .CI(
        \u_decoder/fir_filter/add_298/carry [13]), .CO(
        \u_decoder/fir_filter/add_298/carry [14]), .S(
        \u_decoder/fir_filter/I_data_add_4 [13]) );
  ADD32 \u_decoder/fir_filter/add_299/U1_1  ( .A(
        \u_decoder/fir_filter/I_data_mult_5_buff [1]), .B(
        \u_decoder/fir_filter/I_data_add_6_buff [1]), .CI(
        \u_decoder/fir_filter/add_299/carry [1]), .CO(
        \u_decoder/fir_filter/add_299/carry [2]), .S(
        \u_decoder/fir_filter/I_data_add_5 [1]) );
  ADD32 \u_decoder/fir_filter/add_299/U1_2  ( .A(
        \u_decoder/fir_filter/I_data_mult_5_buff [2]), .B(
        \u_decoder/fir_filter/I_data_add_6_buff [2]), .CI(
        \u_decoder/fir_filter/add_299/carry [2]), .CO(
        \u_decoder/fir_filter/add_299/carry [3]), .S(
        \u_decoder/fir_filter/I_data_add_5 [2]) );
  ADD32 \u_decoder/fir_filter/add_299/U1_3  ( .A(
        \u_decoder/fir_filter/I_data_mult_5_buff [3]), .B(
        \u_decoder/fir_filter/I_data_add_6_buff [3]), .CI(
        \u_decoder/fir_filter/add_299/carry [3]), .CO(
        \u_decoder/fir_filter/add_299/carry [4]), .S(
        \u_decoder/fir_filter/I_data_add_5 [3]) );
  ADD32 \u_decoder/fir_filter/add_299/U1_4  ( .A(
        \u_decoder/fir_filter/I_data_mult_5_buff [4]), .B(
        \u_decoder/fir_filter/I_data_add_6_buff [4]), .CI(
        \u_decoder/fir_filter/add_299/carry [4]), .CO(
        \u_decoder/fir_filter/add_299/carry [5]), .S(
        \u_decoder/fir_filter/I_data_add_5 [4]) );
  ADD32 \u_decoder/fir_filter/add_299/U1_5  ( .A(
        \u_decoder/fir_filter/I_data_mult_5_buff [5]), .B(
        \u_decoder/fir_filter/I_data_add_6_buff [5]), .CI(
        \u_decoder/fir_filter/add_299/carry [5]), .CO(
        \u_decoder/fir_filter/add_299/carry [6]), .S(
        \u_decoder/fir_filter/I_data_add_5 [5]) );
  ADD32 \u_decoder/fir_filter/add_299/U1_6  ( .A(
        \u_decoder/fir_filter/I_data_mult_5_buff [6]), .B(
        \u_decoder/fir_filter/I_data_add_6_buff [6]), .CI(
        \u_decoder/fir_filter/add_299/carry [6]), .CO(
        \u_decoder/fir_filter/add_299/carry [7]), .S(
        \u_decoder/fir_filter/I_data_add_5 [6]) );
  ADD32 \u_decoder/fir_filter/add_299/U1_7  ( .A(
        \u_decoder/fir_filter/I_data_mult_5_buff [7]), .B(
        \u_decoder/fir_filter/I_data_add_6_buff [7]), .CI(
        \u_decoder/fir_filter/add_299/carry [7]), .CO(
        \u_decoder/fir_filter/add_299/carry [8]), .S(
        \u_decoder/fir_filter/I_data_add_5 [7]) );
  ADD32 \u_decoder/fir_filter/add_299/U1_8  ( .A(
        \u_decoder/fir_filter/I_data_mult_5_buff [8]), .B(
        \u_decoder/fir_filter/I_data_add_6_buff [8]), .CI(
        \u_decoder/fir_filter/add_299/carry [8]), .CO(
        \u_decoder/fir_filter/add_299/carry [9]), .S(
        \u_decoder/fir_filter/I_data_add_5 [8]) );
  ADD32 \u_decoder/fir_filter/add_299/U1_9  ( .A(
        \u_decoder/fir_filter/I_data_mult_5_buff [9]), .B(
        \u_decoder/fir_filter/I_data_add_6_buff [9]), .CI(
        \u_decoder/fir_filter/add_299/carry [9]), .CO(
        \u_decoder/fir_filter/add_299/carry [10]), .S(
        \u_decoder/fir_filter/I_data_add_5 [9]) );
  ADD32 \u_decoder/fir_filter/add_299/U1_10  ( .A(
        \u_decoder/fir_filter/I_data_mult_5_buff [10]), .B(
        \u_decoder/fir_filter/I_data_add_6_buff [10]), .CI(
        \u_decoder/fir_filter/add_299/carry [10]), .CO(
        \u_decoder/fir_filter/add_299/carry [11]), .S(
        \u_decoder/fir_filter/I_data_add_5 [10]) );
  ADD32 \u_decoder/fir_filter/add_299/U1_11  ( .A(
        \u_decoder/fir_filter/I_data_mult_5_buff [11]), .B(
        \u_decoder/fir_filter/I_data_add_6_buff [11]), .CI(
        \u_decoder/fir_filter/add_299/carry [11]), .CO(
        \u_decoder/fir_filter/add_299/carry [12]), .S(
        \u_decoder/fir_filter/I_data_add_5 [11]) );
  ADD32 \u_decoder/fir_filter/add_299/U1_12  ( .A(
        \u_decoder/fir_filter/I_data_mult_5_buff [12]), .B(
        \u_decoder/fir_filter/I_data_add_6_buff [12]), .CI(
        \u_decoder/fir_filter/add_299/carry [12]), .CO(
        \u_decoder/fir_filter/add_299/carry [13]), .S(
        \u_decoder/fir_filter/I_data_add_5 [12]) );
  ADD32 \u_decoder/fir_filter/add_299/U1_13  ( .A(
        \u_decoder/fir_filter/I_data_mult_5_buff [13]), .B(
        \u_decoder/fir_filter/I_data_add_6_buff [13]), .CI(
        \u_decoder/fir_filter/add_299/carry [13]), .CO(
        \u_decoder/fir_filter/add_299/carry [14]), .S(
        \u_decoder/fir_filter/I_data_add_5 [13]) );
  ADD32 \u_decoder/fir_filter/add_300/U1_1  ( .A(
        \u_decoder/fir_filter/I_data_mult_6_buff [1]), .B(
        \u_decoder/fir_filter/I_data_add_7_buff [1]), .CI(
        \u_decoder/fir_filter/add_300/carry [1]), .CO(
        \u_decoder/fir_filter/add_300/carry [2]), .S(
        \u_decoder/fir_filter/I_data_add_6 [1]) );
  ADD32 \u_decoder/fir_filter/add_300/U1_2  ( .A(
        \u_decoder/fir_filter/I_data_mult_6_buff [2]), .B(
        \u_decoder/fir_filter/I_data_add_7_buff [2]), .CI(
        \u_decoder/fir_filter/add_300/carry [2]), .CO(
        \u_decoder/fir_filter/add_300/carry [3]), .S(
        \u_decoder/fir_filter/I_data_add_6 [2]) );
  ADD32 \u_decoder/fir_filter/add_300/U1_3  ( .A(
        \u_decoder/fir_filter/I_data_mult_6_buff [3]), .B(
        \u_decoder/fir_filter/I_data_add_7_buff [3]), .CI(
        \u_decoder/fir_filter/add_300/carry [3]), .CO(
        \u_decoder/fir_filter/add_300/carry [4]), .S(
        \u_decoder/fir_filter/I_data_add_6 [3]) );
  ADD32 \u_decoder/fir_filter/add_300/U1_4  ( .A(
        \u_decoder/fir_filter/I_data_mult_6_buff [4]), .B(
        \u_decoder/fir_filter/I_data_add_7_buff [4]), .CI(
        \u_decoder/fir_filter/add_300/carry [4]), .CO(
        \u_decoder/fir_filter/add_300/carry [5]), .S(
        \u_decoder/fir_filter/I_data_add_6 [4]) );
  ADD32 \u_decoder/fir_filter/add_300/U1_5  ( .A(
        \u_decoder/fir_filter/I_data_mult_6_buff [5]), .B(
        \u_decoder/fir_filter/I_data_add_7_buff [5]), .CI(
        \u_decoder/fir_filter/add_300/carry [5]), .CO(
        \u_decoder/fir_filter/add_300/carry [6]), .S(
        \u_decoder/fir_filter/I_data_add_6 [5]) );
  ADD32 \u_decoder/fir_filter/add_300/U1_6  ( .A(
        \u_decoder/fir_filter/I_data_mult_6_buff [6]), .B(
        \u_decoder/fir_filter/I_data_add_7_buff [6]), .CI(
        \u_decoder/fir_filter/add_300/carry [6]), .CO(
        \u_decoder/fir_filter/add_300/carry [7]), .S(
        \u_decoder/fir_filter/I_data_add_6 [6]) );
  ADD32 \u_decoder/fir_filter/add_300/U1_7  ( .A(
        \u_decoder/fir_filter/I_data_mult_6_buff [7]), .B(
        \u_decoder/fir_filter/I_data_add_7_buff [7]), .CI(
        \u_decoder/fir_filter/add_300/carry [7]), .CO(
        \u_decoder/fir_filter/add_300/carry [8]), .S(
        \u_decoder/fir_filter/I_data_add_6 [7]) );
  ADD32 \u_decoder/fir_filter/add_300/U1_8  ( .A(
        \u_decoder/fir_filter/I_data_mult_6_buff [8]), .B(
        \u_decoder/fir_filter/I_data_add_7_buff [8]), .CI(
        \u_decoder/fir_filter/add_300/carry [8]), .CO(
        \u_decoder/fir_filter/add_300/carry [9]), .S(
        \u_decoder/fir_filter/I_data_add_6 [8]) );
  ADD32 \u_decoder/fir_filter/add_300/U1_9  ( .A(
        \u_decoder/fir_filter/I_data_mult_6_buff [9]), .B(
        \u_decoder/fir_filter/I_data_add_7_buff [9]), .CI(
        \u_decoder/fir_filter/add_300/carry [9]), .CO(
        \u_decoder/fir_filter/add_300/carry [10]), .S(
        \u_decoder/fir_filter/I_data_add_6 [9]) );
  ADD32 \u_decoder/fir_filter/add_300/U1_10  ( .A(
        \u_decoder/fir_filter/I_data_mult_6_buff [10]), .B(
        \u_decoder/fir_filter/I_data_add_7_buff [10]), .CI(
        \u_decoder/fir_filter/add_300/carry [10]), .CO(
        \u_decoder/fir_filter/add_300/carry [11]), .S(
        \u_decoder/fir_filter/I_data_add_6 [10]) );
  ADD32 \u_decoder/fir_filter/add_300/U1_11  ( .A(
        \u_decoder/fir_filter/I_data_mult_6_buff [11]), .B(
        \u_decoder/fir_filter/I_data_add_7_buff [11]), .CI(
        \u_decoder/fir_filter/add_300/carry [11]), .CO(
        \u_decoder/fir_filter/add_300/carry [12]), .S(
        \u_decoder/fir_filter/I_data_add_6 [11]) );
  ADD32 \u_decoder/fir_filter/add_300/U1_12  ( .A(
        \u_decoder/fir_filter/I_data_mult_6_buff [12]), .B(
        \u_decoder/fir_filter/I_data_add_7_buff [12]), .CI(
        \u_decoder/fir_filter/add_300/carry [12]), .CO(
        \u_decoder/fir_filter/add_300/carry [13]), .S(
        \u_decoder/fir_filter/I_data_add_6 [12]) );
  ADD32 \u_decoder/fir_filter/add_300/U1_13  ( .A(
        \u_decoder/fir_filter/I_data_mult_6_buff [13]), .B(
        \u_decoder/fir_filter/I_data_add_7_buff [13]), .CI(
        \u_decoder/fir_filter/add_300/carry [13]), .CO(
        \u_decoder/fir_filter/add_300/carry [14]), .S(
        \u_decoder/fir_filter/I_data_add_6 [13]) );
  ADD32 \u_decoder/fir_filter/add_301/U1_1  ( .A(
        \u_decoder/fir_filter/I_data_mult_7_buff [1]), .B(
        \u_decoder/fir_filter/I_data_mult_8_buff [1]), .CI(
        \u_decoder/fir_filter/add_301/carry [1]), .CO(
        \u_decoder/fir_filter/add_301/carry [2]), .S(
        \u_decoder/fir_filter/I_data_add_7 [1]) );
  ADD32 \u_decoder/fir_filter/add_301/U1_2  ( .A(
        \u_decoder/fir_filter/I_data_mult_7_buff [2]), .B(
        \u_decoder/fir_filter/I_data_mult_8_buff [2]), .CI(
        \u_decoder/fir_filter/add_301/carry [2]), .CO(
        \u_decoder/fir_filter/add_301/carry [3]), .S(
        \u_decoder/fir_filter/I_data_add_7 [2]) );
  ADD32 \u_decoder/fir_filter/add_301/U1_3  ( .A(
        \u_decoder/fir_filter/I_data_mult_7_buff [3]), .B(
        \u_decoder/fir_filter/I_data_mult_8_buff [3]), .CI(
        \u_decoder/fir_filter/add_301/carry [3]), .CO(
        \u_decoder/fir_filter/add_301/carry [4]), .S(
        \u_decoder/fir_filter/I_data_add_7 [3]) );
  ADD32 \u_decoder/fir_filter/add_301/U1_4  ( .A(
        \u_decoder/fir_filter/I_data_mult_7_buff [4]), .B(
        \u_decoder/fir_filter/I_data_mult_8_buff [4]), .CI(
        \u_decoder/fir_filter/add_301/carry [4]), .CO(
        \u_decoder/fir_filter/add_301/carry [5]), .S(
        \u_decoder/fir_filter/I_data_add_7 [4]) );
  ADD32 \u_decoder/fir_filter/add_301/U1_5  ( .A(
        \u_decoder/fir_filter/I_data_mult_7_buff [5]), .B(
        \u_decoder/fir_filter/I_data_mult_8_buff [5]), .CI(
        \u_decoder/fir_filter/add_301/carry [5]), .CO(
        \u_decoder/fir_filter/add_301/carry [6]), .S(
        \u_decoder/fir_filter/I_data_add_7 [5]) );
  ADD32 \u_decoder/fir_filter/add_301/U1_6  ( .A(
        \u_decoder/fir_filter/I_data_mult_7_buff [6]), .B(
        \u_decoder/fir_filter/I_data_mult_8_buff [6]), .CI(
        \u_decoder/fir_filter/add_301/carry [6]), .CO(
        \u_decoder/fir_filter/add_301/carry [7]), .S(
        \u_decoder/fir_filter/I_data_add_7 [6]) );
  ADD32 \u_decoder/fir_filter/add_301/U1_7  ( .A(
        \u_decoder/fir_filter/I_data_mult_7_buff [7]), .B(
        \u_decoder/fir_filter/I_data_mult_8_buff [7]), .CI(
        \u_decoder/fir_filter/add_301/carry [7]), .CO(
        \u_decoder/fir_filter/add_301/carry [8]), .S(
        \u_decoder/fir_filter/I_data_add_7 [7]) );
  ADD32 \u_decoder/fir_filter/add_301/U1_8  ( .A(
        \u_decoder/fir_filter/I_data_mult_7_buff [8]), .B(
        \u_decoder/fir_filter/I_data_mult_8_buff [8]), .CI(
        \u_decoder/fir_filter/add_301/carry [8]), .CO(
        \u_decoder/fir_filter/add_301/carry [9]), .S(
        \u_decoder/fir_filter/I_data_add_7 [8]) );
  ADD32 \u_decoder/fir_filter/add_301/U1_9  ( .A(
        \u_decoder/fir_filter/I_data_mult_7_buff [9]), .B(
        \u_decoder/fir_filter/I_data_mult_8_buff [9]), .CI(
        \u_decoder/fir_filter/add_301/carry [9]), .CO(
        \u_decoder/fir_filter/add_301/carry [10]), .S(
        \u_decoder/fir_filter/I_data_add_7 [9]) );
  ADD32 \u_decoder/fir_filter/add_301/U1_10  ( .A(
        \u_decoder/fir_filter/I_data_mult_7_buff [10]), .B(
        \u_decoder/fir_filter/I_data_mult_8_buff [10]), .CI(
        \u_decoder/fir_filter/add_301/carry [10]), .CO(
        \u_decoder/fir_filter/add_301/carry [11]), .S(
        \u_decoder/fir_filter/I_data_add_7 [10]) );
  ADD32 \u_decoder/fir_filter/add_301/U1_11  ( .A(
        \u_decoder/fir_filter/I_data_mult_7_buff [11]), .B(
        \u_decoder/fir_filter/I_data_mult_8_buff [11]), .CI(
        \u_decoder/fir_filter/add_301/carry [11]), .CO(
        \u_decoder/fir_filter/add_301/carry [12]), .S(
        \u_decoder/fir_filter/I_data_add_7 [11]) );
  ADD32 \u_decoder/fir_filter/add_301/U1_12  ( .A(
        \u_decoder/fir_filter/I_data_mult_7_buff [12]), .B(
        \u_decoder/fir_filter/I_data_mult_8_buff [12]), .CI(
        \u_decoder/fir_filter/add_301/carry [12]), .CO(
        \u_decoder/fir_filter/add_301/carry [13]), .S(
        \u_decoder/fir_filter/I_data_add_7 [12]) );
  ADD32 \u_decoder/fir_filter/add_301/U1_13  ( .A(
        \u_decoder/fir_filter/I_data_mult_7_buff [13]), .B(
        \u_decoder/fir_filter/I_data_mult_8_buff [13]), .CI(
        \u_decoder/fir_filter/add_301/carry [13]), .CO(
        \u_decoder/fir_filter/add_301/carry [14]), .S(
        \u_decoder/fir_filter/I_data_add_7 [13]) );
  ADD32 \u_decoder/fir_filter/add_326/U1_11  ( .A(
        \u_decoder/fir_filter/Q_data_mult_0_buff [11]), .B(
        \u_decoder/fir_filter/Q_data_add_1_buff [11]), .CI(
        \u_decoder/fir_filter/add_326/carry [11]), .CO(
        \u_decoder/fir_filter/add_326/carry [12]), .S(
        \u_decoder/fir_filter/Q_data_add_0 [11]) );
  ADD32 \u_decoder/fir_filter/add_326/U1_12  ( .A(
        \u_decoder/fir_filter/Q_data_mult_0_buff [12]), .B(
        \u_decoder/fir_filter/Q_data_add_1_buff [12]), .CI(
        \u_decoder/fir_filter/add_326/carry [12]), .CO(
        \u_decoder/fir_filter/add_326/carry [13]), .S(
        \u_decoder/fir_filter/Q_data_add_0 [12]) );
  ADD32 \u_decoder/fir_filter/add_326/U1_13  ( .A(
        \u_decoder/fir_filter/Q_data_mult_0_buff [13]), .B(
        \u_decoder/fir_filter/Q_data_add_1_buff [13]), .CI(
        \u_decoder/fir_filter/add_326/carry [13]), .CO(
        \u_decoder/fir_filter/add_326/carry [14]), .S(
        \u_decoder/fir_filter/Q_data_add_0 [13]) );
  ADD32 \u_decoder/fir_filter/add_327/U1_1  ( .A(
        \u_decoder/fir_filter/Q_data_mult_1_buff [1]), .B(
        \u_decoder/fir_filter/Q_data_add_2_buff [1]), .CI(
        \u_decoder/fir_filter/add_327/carry [1]), .CO(
        \u_decoder/fir_filter/add_327/carry [2]), .S(
        \u_decoder/fir_filter/Q_data_add_1 [1]) );
  ADD32 \u_decoder/fir_filter/add_327/U1_2  ( .A(
        \u_decoder/fir_filter/Q_data_mult_1_buff [2]), .B(
        \u_decoder/fir_filter/Q_data_add_2_buff [2]), .CI(
        \u_decoder/fir_filter/add_327/carry [2]), .CO(
        \u_decoder/fir_filter/add_327/carry [3]), .S(
        \u_decoder/fir_filter/Q_data_add_1 [2]) );
  ADD32 \u_decoder/fir_filter/add_327/U1_3  ( .A(
        \u_decoder/fir_filter/Q_data_mult_1_buff [3]), .B(
        \u_decoder/fir_filter/Q_data_add_2_buff [3]), .CI(
        \u_decoder/fir_filter/add_327/carry [3]), .CO(
        \u_decoder/fir_filter/add_327/carry [4]), .S(
        \u_decoder/fir_filter/Q_data_add_1 [3]) );
  ADD32 \u_decoder/fir_filter/add_327/U1_4  ( .A(
        \u_decoder/fir_filter/Q_data_mult_1_buff [4]), .B(
        \u_decoder/fir_filter/Q_data_add_2_buff [4]), .CI(
        \u_decoder/fir_filter/add_327/carry [4]), .CO(
        \u_decoder/fir_filter/add_327/carry [5]), .S(
        \u_decoder/fir_filter/Q_data_add_1 [4]) );
  ADD32 \u_decoder/fir_filter/add_327/U1_5  ( .A(
        \u_decoder/fir_filter/Q_data_mult_1_buff [5]), .B(
        \u_decoder/fir_filter/Q_data_add_2_buff [5]), .CI(
        \u_decoder/fir_filter/add_327/carry [5]), .CO(
        \u_decoder/fir_filter/add_327/carry [6]), .S(
        \u_decoder/fir_filter/Q_data_add_1 [5]) );
  ADD32 \u_decoder/fir_filter/add_327/U1_6  ( .A(
        \u_decoder/fir_filter/Q_data_mult_1_buff [6]), .B(
        \u_decoder/fir_filter/Q_data_add_2_buff [6]), .CI(
        \u_decoder/fir_filter/add_327/carry [6]), .CO(
        \u_decoder/fir_filter/add_327/carry [7]), .S(
        \u_decoder/fir_filter/Q_data_add_1 [6]) );
  ADD32 \u_decoder/fir_filter/add_327/U1_7  ( .A(
        \u_decoder/fir_filter/Q_data_mult_1_buff [7]), .B(
        \u_decoder/fir_filter/Q_data_add_2_buff [7]), .CI(
        \u_decoder/fir_filter/add_327/carry [7]), .CO(
        \u_decoder/fir_filter/add_327/carry [8]), .S(
        \u_decoder/fir_filter/Q_data_add_1 [7]) );
  ADD32 \u_decoder/fir_filter/add_327/U1_8  ( .A(
        \u_decoder/fir_filter/Q_data_mult_1_buff [8]), .B(
        \u_decoder/fir_filter/Q_data_add_2_buff [8]), .CI(
        \u_decoder/fir_filter/add_327/carry [8]), .CO(
        \u_decoder/fir_filter/add_327/carry [9]), .S(
        \u_decoder/fir_filter/Q_data_add_1 [8]) );
  ADD32 \u_decoder/fir_filter/add_327/U1_9  ( .A(
        \u_decoder/fir_filter/Q_data_mult_1_buff [9]), .B(
        \u_decoder/fir_filter/Q_data_add_2_buff [9]), .CI(
        \u_decoder/fir_filter/add_327/carry [9]), .CO(
        \u_decoder/fir_filter/add_327/carry [10]), .S(
        \u_decoder/fir_filter/Q_data_add_1 [9]) );
  ADD32 \u_decoder/fir_filter/add_327/U1_10  ( .A(
        \u_decoder/fir_filter/Q_data_mult_1_buff [10]), .B(
        \u_decoder/fir_filter/Q_data_add_2_buff [10]), .CI(
        \u_decoder/fir_filter/add_327/carry [10]), .CO(
        \u_decoder/fir_filter/add_327/carry [11]), .S(
        \u_decoder/fir_filter/Q_data_add_1 [10]) );
  ADD32 \u_decoder/fir_filter/add_327/U1_11  ( .A(
        \u_decoder/fir_filter/Q_data_mult_1_buff [11]), .B(
        \u_decoder/fir_filter/Q_data_add_2_buff [11]), .CI(
        \u_decoder/fir_filter/add_327/carry [11]), .CO(
        \u_decoder/fir_filter/add_327/carry [12]), .S(
        \u_decoder/fir_filter/Q_data_add_1 [11]) );
  ADD32 \u_decoder/fir_filter/add_327/U1_12  ( .A(
        \u_decoder/fir_filter/Q_data_mult_1_buff [12]), .B(
        \u_decoder/fir_filter/Q_data_add_2_buff [12]), .CI(
        \u_decoder/fir_filter/add_327/carry [12]), .CO(
        \u_decoder/fir_filter/add_327/carry [13]), .S(
        \u_decoder/fir_filter/Q_data_add_1 [12]) );
  ADD32 \u_decoder/fir_filter/add_327/U1_13  ( .A(
        \u_decoder/fir_filter/Q_data_mult_1_buff [13]), .B(
        \u_decoder/fir_filter/Q_data_add_2_buff [13]), .CI(
        \u_decoder/fir_filter/add_327/carry [13]), .CO(
        \u_decoder/fir_filter/add_327/carry [14]), .S(
        \u_decoder/fir_filter/Q_data_add_1 [13]) );
  ADD32 \u_decoder/fir_filter/add_328/U1_1  ( .A(
        \u_decoder/fir_filter/Q_data_mult_2_buff [1]), .B(
        \u_decoder/fir_filter/Q_data_add_3_buff [1]), .CI(
        \u_decoder/fir_filter/add_328/carry [1]), .CO(
        \u_decoder/fir_filter/add_328/carry [2]), .S(
        \u_decoder/fir_filter/Q_data_add_2 [1]) );
  ADD32 \u_decoder/fir_filter/add_328/U1_2  ( .A(
        \u_decoder/fir_filter/Q_data_mult_2_buff [2]), .B(
        \u_decoder/fir_filter/Q_data_add_3_buff [2]), .CI(
        \u_decoder/fir_filter/add_328/carry [2]), .CO(
        \u_decoder/fir_filter/add_328/carry [3]), .S(
        \u_decoder/fir_filter/Q_data_add_2 [2]) );
  ADD32 \u_decoder/fir_filter/add_328/U1_3  ( .A(
        \u_decoder/fir_filter/Q_data_mult_2_buff [3]), .B(
        \u_decoder/fir_filter/Q_data_add_3_buff [3]), .CI(
        \u_decoder/fir_filter/add_328/carry [3]), .CO(
        \u_decoder/fir_filter/add_328/carry [4]), .S(
        \u_decoder/fir_filter/Q_data_add_2 [3]) );
  ADD32 \u_decoder/fir_filter/add_328/U1_4  ( .A(
        \u_decoder/fir_filter/Q_data_mult_2_buff [4]), .B(
        \u_decoder/fir_filter/Q_data_add_3_buff [4]), .CI(
        \u_decoder/fir_filter/add_328/carry [4]), .CO(
        \u_decoder/fir_filter/add_328/carry [5]), .S(
        \u_decoder/fir_filter/Q_data_add_2 [4]) );
  ADD32 \u_decoder/fir_filter/add_328/U1_5  ( .A(
        \u_decoder/fir_filter/Q_data_mult_2_buff [5]), .B(
        \u_decoder/fir_filter/Q_data_add_3_buff [5]), .CI(
        \u_decoder/fir_filter/add_328/carry [5]), .CO(
        \u_decoder/fir_filter/add_328/carry [6]), .S(
        \u_decoder/fir_filter/Q_data_add_2 [5]) );
  ADD32 \u_decoder/fir_filter/add_328/U1_6  ( .A(
        \u_decoder/fir_filter/Q_data_mult_2_buff [6]), .B(
        \u_decoder/fir_filter/Q_data_add_3_buff [6]), .CI(
        \u_decoder/fir_filter/add_328/carry [6]), .CO(
        \u_decoder/fir_filter/add_328/carry [7]), .S(
        \u_decoder/fir_filter/Q_data_add_2 [6]) );
  ADD32 \u_decoder/fir_filter/add_328/U1_7  ( .A(
        \u_decoder/fir_filter/Q_data_mult_2_buff [7]), .B(
        \u_decoder/fir_filter/Q_data_add_3_buff [7]), .CI(
        \u_decoder/fir_filter/add_328/carry [7]), .CO(
        \u_decoder/fir_filter/add_328/carry [8]), .S(
        \u_decoder/fir_filter/Q_data_add_2 [7]) );
  ADD32 \u_decoder/fir_filter/add_328/U1_8  ( .A(
        \u_decoder/fir_filter/Q_data_mult_2_buff [8]), .B(
        \u_decoder/fir_filter/Q_data_add_3_buff [8]), .CI(
        \u_decoder/fir_filter/add_328/carry [8]), .CO(
        \u_decoder/fir_filter/add_328/carry [9]), .S(
        \u_decoder/fir_filter/Q_data_add_2 [8]) );
  ADD32 \u_decoder/fir_filter/add_328/U1_9  ( .A(
        \u_decoder/fir_filter/Q_data_mult_2_buff [9]), .B(
        \u_decoder/fir_filter/Q_data_add_3_buff [9]), .CI(
        \u_decoder/fir_filter/add_328/carry [9]), .CO(
        \u_decoder/fir_filter/add_328/carry [10]), .S(
        \u_decoder/fir_filter/Q_data_add_2 [9]) );
  ADD32 \u_decoder/fir_filter/add_328/U1_10  ( .A(
        \u_decoder/fir_filter/Q_data_mult_2_buff [10]), .B(
        \u_decoder/fir_filter/Q_data_add_3_buff [10]), .CI(
        \u_decoder/fir_filter/add_328/carry [10]), .CO(
        \u_decoder/fir_filter/add_328/carry [11]), .S(
        \u_decoder/fir_filter/Q_data_add_2 [10]) );
  ADD32 \u_decoder/fir_filter/add_328/U1_11  ( .A(
        \u_decoder/fir_filter/Q_data_mult_2_buff [11]), .B(
        \u_decoder/fir_filter/Q_data_add_3_buff [11]), .CI(
        \u_decoder/fir_filter/add_328/carry [11]), .CO(
        \u_decoder/fir_filter/add_328/carry [12]), .S(
        \u_decoder/fir_filter/Q_data_add_2 [11]) );
  ADD32 \u_decoder/fir_filter/add_328/U1_12  ( .A(
        \u_decoder/fir_filter/Q_data_mult_2_buff [12]), .B(
        \u_decoder/fir_filter/Q_data_add_3_buff [12]), .CI(
        \u_decoder/fir_filter/add_328/carry [12]), .CO(
        \u_decoder/fir_filter/add_328/carry [13]), .S(
        \u_decoder/fir_filter/Q_data_add_2 [12]) );
  ADD32 \u_decoder/fir_filter/add_328/U1_13  ( .A(
        \u_decoder/fir_filter/Q_data_mult_2_buff [13]), .B(
        \u_decoder/fir_filter/Q_data_add_3_buff [13]), .CI(
        \u_decoder/fir_filter/add_328/carry [13]), .CO(
        \u_decoder/fir_filter/add_328/carry [14]), .S(
        \u_decoder/fir_filter/Q_data_add_2 [13]) );
  ADD32 \u_decoder/fir_filter/add_329/U1_1  ( .A(
        \u_decoder/fir_filter/Q_data_mult_3_buff [1]), .B(
        \u_decoder/fir_filter/Q_data_add_4_buff [1]), .CI(
        \u_decoder/fir_filter/add_329/carry [1]), .CO(
        \u_decoder/fir_filter/add_329/carry [2]), .S(
        \u_decoder/fir_filter/Q_data_add_3 [1]) );
  ADD32 \u_decoder/fir_filter/add_329/U1_2  ( .A(
        \u_decoder/fir_filter/Q_data_mult_3_buff [2]), .B(
        \u_decoder/fir_filter/Q_data_add_4_buff [2]), .CI(
        \u_decoder/fir_filter/add_329/carry [2]), .CO(
        \u_decoder/fir_filter/add_329/carry [3]), .S(
        \u_decoder/fir_filter/Q_data_add_3 [2]) );
  ADD32 \u_decoder/fir_filter/add_329/U1_3  ( .A(
        \u_decoder/fir_filter/Q_data_mult_3_buff [3]), .B(
        \u_decoder/fir_filter/Q_data_add_4_buff [3]), .CI(
        \u_decoder/fir_filter/add_329/carry [3]), .CO(
        \u_decoder/fir_filter/add_329/carry [4]), .S(
        \u_decoder/fir_filter/Q_data_add_3 [3]) );
  ADD32 \u_decoder/fir_filter/add_329/U1_4  ( .A(
        \u_decoder/fir_filter/Q_data_mult_3_buff [4]), .B(
        \u_decoder/fir_filter/Q_data_add_4_buff [4]), .CI(
        \u_decoder/fir_filter/add_329/carry [4]), .CO(
        \u_decoder/fir_filter/add_329/carry [5]), .S(
        \u_decoder/fir_filter/Q_data_add_3 [4]) );
  ADD32 \u_decoder/fir_filter/add_329/U1_5  ( .A(
        \u_decoder/fir_filter/Q_data_mult_3_buff [5]), .B(
        \u_decoder/fir_filter/Q_data_add_4_buff [5]), .CI(
        \u_decoder/fir_filter/add_329/carry [5]), .CO(
        \u_decoder/fir_filter/add_329/carry [6]), .S(
        \u_decoder/fir_filter/Q_data_add_3 [5]) );
  ADD32 \u_decoder/fir_filter/add_329/U1_6  ( .A(
        \u_decoder/fir_filter/Q_data_mult_3_buff [6]), .B(
        \u_decoder/fir_filter/Q_data_add_4_buff [6]), .CI(
        \u_decoder/fir_filter/add_329/carry [6]), .CO(
        \u_decoder/fir_filter/add_329/carry [7]), .S(
        \u_decoder/fir_filter/Q_data_add_3 [6]) );
  ADD32 \u_decoder/fir_filter/add_329/U1_7  ( .A(
        \u_decoder/fir_filter/Q_data_mult_3_buff [7]), .B(
        \u_decoder/fir_filter/Q_data_add_4_buff [7]), .CI(
        \u_decoder/fir_filter/add_329/carry [7]), .CO(
        \u_decoder/fir_filter/add_329/carry [8]), .S(
        \u_decoder/fir_filter/Q_data_add_3 [7]) );
  ADD32 \u_decoder/fir_filter/add_329/U1_8  ( .A(
        \u_decoder/fir_filter/Q_data_mult_3_buff [8]), .B(
        \u_decoder/fir_filter/Q_data_add_4_buff [8]), .CI(
        \u_decoder/fir_filter/add_329/carry [8]), .CO(
        \u_decoder/fir_filter/add_329/carry [9]), .S(
        \u_decoder/fir_filter/Q_data_add_3 [8]) );
  ADD32 \u_decoder/fir_filter/add_329/U1_9  ( .A(
        \u_decoder/fir_filter/Q_data_mult_3_buff [9]), .B(
        \u_decoder/fir_filter/Q_data_add_4_buff [9]), .CI(
        \u_decoder/fir_filter/add_329/carry [9]), .CO(
        \u_decoder/fir_filter/add_329/carry [10]), .S(
        \u_decoder/fir_filter/Q_data_add_3 [9]) );
  ADD32 \u_decoder/fir_filter/add_329/U1_10  ( .A(
        \u_decoder/fir_filter/Q_data_mult_3_buff [10]), .B(
        \u_decoder/fir_filter/Q_data_add_4_buff [10]), .CI(
        \u_decoder/fir_filter/add_329/carry [10]), .CO(
        \u_decoder/fir_filter/add_329/carry [11]), .S(
        \u_decoder/fir_filter/Q_data_add_3 [10]) );
  ADD32 \u_decoder/fir_filter/add_329/U1_11  ( .A(
        \u_decoder/fir_filter/Q_data_mult_3_buff [11]), .B(
        \u_decoder/fir_filter/Q_data_add_4_buff [11]), .CI(
        \u_decoder/fir_filter/add_329/carry [11]), .CO(
        \u_decoder/fir_filter/add_329/carry [12]), .S(
        \u_decoder/fir_filter/Q_data_add_3 [11]) );
  ADD32 \u_decoder/fir_filter/add_329/U1_12  ( .A(
        \u_decoder/fir_filter/Q_data_mult_3_buff [12]), .B(
        \u_decoder/fir_filter/Q_data_add_4_buff [12]), .CI(
        \u_decoder/fir_filter/add_329/carry [12]), .CO(
        \u_decoder/fir_filter/add_329/carry [13]), .S(
        \u_decoder/fir_filter/Q_data_add_3 [12]) );
  ADD32 \u_decoder/fir_filter/add_329/U1_13  ( .A(
        \u_decoder/fir_filter/Q_data_mult_3_buff [13]), .B(
        \u_decoder/fir_filter/Q_data_add_4_buff [13]), .CI(
        \u_decoder/fir_filter/add_329/carry [13]), .CO(
        \u_decoder/fir_filter/add_329/carry [14]), .S(
        \u_decoder/fir_filter/Q_data_add_3 [13]) );
  ADD32 \u_decoder/fir_filter/add_330/U1_1  ( .A(
        \u_decoder/fir_filter/Q_data_mult_4_buff [1]), .B(
        \u_decoder/fir_filter/Q_data_add_5_buff [1]), .CI(
        \u_decoder/fir_filter/add_330/carry [1]), .CO(
        \u_decoder/fir_filter/add_330/carry [2]), .S(
        \u_decoder/fir_filter/Q_data_add_4 [1]) );
  ADD32 \u_decoder/fir_filter/add_330/U1_2  ( .A(
        \u_decoder/fir_filter/Q_data_mult_4_buff [2]), .B(
        \u_decoder/fir_filter/Q_data_add_5_buff [2]), .CI(
        \u_decoder/fir_filter/add_330/carry [2]), .CO(
        \u_decoder/fir_filter/add_330/carry [3]), .S(
        \u_decoder/fir_filter/Q_data_add_4 [2]) );
  ADD32 \u_decoder/fir_filter/add_330/U1_3  ( .A(
        \u_decoder/fir_filter/Q_data_mult_4_buff [3]), .B(
        \u_decoder/fir_filter/Q_data_add_5_buff [3]), .CI(
        \u_decoder/fir_filter/add_330/carry [3]), .CO(
        \u_decoder/fir_filter/add_330/carry [4]), .S(
        \u_decoder/fir_filter/Q_data_add_4 [3]) );
  ADD32 \u_decoder/fir_filter/add_330/U1_4  ( .A(
        \u_decoder/fir_filter/Q_data_mult_4_buff [4]), .B(
        \u_decoder/fir_filter/Q_data_add_5_buff [4]), .CI(
        \u_decoder/fir_filter/add_330/carry [4]), .CO(
        \u_decoder/fir_filter/add_330/carry [5]), .S(
        \u_decoder/fir_filter/Q_data_add_4 [4]) );
  ADD32 \u_decoder/fir_filter/add_330/U1_5  ( .A(
        \u_decoder/fir_filter/Q_data_mult_4_buff [5]), .B(
        \u_decoder/fir_filter/Q_data_add_5_buff [5]), .CI(
        \u_decoder/fir_filter/add_330/carry [5]), .CO(
        \u_decoder/fir_filter/add_330/carry [6]), .S(
        \u_decoder/fir_filter/Q_data_add_4 [5]) );
  ADD32 \u_decoder/fir_filter/add_330/U1_6  ( .A(
        \u_decoder/fir_filter/Q_data_mult_4_buff [6]), .B(
        \u_decoder/fir_filter/Q_data_add_5_buff [6]), .CI(
        \u_decoder/fir_filter/add_330/carry [6]), .CO(
        \u_decoder/fir_filter/add_330/carry [7]), .S(
        \u_decoder/fir_filter/Q_data_add_4 [6]) );
  ADD32 \u_decoder/fir_filter/add_330/U1_7  ( .A(
        \u_decoder/fir_filter/Q_data_mult_4_buff [7]), .B(
        \u_decoder/fir_filter/Q_data_add_5_buff [7]), .CI(
        \u_decoder/fir_filter/add_330/carry [7]), .CO(
        \u_decoder/fir_filter/add_330/carry [8]), .S(
        \u_decoder/fir_filter/Q_data_add_4 [7]) );
  ADD32 \u_decoder/fir_filter/add_330/U1_8  ( .A(
        \u_decoder/fir_filter/Q_data_mult_4_buff [8]), .B(
        \u_decoder/fir_filter/Q_data_add_5_buff [8]), .CI(
        \u_decoder/fir_filter/add_330/carry [8]), .CO(
        \u_decoder/fir_filter/add_330/carry [9]), .S(
        \u_decoder/fir_filter/Q_data_add_4 [8]) );
  ADD32 \u_decoder/fir_filter/add_330/U1_9  ( .A(
        \u_decoder/fir_filter/Q_data_mult_4_buff [9]), .B(
        \u_decoder/fir_filter/Q_data_add_5_buff [9]), .CI(
        \u_decoder/fir_filter/add_330/carry [9]), .CO(
        \u_decoder/fir_filter/add_330/carry [10]), .S(
        \u_decoder/fir_filter/Q_data_add_4 [9]) );
  ADD32 \u_decoder/fir_filter/add_330/U1_10  ( .A(
        \u_decoder/fir_filter/Q_data_mult_4_buff [10]), .B(
        \u_decoder/fir_filter/Q_data_add_5_buff [10]), .CI(
        \u_decoder/fir_filter/add_330/carry [10]), .CO(
        \u_decoder/fir_filter/add_330/carry [11]), .S(
        \u_decoder/fir_filter/Q_data_add_4 [10]) );
  ADD32 \u_decoder/fir_filter/add_330/U1_11  ( .A(
        \u_decoder/fir_filter/Q_data_mult_4_buff [11]), .B(
        \u_decoder/fir_filter/Q_data_add_5_buff [11]), .CI(
        \u_decoder/fir_filter/add_330/carry [11]), .CO(
        \u_decoder/fir_filter/add_330/carry [12]), .S(
        \u_decoder/fir_filter/Q_data_add_4 [11]) );
  ADD32 \u_decoder/fir_filter/add_330/U1_12  ( .A(
        \u_decoder/fir_filter/Q_data_mult_4_buff [12]), .B(
        \u_decoder/fir_filter/Q_data_add_5_buff [12]), .CI(
        \u_decoder/fir_filter/add_330/carry [12]), .CO(
        \u_decoder/fir_filter/add_330/carry [13]), .S(
        \u_decoder/fir_filter/Q_data_add_4 [12]) );
  ADD32 \u_decoder/fir_filter/add_330/U1_13  ( .A(
        \u_decoder/fir_filter/Q_data_mult_4_buff [13]), .B(
        \u_decoder/fir_filter/Q_data_add_5_buff [13]), .CI(
        \u_decoder/fir_filter/add_330/carry [13]), .CO(
        \u_decoder/fir_filter/add_330/carry [14]), .S(
        \u_decoder/fir_filter/Q_data_add_4 [13]) );
  ADD32 \u_decoder/fir_filter/add_331/U1_1  ( .A(
        \u_decoder/fir_filter/Q_data_mult_5_buff [1]), .B(
        \u_decoder/fir_filter/Q_data_add_6_buff [1]), .CI(
        \u_decoder/fir_filter/add_331/carry [1]), .CO(
        \u_decoder/fir_filter/add_331/carry [2]), .S(
        \u_decoder/fir_filter/Q_data_add_5 [1]) );
  ADD32 \u_decoder/fir_filter/add_331/U1_2  ( .A(
        \u_decoder/fir_filter/Q_data_mult_5_buff [2]), .B(
        \u_decoder/fir_filter/Q_data_add_6_buff [2]), .CI(
        \u_decoder/fir_filter/add_331/carry [2]), .CO(
        \u_decoder/fir_filter/add_331/carry [3]), .S(
        \u_decoder/fir_filter/Q_data_add_5 [2]) );
  ADD32 \u_decoder/fir_filter/add_331/U1_3  ( .A(
        \u_decoder/fir_filter/Q_data_mult_5_buff [3]), .B(
        \u_decoder/fir_filter/Q_data_add_6_buff [3]), .CI(
        \u_decoder/fir_filter/add_331/carry [3]), .CO(
        \u_decoder/fir_filter/add_331/carry [4]), .S(
        \u_decoder/fir_filter/Q_data_add_5 [3]) );
  ADD32 \u_decoder/fir_filter/add_331/U1_4  ( .A(
        \u_decoder/fir_filter/Q_data_mult_5_buff [4]), .B(
        \u_decoder/fir_filter/Q_data_add_6_buff [4]), .CI(
        \u_decoder/fir_filter/add_331/carry [4]), .CO(
        \u_decoder/fir_filter/add_331/carry [5]), .S(
        \u_decoder/fir_filter/Q_data_add_5 [4]) );
  ADD32 \u_decoder/fir_filter/add_331/U1_5  ( .A(
        \u_decoder/fir_filter/Q_data_mult_5_buff [5]), .B(
        \u_decoder/fir_filter/Q_data_add_6_buff [5]), .CI(
        \u_decoder/fir_filter/add_331/carry [5]), .CO(
        \u_decoder/fir_filter/add_331/carry [6]), .S(
        \u_decoder/fir_filter/Q_data_add_5 [5]) );
  ADD32 \u_decoder/fir_filter/add_331/U1_6  ( .A(
        \u_decoder/fir_filter/Q_data_mult_5_buff [6]), .B(
        \u_decoder/fir_filter/Q_data_add_6_buff [6]), .CI(
        \u_decoder/fir_filter/add_331/carry [6]), .CO(
        \u_decoder/fir_filter/add_331/carry [7]), .S(
        \u_decoder/fir_filter/Q_data_add_5 [6]) );
  ADD32 \u_decoder/fir_filter/add_331/U1_7  ( .A(
        \u_decoder/fir_filter/Q_data_mult_5_buff [7]), .B(
        \u_decoder/fir_filter/Q_data_add_6_buff [7]), .CI(
        \u_decoder/fir_filter/add_331/carry [7]), .CO(
        \u_decoder/fir_filter/add_331/carry [8]), .S(
        \u_decoder/fir_filter/Q_data_add_5 [7]) );
  ADD32 \u_decoder/fir_filter/add_331/U1_8  ( .A(
        \u_decoder/fir_filter/Q_data_mult_5_buff [8]), .B(
        \u_decoder/fir_filter/Q_data_add_6_buff [8]), .CI(
        \u_decoder/fir_filter/add_331/carry [8]), .CO(
        \u_decoder/fir_filter/add_331/carry [9]), .S(
        \u_decoder/fir_filter/Q_data_add_5 [8]) );
  ADD32 \u_decoder/fir_filter/add_331/U1_9  ( .A(
        \u_decoder/fir_filter/Q_data_mult_5_buff [9]), .B(
        \u_decoder/fir_filter/Q_data_add_6_buff [9]), .CI(
        \u_decoder/fir_filter/add_331/carry [9]), .CO(
        \u_decoder/fir_filter/add_331/carry [10]), .S(
        \u_decoder/fir_filter/Q_data_add_5 [9]) );
  ADD32 \u_decoder/fir_filter/add_331/U1_10  ( .A(
        \u_decoder/fir_filter/Q_data_mult_5_buff [10]), .B(
        \u_decoder/fir_filter/Q_data_add_6_buff [10]), .CI(
        \u_decoder/fir_filter/add_331/carry [10]), .CO(
        \u_decoder/fir_filter/add_331/carry [11]), .S(
        \u_decoder/fir_filter/Q_data_add_5 [10]) );
  ADD32 \u_decoder/fir_filter/add_331/U1_11  ( .A(
        \u_decoder/fir_filter/Q_data_mult_5_buff [11]), .B(
        \u_decoder/fir_filter/Q_data_add_6_buff [11]), .CI(
        \u_decoder/fir_filter/add_331/carry [11]), .CO(
        \u_decoder/fir_filter/add_331/carry [12]), .S(
        \u_decoder/fir_filter/Q_data_add_5 [11]) );
  ADD32 \u_decoder/fir_filter/add_331/U1_12  ( .A(
        \u_decoder/fir_filter/Q_data_mult_5_buff [12]), .B(
        \u_decoder/fir_filter/Q_data_add_6_buff [12]), .CI(
        \u_decoder/fir_filter/add_331/carry [12]), .CO(
        \u_decoder/fir_filter/add_331/carry [13]), .S(
        \u_decoder/fir_filter/Q_data_add_5 [12]) );
  ADD32 \u_decoder/fir_filter/add_331/U1_13  ( .A(
        \u_decoder/fir_filter/Q_data_mult_5_buff [13]), .B(
        \u_decoder/fir_filter/Q_data_add_6_buff [13]), .CI(
        \u_decoder/fir_filter/add_331/carry [13]), .CO(
        \u_decoder/fir_filter/add_331/carry [14]), .S(
        \u_decoder/fir_filter/Q_data_add_5 [13]) );
  ADD32 \u_decoder/fir_filter/add_332/U1_1  ( .A(
        \u_decoder/fir_filter/Q_data_mult_6_buff [1]), .B(
        \u_decoder/fir_filter/Q_data_add_7_buff [1]), .CI(
        \u_decoder/fir_filter/add_332/carry [1]), .CO(
        \u_decoder/fir_filter/add_332/carry [2]), .S(
        \u_decoder/fir_filter/Q_data_add_6 [1]) );
  ADD32 \u_decoder/fir_filter/add_332/U1_2  ( .A(
        \u_decoder/fir_filter/Q_data_mult_6_buff [2]), .B(
        \u_decoder/fir_filter/Q_data_add_7_buff [2]), .CI(
        \u_decoder/fir_filter/add_332/carry [2]), .CO(
        \u_decoder/fir_filter/add_332/carry [3]), .S(
        \u_decoder/fir_filter/Q_data_add_6 [2]) );
  ADD32 \u_decoder/fir_filter/add_332/U1_3  ( .A(
        \u_decoder/fir_filter/Q_data_mult_6_buff [3]), .B(
        \u_decoder/fir_filter/Q_data_add_7_buff [3]), .CI(
        \u_decoder/fir_filter/add_332/carry [3]), .CO(
        \u_decoder/fir_filter/add_332/carry [4]), .S(
        \u_decoder/fir_filter/Q_data_add_6 [3]) );
  ADD32 \u_decoder/fir_filter/add_332/U1_4  ( .A(
        \u_decoder/fir_filter/Q_data_mult_6_buff [4]), .B(
        \u_decoder/fir_filter/Q_data_add_7_buff [4]), .CI(
        \u_decoder/fir_filter/add_332/carry [4]), .CO(
        \u_decoder/fir_filter/add_332/carry [5]), .S(
        \u_decoder/fir_filter/Q_data_add_6 [4]) );
  ADD32 \u_decoder/fir_filter/add_332/U1_5  ( .A(
        \u_decoder/fir_filter/Q_data_mult_6_buff [5]), .B(
        \u_decoder/fir_filter/Q_data_add_7_buff [5]), .CI(
        \u_decoder/fir_filter/add_332/carry [5]), .CO(
        \u_decoder/fir_filter/add_332/carry [6]), .S(
        \u_decoder/fir_filter/Q_data_add_6 [5]) );
  ADD32 \u_decoder/fir_filter/add_332/U1_6  ( .A(
        \u_decoder/fir_filter/Q_data_mult_6_buff [6]), .B(
        \u_decoder/fir_filter/Q_data_add_7_buff [6]), .CI(
        \u_decoder/fir_filter/add_332/carry [6]), .CO(
        \u_decoder/fir_filter/add_332/carry [7]), .S(
        \u_decoder/fir_filter/Q_data_add_6 [6]) );
  ADD32 \u_decoder/fir_filter/add_332/U1_7  ( .A(
        \u_decoder/fir_filter/Q_data_mult_6_buff [7]), .B(
        \u_decoder/fir_filter/Q_data_add_7_buff [7]), .CI(
        \u_decoder/fir_filter/add_332/carry [7]), .CO(
        \u_decoder/fir_filter/add_332/carry [8]), .S(
        \u_decoder/fir_filter/Q_data_add_6 [7]) );
  ADD32 \u_decoder/fir_filter/add_332/U1_8  ( .A(
        \u_decoder/fir_filter/Q_data_mult_6_buff [8]), .B(
        \u_decoder/fir_filter/Q_data_add_7_buff [8]), .CI(
        \u_decoder/fir_filter/add_332/carry [8]), .CO(
        \u_decoder/fir_filter/add_332/carry [9]), .S(
        \u_decoder/fir_filter/Q_data_add_6 [8]) );
  ADD32 \u_decoder/fir_filter/add_332/U1_9  ( .A(
        \u_decoder/fir_filter/Q_data_mult_6_buff [9]), .B(
        \u_decoder/fir_filter/Q_data_add_7_buff [9]), .CI(
        \u_decoder/fir_filter/add_332/carry [9]), .CO(
        \u_decoder/fir_filter/add_332/carry [10]), .S(
        \u_decoder/fir_filter/Q_data_add_6 [9]) );
  ADD32 \u_decoder/fir_filter/add_332/U1_10  ( .A(
        \u_decoder/fir_filter/Q_data_mult_6_buff [10]), .B(
        \u_decoder/fir_filter/Q_data_add_7_buff [10]), .CI(
        \u_decoder/fir_filter/add_332/carry [10]), .CO(
        \u_decoder/fir_filter/add_332/carry [11]), .S(
        \u_decoder/fir_filter/Q_data_add_6 [10]) );
  ADD32 \u_decoder/fir_filter/add_332/U1_11  ( .A(
        \u_decoder/fir_filter/Q_data_mult_6_buff [11]), .B(
        \u_decoder/fir_filter/Q_data_add_7_buff [11]), .CI(
        \u_decoder/fir_filter/add_332/carry [11]), .CO(
        \u_decoder/fir_filter/add_332/carry [12]), .S(
        \u_decoder/fir_filter/Q_data_add_6 [11]) );
  ADD32 \u_decoder/fir_filter/add_332/U1_12  ( .A(
        \u_decoder/fir_filter/Q_data_mult_6_buff [12]), .B(
        \u_decoder/fir_filter/Q_data_add_7_buff [12]), .CI(
        \u_decoder/fir_filter/add_332/carry [12]), .CO(
        \u_decoder/fir_filter/add_332/carry [13]), .S(
        \u_decoder/fir_filter/Q_data_add_6 [12]) );
  ADD32 \u_decoder/fir_filter/add_332/U1_13  ( .A(
        \u_decoder/fir_filter/Q_data_mult_6_buff [13]), .B(
        \u_decoder/fir_filter/Q_data_add_7_buff [13]), .CI(
        \u_decoder/fir_filter/add_332/carry [13]), .CO(
        \u_decoder/fir_filter/add_332/carry [14]), .S(
        \u_decoder/fir_filter/Q_data_add_6 [13]) );
  ADD32 \u_decoder/fir_filter/add_333/U1_1  ( .A(
        \u_decoder/fir_filter/Q_data_mult_7_buff [1]), .B(
        \u_decoder/fir_filter/Q_data_mult_8_buff [1]), .CI(
        \u_decoder/fir_filter/add_333/carry [1]), .CO(
        \u_decoder/fir_filter/add_333/carry [2]), .S(
        \u_decoder/fir_filter/Q_data_add_7 [1]) );
  ADD32 \u_decoder/fir_filter/add_333/U1_2  ( .A(
        \u_decoder/fir_filter/Q_data_mult_7_buff [2]), .B(
        \u_decoder/fir_filter/Q_data_mult_8_buff [2]), .CI(
        \u_decoder/fir_filter/add_333/carry [2]), .CO(
        \u_decoder/fir_filter/add_333/carry [3]), .S(
        \u_decoder/fir_filter/Q_data_add_7 [2]) );
  ADD32 \u_decoder/fir_filter/add_333/U1_3  ( .A(
        \u_decoder/fir_filter/Q_data_mult_7_buff [3]), .B(
        \u_decoder/fir_filter/Q_data_mult_8_buff [3]), .CI(
        \u_decoder/fir_filter/add_333/carry [3]), .CO(
        \u_decoder/fir_filter/add_333/carry [4]), .S(
        \u_decoder/fir_filter/Q_data_add_7 [3]) );
  ADD32 \u_decoder/fir_filter/add_333/U1_4  ( .A(
        \u_decoder/fir_filter/Q_data_mult_7_buff [4]), .B(
        \u_decoder/fir_filter/Q_data_mult_8_buff [4]), .CI(
        \u_decoder/fir_filter/add_333/carry [4]), .CO(
        \u_decoder/fir_filter/add_333/carry [5]), .S(
        \u_decoder/fir_filter/Q_data_add_7 [4]) );
  ADD32 \u_decoder/fir_filter/add_333/U1_5  ( .A(
        \u_decoder/fir_filter/Q_data_mult_7_buff [5]), .B(
        \u_decoder/fir_filter/Q_data_mult_8_buff [5]), .CI(
        \u_decoder/fir_filter/add_333/carry [5]), .CO(
        \u_decoder/fir_filter/add_333/carry [6]), .S(
        \u_decoder/fir_filter/Q_data_add_7 [5]) );
  ADD32 \u_decoder/fir_filter/add_333/U1_6  ( .A(
        \u_decoder/fir_filter/Q_data_mult_7_buff [6]), .B(
        \u_decoder/fir_filter/Q_data_mult_8_buff [6]), .CI(
        \u_decoder/fir_filter/add_333/carry [6]), .CO(
        \u_decoder/fir_filter/add_333/carry [7]), .S(
        \u_decoder/fir_filter/Q_data_add_7 [6]) );
  ADD32 \u_decoder/fir_filter/add_333/U1_7  ( .A(
        \u_decoder/fir_filter/Q_data_mult_7_buff [7]), .B(
        \u_decoder/fir_filter/Q_data_mult_8_buff [7]), .CI(
        \u_decoder/fir_filter/add_333/carry [7]), .CO(
        \u_decoder/fir_filter/add_333/carry [8]), .S(
        \u_decoder/fir_filter/Q_data_add_7 [7]) );
  ADD32 \u_decoder/fir_filter/add_333/U1_8  ( .A(
        \u_decoder/fir_filter/Q_data_mult_7_buff [8]), .B(
        \u_decoder/fir_filter/Q_data_mult_8_buff [8]), .CI(
        \u_decoder/fir_filter/add_333/carry [8]), .CO(
        \u_decoder/fir_filter/add_333/carry [9]), .S(
        \u_decoder/fir_filter/Q_data_add_7 [8]) );
  ADD32 \u_decoder/fir_filter/add_333/U1_9  ( .A(
        \u_decoder/fir_filter/Q_data_mult_7_buff [9]), .B(
        \u_decoder/fir_filter/Q_data_mult_8_buff [9]), .CI(
        \u_decoder/fir_filter/add_333/carry [9]), .CO(
        \u_decoder/fir_filter/add_333/carry [10]), .S(
        \u_decoder/fir_filter/Q_data_add_7 [9]) );
  ADD32 \u_decoder/fir_filter/add_333/U1_10  ( .A(
        \u_decoder/fir_filter/Q_data_mult_7_buff [10]), .B(
        \u_decoder/fir_filter/Q_data_mult_8_buff [10]), .CI(
        \u_decoder/fir_filter/add_333/carry [10]), .CO(
        \u_decoder/fir_filter/add_333/carry [11]), .S(
        \u_decoder/fir_filter/Q_data_add_7 [10]) );
  ADD32 \u_decoder/fir_filter/add_333/U1_11  ( .A(
        \u_decoder/fir_filter/Q_data_mult_7_buff [11]), .B(
        \u_decoder/fir_filter/Q_data_mult_8_buff [11]), .CI(
        \u_decoder/fir_filter/add_333/carry [11]), .CO(
        \u_decoder/fir_filter/add_333/carry [12]), .S(
        \u_decoder/fir_filter/Q_data_add_7 [11]) );
  ADD32 \u_decoder/fir_filter/add_333/U1_12  ( .A(
        \u_decoder/fir_filter/Q_data_mult_7_buff [12]), .B(
        \u_decoder/fir_filter/Q_data_mult_8_buff [12]), .CI(
        \u_decoder/fir_filter/add_333/carry [12]), .CO(
        \u_decoder/fir_filter/add_333/carry [13]), .S(
        \u_decoder/fir_filter/Q_data_add_7 [12]) );
  ADD32 \u_decoder/fir_filter/add_333/U1_13  ( .A(
        \u_decoder/fir_filter/Q_data_mult_7_buff [13]), .B(
        \u_decoder/fir_filter/Q_data_mult_8_buff [13]), .CI(
        \u_decoder/fir_filter/add_333/carry [13]), .CO(
        \u_decoder/fir_filter/add_333/carry [14]), .S(
        \u_decoder/fir_filter/Q_data_add_7 [13]) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/mult_276/S2_2_5  ( .A(n4), .B(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[1][5] ), .CI(n12), 
        .CO(\u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[2][5] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/SUMB[2][5] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/mult_276/S2_3_5  ( .A(n8), .B(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[2][5] ), .CI(n4), 
        .CO(\u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[3][5] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/SUMB[3][5] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/mult_276/S2_3_3  ( .A(n8), .B(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[2][3] ), .CI(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/SUMB[1][5] ), .CO(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[3][3] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/SUMB[3][3] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/mult_276/S2_4_5  ( .A(
        \u_decoder/I_prefilter [4]), .B(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[3][5] ), .CI(n8), 
        .CO(\u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[4][5] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/SUMB[4][5] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/mult_276/S2_4_3  ( .A(
        \u_decoder/I_prefilter [4]), .B(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[3][3] ), .CI(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/SUMB[2][5] ), .CO(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[4][3] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/SUMB[4][3] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/mult_276/S1_4_0  ( .A(
        \u_decoder/I_prefilter [4]), .B(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[3][0] ), .CI(n12), 
        .CO(\u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[4][0] ), .S(
        \u_decoder/fir_filter/I_data_mult_4 [4]) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/mult_276/S2_5_5  ( .A(n10), .B(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[4][5] ), .CI(
        \u_decoder/I_prefilter [4]), .CO(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[5][5] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/SUMB[5][5] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/mult_276/S2_5_3  ( .A(n10), .B(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[4][3] ), .CI(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/SUMB[3][5] ), .CO(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[5][3] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/SUMB[5][3] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/mult_276/S1_5_0  ( .A(n10), .B(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[4][0] ), .CI(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/SUMB[2][3] ), .CO(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[5][0] ), .S(
        \u_decoder/fir_filter/I_data_mult_4 [5]) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/mult_276/S2_6_5  ( .A(n6), .B(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[5][5] ), .CI(n10), 
        .CO(\u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[6][5] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/SUMB[6][5] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/mult_276/S2_6_3  ( .A(n6), .B(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[5][3] ), .CI(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/SUMB[4][5] ), .CO(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[6][3] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/SUMB[6][3] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/mult_276/S1_6_0  ( .A(n6), .B(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[5][0] ), .CI(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/SUMB[3][3] ), .CO(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[6][0] ), .S(
        \u_decoder/fir_filter/I_data_mult_4 [6]) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r167/S1_2_0  ( .A(n4), .B(
        \u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[1][0] ), .CI(n12), .CO(
        \u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[2][0] ), .S(
        \u_decoder/fir_filter/I_data_mult_3 [2]) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r167/S2_3_1  ( .A(n8), .B(
        \u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[2][1] ), .CI(n12), .CO(
        \u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[3][1] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/r167/SUMB[3][1] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r167/S1_3_0  ( .A(n8), .B(
        \u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[2][0] ), .CI(
        \u_decoder/fir_filter/dp_cluster_0/r167/SUMB[2][1] ), .CO(
        \u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[3][0] ), .S(
        \u_decoder/fir_filter/I_data_mult_3 [3]) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r167/S2_4_3  ( .A(
        \u_decoder/I_prefilter [4]), .B(
        \u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[3][3] ), .CI(n12), .CO(
        \u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[4][3] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/r167/SUMB[4][3] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r167/S2_4_1  ( .A(
        \u_decoder/I_prefilter [4]), .B(
        \u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[3][1] ), .CI(n4), .CO(
        \u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[4][1] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/r167/SUMB[4][1] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r167/S1_4_0  ( .A(
        \u_decoder/I_prefilter [4]), .B(
        \u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[3][0] ), .CI(
        \u_decoder/fir_filter/dp_cluster_0/r167/SUMB[3][1] ), .CO(
        \u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[4][0] ), .S(
        \u_decoder/fir_filter/I_data_mult_3 [4]) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r167/S2_5_3  ( .A(n10), .B(
        \u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[4][3] ), .CI(n4), .CO(
        \u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[5][3] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/r167/SUMB[5][3] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r167/S2_5_1  ( .A(n10), .B(
        \u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[4][1] ), .CI(
        \u_decoder/fir_filter/dp_cluster_0/r167/SUMB[3][3] ), .CO(
        \u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[5][1] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/r167/SUMB[5][1] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r167/S1_5_0  ( .A(n10), .B(
        \u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[4][0] ), .CI(
        \u_decoder/fir_filter/dp_cluster_0/r167/SUMB[4][1] ), .CO(
        \u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[5][0] ), .S(
        \u_decoder/fir_filter/I_data_mult_3 [5]) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r167/S2_6_3  ( .A(n6), .B(
        \u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[5][3] ), .CI(n8), .CO(
        \u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[6][3] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/r167/SUMB[6][3] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r167/S2_6_1  ( .A(n6), .B(
        \u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[5][1] ), .CI(
        \u_decoder/fir_filter/dp_cluster_0/r167/SUMB[4][3] ), .CO(
        \u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[6][1] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/r167/SUMB[6][1] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r167/S1_6_0  ( .A(n6), .B(
        \u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[5][0] ), .CI(
        \u_decoder/fir_filter/dp_cluster_0/r167/SUMB[5][1] ), .CO(
        \u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[6][0] ), .S(
        \u_decoder/fir_filter/I_data_mult_3 [6]) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r166/S2_2_3  ( .A(n4), .B(
        \u_decoder/fir_filter/dp_cluster_0/r166/CARRYB[1][3] ), .CI(n12), .CO(
        \u_decoder/fir_filter/dp_cluster_0/r166/CARRYB[2][3] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/r166/SUMB[2][3] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r166/S2_3_3  ( .A(n8), .B(
        \u_decoder/fir_filter/dp_cluster_0/r166/CARRYB[2][3] ), .CI(n4), .CO(
        \u_decoder/fir_filter/dp_cluster_0/r166/CARRYB[3][3] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/r166/SUMB[3][3] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r166/S2_3_1  ( .A(n8), .B(
        \u_decoder/fir_filter/dp_cluster_0/r166/CARRYB[2][1] ), .CI(
        \u_decoder/fir_filter/dp_cluster_0/r166/SUMB[1][3] ), .CO(
        \u_decoder/fir_filter/dp_cluster_0/r166/CARRYB[3][1] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/r166/SUMB[3][1] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r166/S2_4_3  ( .A(
        \u_decoder/I_prefilter [4]), .B(
        \u_decoder/fir_filter/dp_cluster_0/r166/CARRYB[3][3] ), .CI(n8), .CO(
        \u_decoder/fir_filter/dp_cluster_0/r166/CARRYB[4][3] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/r166/SUMB[4][3] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r166/S2_4_1  ( .A(
        \u_decoder/I_prefilter [4]), .B(
        \u_decoder/fir_filter/dp_cluster_0/r166/CARRYB[3][1] ), .CI(
        \u_decoder/fir_filter/dp_cluster_0/r166/SUMB[2][3] ), .CO(
        \u_decoder/fir_filter/dp_cluster_0/r166/CARRYB[4][1] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/r166/SUMB[4][1] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r166/S2_5_3  ( .A(n10), .B(
        \u_decoder/fir_filter/dp_cluster_0/r166/CARRYB[4][3] ), .CI(
        \u_decoder/I_prefilter [4]), .CO(
        \u_decoder/fir_filter/dp_cluster_0/r166/CARRYB[5][3] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/r166/SUMB[5][3] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r166/S2_5_1  ( .A(n10), .B(
        \u_decoder/fir_filter/dp_cluster_0/r166/CARRYB[4][1] ), .CI(
        \u_decoder/fir_filter/dp_cluster_0/r166/SUMB[3][3] ), .CO(
        \u_decoder/fir_filter/dp_cluster_0/r166/CARRYB[5][1] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/r166/SUMB[5][1] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r166/S2_6_3  ( .A(n6), .B(
        \u_decoder/fir_filter/dp_cluster_0/r166/CARRYB[5][3] ), .CI(n10), .CO(
        \u_decoder/fir_filter/dp_cluster_0/r166/CARRYB[6][3] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/r166/SUMB[6][3] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r166/S2_6_1  ( .A(n6), .B(
        \u_decoder/fir_filter/dp_cluster_0/r166/CARRYB[5][1] ), .CI(
        \u_decoder/fir_filter/dp_cluster_0/r166/SUMB[4][3] ), .CO(
        \u_decoder/fir_filter/dp_cluster_0/r166/CARRYB[6][1] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/r166/SUMB[6][1] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r165/S2_3_3  ( .A(n8), .B(
        \u_decoder/fir_filter/dp_cluster_0/r165/CARRYB[2][3] ), .CI(n74), .CO(
        \u_decoder/fir_filter/dp_cluster_0/r165/CARRYB[3][3] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/r165/SUMB[3][3] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r165/S2_4_3  ( .A(
        \u_decoder/I_prefilter [4]), .B(
        \u_decoder/fir_filter/dp_cluster_0/r165/CARRYB[3][3] ), .CI(n89), .CO(
        \u_decoder/fir_filter/dp_cluster_0/r165/CARRYB[4][3] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/r165/SUMB[4][3] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r165/S1_4_0  ( .A(
        \u_decoder/I_prefilter [4]), .B(
        \u_decoder/fir_filter/dp_cluster_0/r165/CARRYB[3][0] ), .CI(n12), .CO(
        \u_decoder/fir_filter/dp_cluster_0/r165/CARRYB[4][0] ), .S(
        \u_decoder/fir_filter/I_data_mult_1[4] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r165/S2_5_3  ( .A(n10), .B(
        \u_decoder/fir_filter/dp_cluster_0/r165/CARRYB[4][3] ), .CI(n80), .CO(
        \u_decoder/fir_filter/dp_cluster_0/r165/CARRYB[5][3] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/r165/SUMB[5][3] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r165/S1_5_0  ( .A(n10), .B(
        \u_decoder/fir_filter/dp_cluster_0/r165/CARRYB[4][0] ), .CI(
        \u_decoder/fir_filter/dp_cluster_0/r165/SUMB[2][3] ), .CO(
        \u_decoder/fir_filter/dp_cluster_0/r165/CARRYB[5][0] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/r165/PROD1[5] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r165/S2_6_3  ( .A(n6), .B(
        \u_decoder/fir_filter/dp_cluster_0/r165/CARRYB[5][3] ), .CI(n164), 
        .CO(\u_decoder/fir_filter/dp_cluster_0/r165/CARRYB[6][3] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/r165/SUMB[6][3] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r165/S1_6_0  ( .A(n6), .B(
        \u_decoder/fir_filter/dp_cluster_0/r165/CARRYB[5][0] ), .CI(
        \u_decoder/fir_filter/dp_cluster_0/r165/SUMB[3][3] ), .CO(
        \u_decoder/fir_filter/dp_cluster_0/r165/CARRYB[6][0] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/r165/A1[4] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r164/S2_3_2  ( .A(n8), .B(
        \u_decoder/fir_filter/dp_cluster_0/r164/CARRYB[2][2] ), .CI(n74), .CO(
        \u_decoder/fir_filter/dp_cluster_0/r164/CARRYB[3][2] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/r164/SUMB[3][2] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r164/S1_3_0  ( .A(n8), .B(
        \u_decoder/fir_filter/dp_cluster_0/r164/CARRYB[2][0] ), .CI(n12), .CO(
        \u_decoder/fir_filter/dp_cluster_0/r164/CARRYB[3][0] ), .S(
        \u_decoder/fir_filter/I_data_mult_0 [3]) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r164/S2_4_2  ( .A(
        \u_decoder/I_prefilter [4]), .B(
        \u_decoder/fir_filter/dp_cluster_0/r164/CARRYB[3][2] ), .CI(n89), .CO(
        \u_decoder/fir_filter/dp_cluster_0/r164/CARRYB[4][2] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/r164/SUMB[4][2] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r164/S1_4_0  ( .A(
        \u_decoder/I_prefilter [4]), .B(
        \u_decoder/fir_filter/dp_cluster_0/r164/CARRYB[3][0] ), .CI(
        \u_decoder/fir_filter/dp_cluster_0/r164/SUMB[2][2] ), .CO(
        \u_decoder/fir_filter/dp_cluster_0/r164/CARRYB[4][0] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/r164/PROD1[4] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r164/S2_5_2  ( .A(n10), .B(
        \u_decoder/fir_filter/dp_cluster_0/r164/CARRYB[4][2] ), .CI(n80), .CO(
        \u_decoder/fir_filter/dp_cluster_0/r164/CARRYB[5][2] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/r164/SUMB[5][2] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r164/S1_5_0  ( .A(n10), .B(
        \u_decoder/fir_filter/dp_cluster_0/r164/CARRYB[4][0] ), .CI(
        \u_decoder/fir_filter/dp_cluster_0/r164/SUMB[3][2] ), .CO(
        \u_decoder/fir_filter/dp_cluster_0/r164/CARRYB[5][0] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/r164/A1[3] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r164/S2_6_2  ( .A(n6), .B(
        \u_decoder/fir_filter/dp_cluster_0/r164/CARRYB[5][2] ), .CI(n164), 
        .CO(\u_decoder/fir_filter/dp_cluster_0/r164/CARRYB[6][2] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/r164/SUMB[6][2] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r164/S1_6_0  ( .A(n6), .B(
        \u_decoder/fir_filter/dp_cluster_0/r164/CARRYB[5][0] ), .CI(
        \u_decoder/fir_filter/dp_cluster_0/r164/SUMB[4][2] ), .CO(
        \u_decoder/fir_filter/dp_cluster_0/r164/CARRYB[6][0] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/r164/A1[4] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/mult_308/S2_2_5  ( .A(n3), .B(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[1][5] ), .CI(n11), 
        .CO(\u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[2][5] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/SUMB[2][5] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/mult_308/S2_3_5  ( .A(n7), .B(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[2][5] ), .CI(n3), 
        .CO(\u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[3][5] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/SUMB[3][5] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/mult_308/S2_3_3  ( .A(n7), .B(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[2][3] ), .CI(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/SUMB[1][5] ), .CO(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[3][3] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/SUMB[3][3] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/mult_308/S2_4_5  ( .A(
        \u_decoder/Q_prefilter [4]), .B(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[3][5] ), .CI(n7), 
        .CO(\u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[4][5] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/SUMB[4][5] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/mult_308/S2_4_3  ( .A(
        \u_decoder/Q_prefilter [4]), .B(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[3][3] ), .CI(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/SUMB[2][5] ), .CO(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[4][3] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/SUMB[4][3] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/mult_308/S1_4_0  ( .A(
        \u_decoder/Q_prefilter [4]), .B(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[3][0] ), .CI(n11), 
        .CO(\u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[4][0] ), .S(
        \u_decoder/fir_filter/Q_data_mult_4 [4]) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/mult_308/S2_5_5  ( .A(n9), .B(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[4][5] ), .CI(
        \u_decoder/Q_prefilter [4]), .CO(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[5][5] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/SUMB[5][5] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/mult_308/S2_5_3  ( .A(n9), .B(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[4][3] ), .CI(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/SUMB[3][5] ), .CO(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[5][3] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/SUMB[5][3] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/mult_308/S1_5_0  ( .A(n9), .B(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[4][0] ), .CI(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/SUMB[2][3] ), .CO(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[5][0] ), .S(
        \u_decoder/fir_filter/Q_data_mult_4 [5]) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/mult_308/S2_6_5  ( .A(n5), .B(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[5][5] ), .CI(n9), 
        .CO(\u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[6][5] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/SUMB[6][5] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/mult_308/S2_6_3  ( .A(n5), .B(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[5][3] ), .CI(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/SUMB[4][5] ), .CO(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[6][3] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/SUMB[6][3] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/mult_308/S1_6_0  ( .A(n5), .B(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[5][0] ), .CI(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/SUMB[3][3] ), .CO(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[6][0] ), .S(
        \u_decoder/fir_filter/Q_data_mult_4 [6]) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r180/S1_2_0  ( .A(n3), .B(
        \u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[1][0] ), .CI(n11), .CO(
        \u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[2][0] ), .S(
        \u_decoder/fir_filter/Q_data_mult_3 [2]) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r180/S2_3_1  ( .A(n7), .B(
        \u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[2][1] ), .CI(n11), .CO(
        \u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[3][1] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/r180/SUMB[3][1] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r180/S1_3_0  ( .A(n7), .B(
        \u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[2][0] ), .CI(
        \u_decoder/fir_filter/dp_cluster_0/r180/SUMB[2][1] ), .CO(
        \u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[3][0] ), .S(
        \u_decoder/fir_filter/Q_data_mult_3 [3]) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r180/S2_4_3  ( .A(
        \u_decoder/Q_prefilter [4]), .B(
        \u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[3][3] ), .CI(n11), .CO(
        \u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[4][3] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/r180/SUMB[4][3] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r180/S2_4_1  ( .A(
        \u_decoder/Q_prefilter [4]), .B(
        \u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[3][1] ), .CI(n3), .CO(
        \u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[4][1] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/r180/SUMB[4][1] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r180/S1_4_0  ( .A(
        \u_decoder/Q_prefilter [4]), .B(
        \u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[3][0] ), .CI(
        \u_decoder/fir_filter/dp_cluster_0/r180/SUMB[3][1] ), .CO(
        \u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[4][0] ), .S(
        \u_decoder/fir_filter/Q_data_mult_3 [4]) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r180/S2_5_3  ( .A(n9), .B(
        \u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[4][3] ), .CI(n3), .CO(
        \u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[5][3] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/r180/SUMB[5][3] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r180/S2_5_1  ( .A(n9), .B(
        \u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[4][1] ), .CI(
        \u_decoder/fir_filter/dp_cluster_0/r180/SUMB[3][3] ), .CO(
        \u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[5][1] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/r180/SUMB[5][1] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r180/S1_5_0  ( .A(n9), .B(
        \u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[4][0] ), .CI(
        \u_decoder/fir_filter/dp_cluster_0/r180/SUMB[4][1] ), .CO(
        \u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[5][0] ), .S(
        \u_decoder/fir_filter/Q_data_mult_3 [5]) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r180/S2_6_3  ( .A(n5), .B(
        \u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[5][3] ), .CI(n7), .CO(
        \u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[6][3] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/r180/SUMB[6][3] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r180/S2_6_1  ( .A(n5), .B(
        \u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[5][1] ), .CI(
        \u_decoder/fir_filter/dp_cluster_0/r180/SUMB[4][3] ), .CO(
        \u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[6][1] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/r180/SUMB[6][1] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r180/S1_6_0  ( .A(n5), .B(
        \u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[5][0] ), .CI(
        \u_decoder/fir_filter/dp_cluster_0/r180/SUMB[5][1] ), .CO(
        \u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[6][0] ), .S(
        \u_decoder/fir_filter/Q_data_mult_3 [6]) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r179/S2_2_3  ( .A(n3), .B(
        \u_decoder/fir_filter/dp_cluster_0/r179/CARRYB[1][3] ), .CI(n11), .CO(
        \u_decoder/fir_filter/dp_cluster_0/r179/CARRYB[2][3] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/r179/SUMB[2][3] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r179/S2_3_3  ( .A(n7), .B(
        \u_decoder/fir_filter/dp_cluster_0/r179/CARRYB[2][3] ), .CI(n3), .CO(
        \u_decoder/fir_filter/dp_cluster_0/r179/CARRYB[3][3] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/r179/SUMB[3][3] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r179/S2_3_1  ( .A(n7), .B(
        \u_decoder/fir_filter/dp_cluster_0/r179/CARRYB[2][1] ), .CI(
        \u_decoder/fir_filter/dp_cluster_0/r179/SUMB[1][3] ), .CO(
        \u_decoder/fir_filter/dp_cluster_0/r179/CARRYB[3][1] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/r179/SUMB[3][1] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r179/S2_4_3  ( .A(
        \u_decoder/Q_prefilter [4]), .B(
        \u_decoder/fir_filter/dp_cluster_0/r179/CARRYB[3][3] ), .CI(n7), .CO(
        \u_decoder/fir_filter/dp_cluster_0/r179/CARRYB[4][3] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/r179/SUMB[4][3] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r179/S2_4_1  ( .A(
        \u_decoder/Q_prefilter [4]), .B(
        \u_decoder/fir_filter/dp_cluster_0/r179/CARRYB[3][1] ), .CI(
        \u_decoder/fir_filter/dp_cluster_0/r179/SUMB[2][3] ), .CO(
        \u_decoder/fir_filter/dp_cluster_0/r179/CARRYB[4][1] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/r179/SUMB[4][1] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r179/S2_5_3  ( .A(n9), .B(
        \u_decoder/fir_filter/dp_cluster_0/r179/CARRYB[4][3] ), .CI(
        \u_decoder/Q_prefilter [4]), .CO(
        \u_decoder/fir_filter/dp_cluster_0/r179/CARRYB[5][3] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/r179/SUMB[5][3] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r179/S2_5_1  ( .A(n9), .B(
        \u_decoder/fir_filter/dp_cluster_0/r179/CARRYB[4][1] ), .CI(
        \u_decoder/fir_filter/dp_cluster_0/r179/SUMB[3][3] ), .CO(
        \u_decoder/fir_filter/dp_cluster_0/r179/CARRYB[5][1] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/r179/SUMB[5][1] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r179/S2_6_3  ( .A(n5), .B(
        \u_decoder/fir_filter/dp_cluster_0/r179/CARRYB[5][3] ), .CI(n9), .CO(
        \u_decoder/fir_filter/dp_cluster_0/r179/CARRYB[6][3] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/r179/SUMB[6][3] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r179/S2_6_1  ( .A(n5), .B(
        \u_decoder/fir_filter/dp_cluster_0/r179/CARRYB[5][1] ), .CI(
        \u_decoder/fir_filter/dp_cluster_0/r179/SUMB[4][3] ), .CO(
        \u_decoder/fir_filter/dp_cluster_0/r179/CARRYB[6][1] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/r179/SUMB[6][1] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r178/S2_3_3  ( .A(n7), .B(
        \u_decoder/fir_filter/dp_cluster_0/r178/CARRYB[2][3] ), .CI(n75), .CO(
        \u_decoder/fir_filter/dp_cluster_0/r178/CARRYB[3][3] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/r178/SUMB[3][3] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r178/S2_4_3  ( .A(
        \u_decoder/Q_prefilter [4]), .B(
        \u_decoder/fir_filter/dp_cluster_0/r178/CARRYB[3][3] ), .CI(n90), .CO(
        \u_decoder/fir_filter/dp_cluster_0/r178/CARRYB[4][3] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/r178/SUMB[4][3] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r178/S1_4_0  ( .A(
        \u_decoder/Q_prefilter [4]), .B(
        \u_decoder/fir_filter/dp_cluster_0/r178/CARRYB[3][0] ), .CI(n11), .CO(
        \u_decoder/fir_filter/dp_cluster_0/r178/CARRYB[4][0] ), .S(
        \u_decoder/fir_filter/Q_data_mult_1[4] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r178/S2_5_3  ( .A(n9), .B(
        \u_decoder/fir_filter/dp_cluster_0/r178/CARRYB[4][3] ), .CI(n81), .CO(
        \u_decoder/fir_filter/dp_cluster_0/r178/CARRYB[5][3] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/r178/SUMB[5][3] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r178/S1_5_0  ( .A(n9), .B(
        \u_decoder/fir_filter/dp_cluster_0/r178/CARRYB[4][0] ), .CI(
        \u_decoder/fir_filter/dp_cluster_0/r178/SUMB[2][3] ), .CO(
        \u_decoder/fir_filter/dp_cluster_0/r178/CARRYB[5][0] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/r178/PROD1[5] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r178/S2_6_3  ( .A(n5), .B(
        \u_decoder/fir_filter/dp_cluster_0/r178/CARRYB[5][3] ), .CI(n165), 
        .CO(\u_decoder/fir_filter/dp_cluster_0/r178/CARRYB[6][3] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/r178/SUMB[6][3] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r178/S1_6_0  ( .A(n5), .B(
        \u_decoder/fir_filter/dp_cluster_0/r178/CARRYB[5][0] ), .CI(
        \u_decoder/fir_filter/dp_cluster_0/r178/SUMB[3][3] ), .CO(
        \u_decoder/fir_filter/dp_cluster_0/r178/CARRYB[6][0] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/r178/A1[4] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r177/S2_3_2  ( .A(n7), .B(
        \u_decoder/fir_filter/dp_cluster_0/r177/CARRYB[2][2] ), .CI(n75), .CO(
        \u_decoder/fir_filter/dp_cluster_0/r177/CARRYB[3][2] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/r177/SUMB[3][2] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r177/S1_3_0  ( .A(n7), .B(
        \u_decoder/fir_filter/dp_cluster_0/r177/CARRYB[2][0] ), .CI(n11), .CO(
        \u_decoder/fir_filter/dp_cluster_0/r177/CARRYB[3][0] ), .S(
        \u_decoder/fir_filter/Q_data_mult_0 [3]) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r177/S2_4_2  ( .A(
        \u_decoder/Q_prefilter [4]), .B(
        \u_decoder/fir_filter/dp_cluster_0/r177/CARRYB[3][2] ), .CI(n90), .CO(
        \u_decoder/fir_filter/dp_cluster_0/r177/CARRYB[4][2] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/r177/SUMB[4][2] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r177/S1_4_0  ( .A(
        \u_decoder/Q_prefilter [4]), .B(
        \u_decoder/fir_filter/dp_cluster_0/r177/CARRYB[3][0] ), .CI(
        \u_decoder/fir_filter/dp_cluster_0/r177/SUMB[2][2] ), .CO(
        \u_decoder/fir_filter/dp_cluster_0/r177/CARRYB[4][0] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/r177/PROD1[4] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r177/S2_5_2  ( .A(n9), .B(
        \u_decoder/fir_filter/dp_cluster_0/r177/CARRYB[4][2] ), .CI(n81), .CO(
        \u_decoder/fir_filter/dp_cluster_0/r177/CARRYB[5][2] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/r177/SUMB[5][2] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r177/S1_5_0  ( .A(n9), .B(
        \u_decoder/fir_filter/dp_cluster_0/r177/CARRYB[4][0] ), .CI(
        \u_decoder/fir_filter/dp_cluster_0/r177/SUMB[3][2] ), .CO(
        \u_decoder/fir_filter/dp_cluster_0/r177/CARRYB[5][0] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/r177/A1[3] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r177/S2_6_2  ( .A(n5), .B(
        \u_decoder/fir_filter/dp_cluster_0/r177/CARRYB[5][2] ), .CI(n165), 
        .CO(\u_decoder/fir_filter/dp_cluster_0/r177/CARRYB[6][2] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/r177/SUMB[6][2] ) );
  ADD32 \u_decoder/fir_filter/dp_cluster_0/r177/S1_6_0  ( .A(n5), .B(
        \u_decoder/fir_filter/dp_cluster_0/r177/CARRYB[5][0] ), .CI(
        \u_decoder/fir_filter/dp_cluster_0/r177/SUMB[4][2] ), .CO(
        \u_decoder/fir_filter/dp_cluster_0/r177/CARRYB[6][0] ), .S(
        \u_decoder/fir_filter/dp_cluster_0/r177/A1[4] ) );
  ADD32 \u_decoder/iq_demod/dp_cluster_0/mult_151/S3_2_2  ( .A(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/ab[2][2] ), .B(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/CARRYB[1][2] ), .CI(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/ab[1][3] ), .CO(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/CARRYB[2][2] ), .S(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/SUMB[2][2] ) );
  ADD32 \u_decoder/iq_demod/dp_cluster_0/mult_151/S2_2_1  ( .A(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/ab[2][1] ), .B(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/CARRYB[1][1] ), .CI(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/SUMB[1][2] ), .CO(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/CARRYB[2][1] ), .S(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/SUMB[2][1] ) );
  ADD32 \u_decoder/iq_demod/dp_cluster_0/mult_151/S1_2_0  ( .A(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/ab[2][0] ), .B(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/CARRYB[1][0] ), .CI(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/SUMB[1][1] ), .CO(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/CARRYB[2][0] ), .S(
        \u_decoder/iq_demod/dp_cluster_0/mult_Q_sin_out [2]) );
  ADD32 \u_decoder/iq_demod/dp_cluster_0/mult_151/S14_3  ( .A(
        \u_decoder/iq_demod/Q_if_buff[3] ), .B(n23), .CI(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/ab[3][3] ), .CO(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/CARRYB[3][3] ), .S(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/SUMB[3][3] ) );
  ADD32 \u_decoder/iq_demod/dp_cluster_0/mult_151/S5_2  ( .A(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/ab[3][2] ), .B(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/CARRYB[2][2] ), .CI(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/ab[2][3] ), .CO(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/CARRYB[3][2] ), .S(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/SUMB[3][2] ) );
  ADD32 \u_decoder/iq_demod/dp_cluster_0/mult_151/S4_1  ( .A(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/ab[3][1] ), .B(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/CARRYB[2][1] ), .CI(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/SUMB[2][2] ), .CO(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/CARRYB[3][1] ), .S(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/SUMB[3][1] ) );
  ADD32 \u_decoder/iq_demod/dp_cluster_0/mult_151/S4_0  ( .A(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/ab[3][0] ), .B(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/CARRYB[2][0] ), .CI(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/SUMB[2][1] ), .CO(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/CARRYB[3][0] ), .S(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/SUMB[3][0] ) );
  ADD32 \u_decoder/iq_demod/dp_cluster_0/mult_151/S14_3_0  ( .A(
        \u_decoder/iq_demod/Q_if_signed [3]), .B(
        \u_decoder/iq_demod/sin_out [3]), .CI(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/SUMB[3][0] ), .CO(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/A2[2] ), .S(
        \u_decoder/iq_demod/dp_cluster_0/mult_Q_sin_out [3]) );
  ADD32 \u_decoder/iq_demod/dp_cluster_0/mult_148/S3_2_2  ( .A(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/ab[2][2] ), .B(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/CARRYB[1][2] ), .CI(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/ab[1][3] ), .CO(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/CARRYB[2][2] ), .S(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/SUMB[2][2] ) );
  ADD32 \u_decoder/iq_demod/dp_cluster_0/mult_148/S2_2_1  ( .A(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/ab[2][1] ), .B(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/CARRYB[1][1] ), .CI(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/SUMB[1][2] ), .CO(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/CARRYB[2][1] ), .S(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/SUMB[2][1] ) );
  ADD32 \u_decoder/iq_demod/dp_cluster_0/mult_148/S1_2_0  ( .A(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/ab[2][0] ), .B(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/CARRYB[1][0] ), .CI(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/SUMB[1][1] ), .CO(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/CARRYB[2][0] ), .S(
        \u_decoder/iq_demod/dp_cluster_0/mult_I_cos_out [2]) );
  ADD32 \u_decoder/iq_demod/dp_cluster_0/mult_148/S14_3  ( .A(
        \u_decoder/iq_demod/I_if_buff[3] ), .B(n22), .CI(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/ab[3][3] ), .CO(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/CARRYB[3][3] ), .S(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/SUMB[3][3] ) );
  ADD32 \u_decoder/iq_demod/dp_cluster_0/mult_148/S5_2  ( .A(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/ab[3][2] ), .B(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/CARRYB[2][2] ), .CI(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/ab[2][3] ), .CO(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/CARRYB[3][2] ), .S(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/SUMB[3][2] ) );
  ADD32 \u_decoder/iq_demod/dp_cluster_0/mult_148/S4_1  ( .A(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/ab[3][1] ), .B(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/CARRYB[2][1] ), .CI(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/SUMB[2][2] ), .CO(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/CARRYB[3][1] ), .S(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/SUMB[3][1] ) );
  ADD32 \u_decoder/iq_demod/dp_cluster_0/mult_148/S4_0  ( .A(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/ab[3][0] ), .B(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/CARRYB[2][0] ), .CI(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/SUMB[2][1] ), .CO(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/CARRYB[3][0] ), .S(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/SUMB[3][0] ) );
  ADD32 \u_decoder/iq_demod/dp_cluster_0/mult_148/S14_3_0  ( .A(
        \u_decoder/iq_demod/I_if_signed [3]), .B(
        \u_decoder/iq_demod/cos_out [3]), .CI(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/SUMB[3][0] ), .CO(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/A2[2] ), .S(
        \u_decoder/iq_demod/dp_cluster_0/mult_I_cos_out [3]) );
  ADD32 \u_decoder/iq_demod/dp_cluster_0/sub_153/U2_1  ( .A(
        \u_decoder/iq_demod/dp_cluster_0/mult_I_cos_out [1]), .B(n170), .CI(
        \u_decoder/iq_demod/dp_cluster_0/sub_153/carry [1]), .CO(
        \u_decoder/iq_demod/dp_cluster_0/sub_153/carry [2]), .S(
        \u_decoder/iq_demod/add_I_out [1]) );
  ADD32 \u_decoder/iq_demod/dp_cluster_0/sub_153/U2_2  ( .A(
        \u_decoder/iq_demod/dp_cluster_0/mult_I_cos_out [2]), .B(n2388), .CI(
        \u_decoder/iq_demod/dp_cluster_0/sub_153/carry [2]), .CO(
        \u_decoder/iq_demod/dp_cluster_0/sub_153/carry [3]), .S(
        \u_decoder/iq_demod/add_I_out [2]) );
  ADD32 \u_decoder/iq_demod/dp_cluster_0/sub_153/U2_3  ( .A(
        \u_decoder/iq_demod/dp_cluster_0/mult_I_cos_out [3]), .B(n2387), .CI(
        \u_decoder/iq_demod/dp_cluster_0/sub_153/carry [3]), .CO(
        \u_decoder/iq_demod/dp_cluster_0/sub_153/carry [4]), .S(
        \u_decoder/iq_demod/add_I_out [3]) );
  ADD32 \u_decoder/iq_demod/dp_cluster_0/sub_153/U2_4  ( .A(
        \u_decoder/iq_demod/dp_cluster_0/mult_I_cos_out [4]), .B(n83), .CI(
        \u_decoder/iq_demod/dp_cluster_0/sub_153/carry [4]), .CO(
        \u_decoder/iq_demod/dp_cluster_0/sub_153/carry [5]), .S(
        \u_decoder/iq_demod/add_I_out [4]) );
  ADD32 \u_decoder/iq_demod/dp_cluster_0/sub_153/U2_5  ( .A(
        \u_decoder/iq_demod/dp_cluster_0/mult_I_cos_out [5]), .B(n82), .CI(
        \u_decoder/iq_demod/dp_cluster_0/sub_153/carry [5]), .CO(
        \u_decoder/iq_demod/dp_cluster_0/sub_153/carry [6]), .S(
        \u_decoder/iq_demod/add_I_out [5]) );
  ADD32 \u_decoder/iq_demod/dp_cluster_0/sub_153/U2_6  ( .A(
        \u_decoder/iq_demod/dp_cluster_0/mult_I_cos_out [6]), .B(n349), .CI(
        \u_decoder/iq_demod/dp_cluster_0/sub_153/carry [6]), .CO(
        \u_decoder/iq_demod/dp_cluster_0/sub_153/carry [7]), .S(
        \u_decoder/iq_demod/add_I_out [6]) );
  ADD32 \u_decoder/iq_demod/dp_cluster_1/mult_150/S3_2_2  ( .A(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/ab[2][2] ), .B(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/CARRYB[1][2] ), .CI(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/ab[1][3] ), .CO(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/CARRYB[2][2] ), .S(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/SUMB[2][2] ) );
  ADD32 \u_decoder/iq_demod/dp_cluster_1/mult_150/S2_2_1  ( .A(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/ab[2][1] ), .B(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/CARRYB[1][1] ), .CI(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/SUMB[1][2] ), .CO(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/CARRYB[2][1] ), .S(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/SUMB[2][1] ) );
  ADD32 \u_decoder/iq_demod/dp_cluster_1/mult_150/S1_2_0  ( .A(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/ab[2][0] ), .B(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/CARRYB[1][0] ), .CI(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/SUMB[1][1] ), .CO(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/CARRYB[2][0] ), .S(
        \u_decoder/iq_demod/dp_cluster_1/mult_Q_cos_out [2]) );
  ADD32 \u_decoder/iq_demod/dp_cluster_1/mult_150/S14_3  ( .A(
        \u_decoder/iq_demod/Q_if_buff[3] ), .B(n22), .CI(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/ab[3][3] ), .CO(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/CARRYB[3][3] ), .S(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/SUMB[3][3] ) );
  ADD32 \u_decoder/iq_demod/dp_cluster_1/mult_150/S5_2  ( .A(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/ab[3][2] ), .B(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/CARRYB[2][2] ), .CI(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/ab[2][3] ), .CO(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/CARRYB[3][2] ), .S(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/SUMB[3][2] ) );
  ADD32 \u_decoder/iq_demod/dp_cluster_1/mult_150/S4_1  ( .A(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/ab[3][1] ), .B(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/CARRYB[2][1] ), .CI(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/SUMB[2][2] ), .CO(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/CARRYB[3][1] ), .S(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/SUMB[3][1] ) );
  ADD32 \u_decoder/iq_demod/dp_cluster_1/mult_150/S4_0  ( .A(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/ab[3][0] ), .B(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/CARRYB[2][0] ), .CI(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/SUMB[2][1] ), .CO(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/CARRYB[3][0] ), .S(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/SUMB[3][0] ) );
  ADD32 \u_decoder/iq_demod/dp_cluster_1/mult_150/S14_3_0  ( .A(
        \u_decoder/iq_demod/Q_if_signed [3]), .B(
        \u_decoder/iq_demod/cos_out [3]), .CI(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/SUMB[3][0] ), .CO(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/A2[2] ), .S(
        \u_decoder/iq_demod/dp_cluster_1/mult_Q_cos_out [3]) );
  ADD32 \u_decoder/iq_demod/dp_cluster_1/mult_149/S3_2_2  ( .A(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/ab[2][2] ), .B(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/CARRYB[1][2] ), .CI(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/ab[1][3] ), .CO(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/CARRYB[2][2] ), .S(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/SUMB[2][2] ) );
  ADD32 \u_decoder/iq_demod/dp_cluster_1/mult_149/S2_2_1  ( .A(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/ab[2][1] ), .B(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/CARRYB[1][1] ), .CI(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/SUMB[1][2] ), .CO(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/CARRYB[2][1] ), .S(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/SUMB[2][1] ) );
  ADD32 \u_decoder/iq_demod/dp_cluster_1/mult_149/S1_2_0  ( .A(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/ab[2][0] ), .B(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/CARRYB[1][0] ), .CI(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/SUMB[1][1] ), .CO(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/CARRYB[2][0] ), .S(
        \u_decoder/iq_demod/dp_cluster_1/mult_I_sin_out [2]) );
  ADD32 \u_decoder/iq_demod/dp_cluster_1/mult_149/S14_3  ( .A(
        \u_decoder/iq_demod/I_if_buff[3] ), .B(n23), .CI(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/ab[3][3] ), .CO(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/CARRYB[3][3] ), .S(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/SUMB[3][3] ) );
  ADD32 \u_decoder/iq_demod/dp_cluster_1/mult_149/S5_2  ( .A(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/ab[3][2] ), .B(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/CARRYB[2][2] ), .CI(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/ab[2][3] ), .CO(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/CARRYB[3][2] ), .S(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/SUMB[3][2] ) );
  ADD32 \u_decoder/iq_demod/dp_cluster_1/mult_149/S4_1  ( .A(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/ab[3][1] ), .B(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/CARRYB[2][1] ), .CI(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/SUMB[2][2] ), .CO(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/CARRYB[3][1] ), .S(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/SUMB[3][1] ) );
  ADD32 \u_decoder/iq_demod/dp_cluster_1/mult_149/S4_0  ( .A(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/ab[3][0] ), .B(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/CARRYB[2][0] ), .CI(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/SUMB[2][1] ), .CO(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/CARRYB[3][0] ), .S(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/SUMB[3][0] ) );
  ADD32 \u_decoder/iq_demod/dp_cluster_1/mult_149/S14_3_0  ( .A(
        \u_decoder/iq_demod/I_if_signed [3]), .B(
        \u_decoder/iq_demod/sin_out [3]), .CI(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/SUMB[3][0] ), .CO(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/A2[2] ), .S(
        \u_decoder/iq_demod/dp_cluster_1/mult_I_sin_out [3]) );
  ADD32 \u_decoder/iq_demod/dp_cluster_1/add_154/U1_1  ( .A(
        \u_decoder/iq_demod/dp_cluster_1/mult_I_sin_out [1]), .B(
        \u_decoder/iq_demod/dp_cluster_1/mult_Q_cos_out [1]), .CI(
        \u_decoder/iq_demod/dp_cluster_1/add_154/carry [1]), .CO(
        \u_decoder/iq_demod/dp_cluster_1/add_154/carry [2]), .S(
        \u_decoder/iq_demod/add_Q_out [1]) );
  ADD32 \u_decoder/iq_demod/dp_cluster_1/add_154/U1_2  ( .A(
        \u_decoder/iq_demod/dp_cluster_1/mult_I_sin_out [2]), .B(
        \u_decoder/iq_demod/dp_cluster_1/mult_Q_cos_out [2]), .CI(
        \u_decoder/iq_demod/dp_cluster_1/add_154/carry [2]), .CO(
        \u_decoder/iq_demod/dp_cluster_1/add_154/carry [3]), .S(
        \u_decoder/iq_demod/add_Q_out [2]) );
  ADD32 \u_decoder/iq_demod/dp_cluster_1/add_154/U1_3  ( .A(
        \u_decoder/iq_demod/dp_cluster_1/mult_I_sin_out [3]), .B(
        \u_decoder/iq_demod/dp_cluster_1/mult_Q_cos_out [3]), .CI(
        \u_decoder/iq_demod/dp_cluster_1/add_154/carry [3]), .CO(
        \u_decoder/iq_demod/dp_cluster_1/add_154/carry [4]), .S(
        \u_decoder/iq_demod/add_Q_out [3]) );
  ADD32 \u_decoder/iq_demod/dp_cluster_1/add_154/U1_4  ( .A(
        \u_decoder/iq_demod/dp_cluster_1/mult_I_sin_out [4]), .B(
        \u_decoder/iq_demod/dp_cluster_1/mult_Q_cos_out [4]), .CI(
        \u_decoder/iq_demod/dp_cluster_1/add_154/carry [4]), .CO(
        \u_decoder/iq_demod/dp_cluster_1/add_154/carry [5]), .S(
        \u_decoder/iq_demod/add_Q_out [4]) );
  ADD32 \u_decoder/iq_demod/dp_cluster_1/add_154/U1_5  ( .A(
        \u_decoder/iq_demod/dp_cluster_1/mult_I_sin_out [5]), .B(
        \u_decoder/iq_demod/dp_cluster_1/mult_Q_cos_out [5]), .CI(
        \u_decoder/iq_demod/dp_cluster_1/add_154/carry [5]), .CO(
        \u_decoder/iq_demod/dp_cluster_1/add_154/carry [6]), .S(
        \u_decoder/iq_demod/add_Q_out [5]) );
  ADD32 \u_decoder/iq_demod/dp_cluster_1/add_154/U1_6  ( .A(
        \u_decoder/iq_demod/dp_cluster_1/mult_I_sin_out [6]), .B(
        \u_decoder/iq_demod/dp_cluster_1/mult_Q_cos_out [6]), .CI(
        \u_decoder/iq_demod/dp_cluster_1/add_154/carry [6]), .CO(
        \u_decoder/iq_demod/dp_cluster_1/add_154/carry [7]), .S(
        \u_decoder/iq_demod/add_Q_out [6]) );
  ADD32 \u_outFIFO/r98/U2_1  ( .A(\u_outFIFO/outWriteCount[1] ), .B(n161), 
        .CI(\u_outFIFO/r98/carry [1]), .CO(\u_outFIFO/r98/carry [2]), .S(
        \u_outFIFO/N144 ) );
  ADD32 \u_outFIFO/r98/U2_2  ( .A(\u_outFIFO/outWriteCount[2] ), .B(n167), 
        .CI(\u_outFIFO/r98/carry [2]), .CO(\u_outFIFO/r98/carry [3]), .S(
        \u_outFIFO/N145 ) );
  ADD32 \u_outFIFO/r98/U2_3  ( .A(\u_outFIFO/outWriteCount[3] ), .B(n169), 
        .CI(\u_outFIFO/r98/carry [3]), .CO(\u_outFIFO/r98/carry [4]), .S(
        \u_outFIFO/N146 ) );
  ADD32 \u_outFIFO/r98/U2_4  ( .A(\u_outFIFO/outWriteCount[4] ), .B(n196), 
        .CI(\u_outFIFO/r98/carry [4]), .CO(\u_outFIFO/r98/carry [5]), .S(
        \u_outFIFO/N147 ) );
  ADD32 \u_outFIFO/r98/U2_5  ( .A(\u_outFIFO/outWriteCount[5] ), .B(n220), 
        .CI(\u_outFIFO/r98/carry [5]), .CO(\u_outFIFO/r98/carry [6]), .S(
        \u_outFIFO/N148 ) );
  ADD32 \u_outFIFO/r98/U2_6  ( .A(\u_outFIFO/outWriteCount[6] ), .B(n218), 
        .CI(\u_outFIFO/r98/carry [6]), .CO(\u_outFIFO/r98/carry [7]), .S(
        \u_outFIFO/N149 ) );
  ADD22 \u_outFIFO/add_255/U1_1_1  ( .A(\u_outFIFO/outWriteCount[1] ), .B(
        \u_outFIFO/outWriteCount[0] ), .CO(\u_outFIFO/add_255/carry [2]), .S(
        \u_outFIFO/N120 ) );
  ADD22 \u_outFIFO/add_255/U1_1_2  ( .A(\u_outFIFO/outWriteCount[2] ), .B(
        \u_outFIFO/add_255/carry [2]), .CO(\u_outFIFO/add_255/carry [3]), .S(
        \u_outFIFO/N121 ) );
  ADD22 \u_outFIFO/add_255/U1_1_3  ( .A(\u_outFIFO/outWriteCount[3] ), .B(
        \u_outFIFO/add_255/carry [3]), .CO(\u_outFIFO/add_255/carry [4]), .S(
        \u_outFIFO/N122 ) );
  ADD22 \u_outFIFO/add_255/U1_1_4  ( .A(\u_outFIFO/outWriteCount[4] ), .B(
        \u_outFIFO/add_255/carry [4]), .CO(\u_outFIFO/add_255/carry [5]), .S(
        \u_outFIFO/N123 ) );
  ADD22 \u_outFIFO/add_255/U1_1_5  ( .A(\u_outFIFO/outWriteCount[5] ), .B(
        \u_outFIFO/add_255/carry [5]), .CO(\u_outFIFO/add_255/carry [6]), .S(
        \u_outFIFO/N124 ) );
  ADD22 \u_outFIFO/add_255/U1_1_6  ( .A(\u_outFIFO/outWriteCount[6] ), .B(
        \u_outFIFO/add_255/carry [6]), .CO(\u_outFIFO/add_255/carry [7]), .S(
        \u_outFIFO/N125 ) );
  ADD22 \u_outFIFO/add_256/U1_1_1  ( .A(\u_outFIFO/i_FIFO [1]), .B(
        \u_outFIFO/i_FIFO [0]), .CO(\u_outFIFO/add_256/carry [2]), .S(
        \u_outFIFO/N128 ) );
  ADD22 \u_outFIFO/add_256/U1_1_2  ( .A(\u_outFIFO/i_FIFO [2]), .B(
        \u_outFIFO/add_256/carry [2]), .CO(\u_outFIFO/add_256/carry [3]), .S(
        \u_outFIFO/N129 ) );
  ADD22 \u_outFIFO/add_256/U1_1_3  ( .A(\u_outFIFO/i_FIFO [3]), .B(
        \u_outFIFO/add_256/carry [3]), .CO(\u_outFIFO/add_256/carry [4]), .S(
        \u_outFIFO/N130 ) );
  ADD22 \u_outFIFO/add_256/U1_1_4  ( .A(\u_outFIFO/i_FIFO [4]), .B(
        \u_outFIFO/add_256/carry [4]), .CO(\u_outFIFO/add_256/carry [5]), .S(
        \u_outFIFO/N131 ) );
  ADD22 \u_outFIFO/add_256/U1_1_5  ( .A(\u_outFIFO/i_FIFO [5]), .B(
        \u_outFIFO/add_256/carry [5]), .CO(\u_outFIFO/add_256/carry [6]), .S(
        \u_outFIFO/N132 ) );
  ADD22 \u_outFIFO/add_260/U1_1_1  ( .A(\u_outFIFO/outReadCount[1] ), .B(
        \u_outFIFO/outReadCount[0] ), .CO(\u_outFIFO/add_260/carry [2]), .S(
        \u_outFIFO/N136 ) );
  ADD22 \u_outFIFO/add_260/U1_1_2  ( .A(\u_outFIFO/outReadCount[2] ), .B(
        \u_outFIFO/add_260/carry [2]), .CO(\u_outFIFO/add_260/carry [3]), .S(
        \u_outFIFO/N137 ) );
  ADD22 \u_outFIFO/add_260/U1_1_3  ( .A(\u_outFIFO/outReadCount[3] ), .B(
        \u_outFIFO/add_260/carry [3]), .CO(\u_outFIFO/add_260/carry [4]), .S(
        \u_outFIFO/N138 ) );
  ADD22 \u_outFIFO/add_260/U1_1_4  ( .A(\u_outFIFO/outReadCount[4] ), .B(
        \u_outFIFO/add_260/carry [4]), .CO(\u_outFIFO/add_260/carry [5]), .S(
        \u_outFIFO/N139 ) );
  ADD22 \u_outFIFO/add_260/U1_1_5  ( .A(\u_outFIFO/outReadCount[5] ), .B(
        \u_outFIFO/add_260/carry [5]), .CO(\u_outFIFO/add_260/carry [6]), .S(
        \u_outFIFO/N140 ) );
  ADD22 \u_outFIFO/add_360/U1_1_1  ( .A(\u_outFIFO/N40 ), .B(n1180), .CO(
        \u_outFIFO/add_360/carry [2]), .S(\u_outFIFO/N216 ) );
  ADD22 \u_outFIFO/add_360/U1_1_2  ( .A(n14), .B(\u_outFIFO/add_360/carry [2]), 
        .CO(\u_outFIFO/add_360/carry [3]), .S(\u_outFIFO/N217 ) );
  ADD22 \u_outFIFO/add_360/U1_1_3  ( .A(n1183), .B(
        \u_outFIFO/add_360/carry [3]), .CO(\u_outFIFO/add_360/carry [4]), .S(
        \u_outFIFO/N218 ) );
  ADD22 \u_outFIFO/add_360/U1_1_4  ( .A(\u_outFIFO/N43 ), .B(
        \u_outFIFO/add_360/carry [4]), .CO(\u_outFIFO/add_360/carry [5]), .S(
        \u_outFIFO/N219 ) );
  ADD22 \u_outFIFO/add_360/U1_1_5  ( .A(n761), .B(\u_outFIFO/add_360/carry [5]), .CO(\u_outFIFO/add_360/carry [6]), .S(\u_outFIFO/N220 ) );
  ADD22 \u_coder/add_93/U1_1_1  ( .A(\u_coder/c [1]), .B(\u_coder/c [0]), .CO(
        \u_coder/add_93/carry [2]), .S(\u_coder/N459 ) );
  ADD22 \u_coder/add_93/U1_1_2  ( .A(\u_coder/c [2]), .B(
        \u_coder/add_93/carry [2]), .CO(\u_coder/add_93/carry [3]), .S(
        \u_coder/N460 ) );
  ADD22 \u_coder/add_93/U1_1_3  ( .A(\u_coder/c [3]), .B(
        \u_coder/add_93/carry [3]), .CO(\u_coder/add_93/carry [4]), .S(
        \u_coder/N461 ) );
  ADD22 \u_coder/add_93/U1_1_4  ( .A(\u_coder/c [4]), .B(
        \u_coder/add_93/carry [4]), .CO(\u_coder/add_93/carry [5]), .S(
        \u_coder/N462 ) );
  ADD22 \u_coder/add_93/U1_1_5  ( .A(\u_coder/c [5]), .B(
        \u_coder/add_93/carry [5]), .CO(\u_coder/add_93/carry [6]), .S(
        \u_coder/N463 ) );
  ADD22 \u_coder/add_93/U1_1_6  ( .A(\u_coder/c [6]), .B(
        \u_coder/add_93/carry [6]), .CO(\u_coder/add_93/carry [7]), .S(
        \u_coder/N464 ) );
  ADD22 \u_coder/add_93/U1_1_7  ( .A(\u_coder/c [7]), .B(
        \u_coder/add_93/carry [7]), .CO(\u_coder/add_93/carry [8]), .S(
        \u_coder/N465 ) );
  ADD22 \u_coder/add_93/U1_1_8  ( .A(\u_coder/c [8]), .B(
        \u_coder/add_93/carry [8]), .CO(\u_coder/add_93/carry [9]), .S(
        \u_coder/N466 ) );
  ADD22 \u_coder/add_93/U1_1_9  ( .A(\u_coder/c [9]), .B(
        \u_coder/add_93/carry [9]), .CO(\u_coder/add_93/carry [10]), .S(
        \u_coder/N467 ) );
  ADD22 \u_coder/add_93/U1_1_10  ( .A(\u_coder/c [10]), .B(
        \u_coder/add_93/carry [10]), .CO(\u_coder/add_93/carry [11]), .S(
        \u_coder/N468 ) );
  ADD22 \u_coder/add_93/U1_1_11  ( .A(\u_coder/c [11]), .B(
        \u_coder/add_93/carry [11]), .CO(\u_coder/add_93/carry [12]), .S(
        \u_coder/N469 ) );
  ADD22 \u_coder/add_93/U1_1_12  ( .A(\u_coder/c [12]), .B(
        \u_coder/add_93/carry [12]), .CO(\u_coder/add_93/carry [13]), .S(
        \u_coder/N470 ) );
  ADD22 \u_coder/add_93/U1_1_13  ( .A(\u_coder/c [13]), .B(
        \u_coder/add_93/carry [13]), .CO(\u_coder/add_93/carry [14]), .S(
        \u_coder/N471 ) );
  ADD22 \u_coder/add_93/U1_1_14  ( .A(\u_coder/c [14]), .B(
        \u_coder/add_93/carry [14]), .CO(\u_coder/add_93/carry [15]), .S(
        \u_coder/N472 ) );
  ADD22 \u_coder/add_93/U1_1_15  ( .A(\u_coder/c [15]), .B(
        \u_coder/add_93/carry [15]), .CO(\u_coder/add_93/carry [16]), .S(
        \u_coder/N473 ) );
  ADD22 \u_coder/add_93/U1_1_16  ( .A(\u_coder/c [16]), .B(
        \u_coder/add_93/carry [16]), .CO(\u_coder/add_93/carry [17]), .S(
        \u_coder/N474 ) );
  ADD22 \u_coder/add_93/U1_1_17  ( .A(\u_coder/c [17]), .B(
        \u_coder/add_93/carry [17]), .CO(\u_coder/add_93/carry [18]), .S(
        \u_coder/N475 ) );
  ADD22 \u_coder/add_93/U1_1_18  ( .A(\u_coder/c [18]), .B(
        \u_coder/add_93/carry [18]), .CO(\u_coder/add_93/carry [19]), .S(
        \u_coder/N476 ) );
  ADD22 \u_coder/add_206/U1_1_1  ( .A(\u_coder/i [1]), .B(n763), .CO(
        \u_coder/add_206/carry [2]), .S(\u_coder/N708 ) );
  ADD22 \u_coder/add_206/U1_1_2  ( .A(\u_coder/i [2]), .B(
        \u_coder/add_206/carry [2]), .CO(\u_coder/add_206/carry [3]), .S(
        \u_coder/N709 ) );
  ADD22 \u_coder/add_206/U1_1_3  ( .A(\u_coder/i [3]), .B(
        \u_coder/add_206/carry [3]), .CO(\u_coder/add_206/carry [4]), .S(
        \u_coder/N710 ) );
  ADD22 \u_coder/add_206/U1_1_4  ( .A(\u_coder/i [4]), .B(
        \u_coder/add_206/carry [4]), .CO(\u_coder/add_206/carry [5]), .S(
        \u_coder/N711 ) );
  ADD22 \u_coder/add_206/U1_1_5  ( .A(\u_coder/i [5]), .B(
        \u_coder/add_206/carry [5]), .CO(\u_coder/add_206/carry [6]), .S(
        \u_coder/N712 ) );
  ADD22 \u_coder/add_206/U1_1_6  ( .A(\u_coder/i [6]), .B(
        \u_coder/add_206/carry [6]), .CO(\u_coder/add_206/carry [7]), .S(
        \u_coder/N713 ) );
  ADD22 \u_coder/add_206/U1_1_7  ( .A(\u_coder/i [7]), .B(
        \u_coder/add_206/carry [7]), .CO(\u_coder/add_206/carry [8]), .S(
        \u_coder/N714 ) );
  ADD22 \u_coder/add_206/U1_1_8  ( .A(\u_coder/i [8]), .B(
        \u_coder/add_206/carry [8]), .CO(\u_coder/add_206/carry [9]), .S(
        \u_coder/N715 ) );
  ADD22 \u_coder/add_206/U1_1_9  ( .A(\u_coder/i [9]), .B(
        \u_coder/add_206/carry [9]), .CO(\u_coder/add_206/carry [10]), .S(
        \u_coder/N716 ) );
  ADD22 \u_coder/add_206/U1_1_10  ( .A(\u_coder/i [10]), .B(
        \u_coder/add_206/carry [10]), .CO(\u_coder/add_206/carry [11]), .S(
        \u_coder/N717 ) );
  ADD22 \u_coder/add_206/U1_1_11  ( .A(\u_coder/i [11]), .B(
        \u_coder/add_206/carry [11]), .CO(\u_coder/add_206/carry [12]), .S(
        \u_coder/N718 ) );
  ADD22 \u_coder/add_206/U1_1_12  ( .A(\u_coder/i [12]), .B(
        \u_coder/add_206/carry [12]), .CO(\u_coder/add_206/carry [13]), .S(
        \u_coder/N719 ) );
  ADD22 \u_coder/add_206/U1_1_13  ( .A(\u_coder/i [13]), .B(
        \u_coder/add_206/carry [13]), .CO(\u_coder/add_206/carry [14]), .S(
        \u_coder/N720 ) );
  ADD22 \u_coder/add_206/U1_1_14  ( .A(\u_coder/i [14]), .B(
        \u_coder/add_206/carry [14]), .CO(\u_coder/add_206/carry [15]), .S(
        \u_coder/N721 ) );
  ADD22 \u_coder/add_206/U1_1_15  ( .A(\u_coder/i [15]), .B(
        \u_coder/add_206/carry [15]), .CO(\u_coder/add_206/carry [16]), .S(
        \u_coder/N722 ) );
  ADD22 \u_coder/add_206/U1_1_16  ( .A(\u_coder/i [16]), .B(
        \u_coder/add_206/carry [16]), .CO(\u_coder/add_206/carry [17]), .S(
        \u_coder/N723 ) );
  ADD22 \u_coder/add_206/U1_1_17  ( .A(\u_coder/i [17]), .B(
        \u_coder/add_206/carry [17]), .CO(\u_coder/add_206/carry [18]), .S(
        \u_coder/N724 ) );
  ADD22 \u_coder/add_206/U1_1_18  ( .A(\u_coder/i [18]), .B(
        \u_coder/add_206/carry [18]), .CO(\u_coder/add_206/carry [19]), .S(
        \u_coder/N725 ) );
  ADD22 \u_coder/add_282/U1_1_1  ( .A(n762), .B(\u_coder/j [0]), .CO(
        \u_coder/add_282/carry [2]), .S(\u_coder/N1014 ) );
  ADD22 \u_coder/add_282/U1_1_2  ( .A(\u_coder/j [2]), .B(
        \u_coder/add_282/carry [2]), .CO(\u_coder/add_282/carry [3]), .S(
        \u_coder/N1015 ) );
  ADD22 \u_coder/add_282/U1_1_3  ( .A(\u_coder/j [3]), .B(
        \u_coder/add_282/carry [3]), .CO(\u_coder/add_282/carry [4]), .S(
        \u_coder/N1016 ) );
  ADD22 \u_coder/add_282/U1_1_4  ( .A(\u_coder/j [4]), .B(
        \u_coder/add_282/carry [4]), .CO(\u_coder/add_282/carry [5]), .S(
        \u_coder/N1017 ) );
  ADD22 \u_coder/add_282/U1_1_5  ( .A(\u_coder/j [5]), .B(
        \u_coder/add_282/carry [5]), .CO(\u_coder/add_282/carry [6]), .S(
        \u_coder/N1018 ) );
  ADD22 \u_coder/add_282/U1_1_6  ( .A(\u_coder/j [6]), .B(
        \u_coder/add_282/carry [6]), .CO(\u_coder/add_282/carry [7]), .S(
        \u_coder/N1019 ) );
  ADD22 \u_coder/add_282/U1_1_7  ( .A(\u_coder/j [7]), .B(
        \u_coder/add_282/carry [7]), .CO(\u_coder/add_282/carry [8]), .S(
        \u_coder/N1020 ) );
  ADD22 \u_coder/add_282/U1_1_8  ( .A(\u_coder/j [8]), .B(
        \u_coder/add_282/carry [8]), .CO(\u_coder/add_282/carry [9]), .S(
        \u_coder/N1021 ) );
  ADD22 \u_coder/add_282/U1_1_9  ( .A(\u_coder/j [9]), .B(
        \u_coder/add_282/carry [9]), .CO(\u_coder/add_282/carry [10]), .S(
        \u_coder/N1022 ) );
  ADD22 \u_coder/add_282/U1_1_10  ( .A(\u_coder/j [10]), .B(
        \u_coder/add_282/carry [10]), .CO(\u_coder/add_282/carry [11]), .S(
        \u_coder/N1023 ) );
  ADD22 \u_coder/add_282/U1_1_11  ( .A(\u_coder/j [11]), .B(
        \u_coder/add_282/carry [11]), .CO(\u_coder/add_282/carry [12]), .S(
        \u_coder/N1024 ) );
  ADD22 \u_coder/add_282/U1_1_12  ( .A(\u_coder/j [12]), .B(
        \u_coder/add_282/carry [12]), .CO(\u_coder/add_282/carry [13]), .S(
        \u_coder/N1025 ) );
  ADD22 \u_coder/add_282/U1_1_13  ( .A(\u_coder/j [13]), .B(
        \u_coder/add_282/carry [13]), .CO(\u_coder/add_282/carry [14]), .S(
        \u_coder/N1026 ) );
  ADD22 \u_coder/add_282/U1_1_14  ( .A(\u_coder/j [14]), .B(
        \u_coder/add_282/carry [14]), .CO(\u_coder/add_282/carry [15]), .S(
        \u_coder/N1027 ) );
  ADD22 \u_coder/add_282/U1_1_15  ( .A(\u_coder/j [15]), .B(
        \u_coder/add_282/carry [15]), .CO(\u_coder/add_282/carry [16]), .S(
        \u_coder/N1028 ) );
  ADD22 \u_coder/add_282/U1_1_16  ( .A(\u_coder/j [16]), .B(
        \u_coder/add_282/carry [16]), .CO(\u_coder/add_282/carry [17]), .S(
        \u_coder/N1029 ) );
  ADD22 \u_coder/add_282/U1_1_17  ( .A(\u_coder/j [17]), .B(
        \u_coder/add_282/carry [17]), .CO(\u_coder/add_282/carry [18]), .S(
        \u_coder/N1030 ) );
  ADD22 \u_coder/add_282/U1_1_18  ( .A(\u_coder/j [18]), .B(
        \u_coder/add_282/carry [18]), .CO(\u_coder/add_282/carry [19]), .S(
        \u_coder/N1031 ) );
  ADD32 \u_inFIFO/r96/U2_1  ( .A(\u_inFIFO/outWriteCount[1] ), .B(n126), .CI(
        \u_inFIFO/r96/carry [1]), .CO(\u_inFIFO/r96/carry [2]), .S(
        \u_inFIFO/N134 ) );
  ADD32 \u_inFIFO/r96/U2_2  ( .A(\u_inFIFO/outWriteCount[2] ), .B(n166), .CI(
        \u_inFIFO/r96/carry [2]), .CO(\u_inFIFO/r96/carry [3]), .S(
        \u_inFIFO/N135 ) );
  ADD32 \u_inFIFO/r96/U2_3  ( .A(\u_inFIFO/outWriteCount[3] ), .B(n168), .CI(
        \u_inFIFO/r96/carry [3]), .CO(\u_inFIFO/r96/carry [4]), .S(
        \u_inFIFO/N136 ) );
  ADD32 \u_inFIFO/r96/U2_4  ( .A(\u_inFIFO/outWriteCount[4] ), .B(n162), .CI(
        \u_inFIFO/r96/carry [4]), .CO(\u_inFIFO/r96/carry [5]), .S(
        \u_inFIFO/N137 ) );
  ADD32 \u_inFIFO/r96/U2_5  ( .A(\u_inFIFO/outWriteCount[5] ), .B(n219), .CI(
        \u_inFIFO/r96/carry [5]), .CO(\u_inFIFO/r96/carry [6]), .S(
        \u_inFIFO/N138 ) );
  ADD32 \u_inFIFO/r96/U2_6  ( .A(\u_inFIFO/outWriteCount[6] ), .B(n217), .CI(
        \u_inFIFO/r96/carry [6]), .CO(\u_inFIFO/r96/carry [7]), .S(
        \u_inFIFO/N139 ) );
  ADD22 \u_inFIFO/add_252/U1_1_1  ( .A(\u_inFIFO/outReadCount[1] ), .B(
        \u_inFIFO/outReadCount[0] ), .CO(\u_inFIFO/add_252/carry [2]), .S(
        \u_inFIFO/N119 ) );
  ADD22 \u_inFIFO/add_252/U1_1_2  ( .A(\u_inFIFO/outReadCount[2] ), .B(
        \u_inFIFO/add_252/carry [2]), .CO(\u_inFIFO/add_252/carry [3]), .S(
        \u_inFIFO/N120 ) );
  ADD22 \u_inFIFO/add_252/U1_1_3  ( .A(\u_inFIFO/outReadCount[3] ), .B(
        \u_inFIFO/add_252/carry [3]), .CO(\u_inFIFO/add_252/carry [4]), .S(
        \u_inFIFO/N121 ) );
  ADD22 \u_inFIFO/add_252/U1_1_4  ( .A(\u_inFIFO/outReadCount[4] ), .B(
        \u_inFIFO/add_252/carry [4]), .CO(\u_inFIFO/add_252/carry [5]), .S(
        \u_inFIFO/N122 ) );
  ADD22 \u_inFIFO/add_252/U1_1_5  ( .A(\u_inFIFO/outReadCount[5] ), .B(
        \u_inFIFO/add_252/carry [5]), .CO(\u_inFIFO/add_252/carry [6]), .S(
        \u_inFIFO/N123 ) );
  ADD22 \u_inFIFO/add_253/U1_1_1  ( .A(\u_inFIFO/N38 ), .B(n13), .CO(
        \u_inFIFO/add_253/carry [2]), .S(\u_inFIFO/N126 ) );
  ADD22 \u_inFIFO/add_253/U1_1_2  ( .A(n15), .B(\u_inFIFO/add_253/carry [2]), 
        .CO(\u_inFIFO/add_253/carry [3]), .S(\u_inFIFO/N127 ) );
  ADD22 \u_inFIFO/add_253/U1_1_3  ( .A(n1202), .B(\u_inFIFO/add_253/carry [3]), 
        .CO(\u_inFIFO/add_253/carry [4]), .S(\u_inFIFO/N128 ) );
  ADD22 \u_inFIFO/add_253/U1_1_4  ( .A(n765), .B(\u_inFIFO/add_253/carry [4]), 
        .CO(\u_inFIFO/add_253/carry [5]), .S(\u_inFIFO/N129 ) );
  ADD22 \u_inFIFO/add_253/U1_1_5  ( .A(n49), .B(\u_inFIFO/add_253/carry [5]), 
        .CO(\u_inFIFO/add_253/carry [6]), .S(\u_inFIFO/N130 ) );
  ADD22 \u_inFIFO/add_263/U1_1_1  ( .A(\u_inFIFO/outWriteCount[1] ), .B(
        \u_inFIFO/outWriteCount[0] ), .CO(\u_inFIFO/add_263/carry [2]), .S(
        \u_inFIFO/N143 ) );
  ADD22 \u_inFIFO/add_263/U1_1_2  ( .A(\u_inFIFO/outWriteCount[2] ), .B(
        \u_inFIFO/add_263/carry [2]), .CO(\u_inFIFO/add_263/carry [3]), .S(
        \u_inFIFO/N144 ) );
  ADD22 \u_inFIFO/add_263/U1_1_3  ( .A(\u_inFIFO/outWriteCount[3] ), .B(
        \u_inFIFO/add_263/carry [3]), .CO(\u_inFIFO/add_263/carry [4]), .S(
        \u_inFIFO/N145 ) );
  ADD22 \u_inFIFO/add_263/U1_1_4  ( .A(\u_inFIFO/outWriteCount[4] ), .B(
        \u_inFIFO/add_263/carry [4]), .CO(\u_inFIFO/add_263/carry [5]), .S(
        \u_inFIFO/N146 ) );
  ADD22 \u_inFIFO/add_263/U1_1_5  ( .A(\u_inFIFO/outWriteCount[5] ), .B(
        \u_inFIFO/add_263/carry [5]), .CO(\u_inFIFO/add_263/carry [6]), .S(
        \u_inFIFO/N147 ) );
  ADD22 \u_inFIFO/add_263/U1_1_6  ( .A(\u_inFIFO/outWriteCount[6] ), .B(
        \u_inFIFO/add_263/carry [6]), .CO(\u_inFIFO/add_263/carry [7]), .S(
        \u_inFIFO/N148 ) );
  ADD22 \u_inFIFO/add_357/U1_1_1  ( .A(\u_inFIFO/j_FIFO [1]), .B(
        \u_inFIFO/j_FIFO [0]), .CO(\u_inFIFO/add_357/carry [2]), .S(
        \u_inFIFO/N212 ) );
  ADD22 \u_inFIFO/add_357/U1_1_2  ( .A(\u_inFIFO/j_FIFO [2]), .B(
        \u_inFIFO/add_357/carry [2]), .CO(\u_inFIFO/add_357/carry [3]), .S(
        \u_inFIFO/N213 ) );
  ADD22 \u_inFIFO/add_357/U1_1_3  ( .A(\u_inFIFO/j_FIFO [3]), .B(
        \u_inFIFO/add_357/carry [3]), .CO(\u_inFIFO/add_357/carry [4]), .S(
        \u_inFIFO/N214 ) );
  ADD22 \u_inFIFO/add_357/U1_1_4  ( .A(\u_inFIFO/j_FIFO [4]), .B(
        \u_inFIFO/add_357/carry [4]), .CO(\u_inFIFO/add_357/carry [5]), .S(
        \u_inFIFO/N215 ) );
  ADD22 \u_inFIFO/add_357/U1_1_5  ( .A(\u_inFIFO/j_FIFO [5]), .B(
        \u_inFIFO/add_357/carry [5]), .CO(\u_inFIFO/add_357/carry [6]), .S(
        \u_inFIFO/N216 ) );
  DF3 \u_inFIFO/sigOutData_reg  ( .D(\u_inFIFO/n572 ), .C(inClock), .Q(
        \sig_MUX_inMUX4[0] ), .QN(\u_inFIFO/n200 ) );
  DF3 \u_inFIFO/j_FIFO_reg[6]  ( .D(n1965), .C(inClock), .Q(
        \u_inFIFO/j_FIFO [6]), .QN(\u_inFIFO/n201 ) );
  DF3 \u_inFIFO/j_FIFO_reg[5]  ( .D(n1964), .C(inClock), .Q(
        \u_inFIFO/j_FIFO [5]), .QN(\u_inFIFO/n202 ) );
  DF3 \u_inFIFO/j_FIFO_reg[4]  ( .D(n1963), .C(inClock), .Q(
        \u_inFIFO/j_FIFO [4]), .QN(\u_inFIFO/n203 ) );
  DF3 \u_inFIFO/j_FIFO_reg[3]  ( .D(n1962), .C(inClock), .Q(
        \u_inFIFO/j_FIFO [3]), .QN(\u_inFIFO/n204 ) );
  DF3 \u_inFIFO/j_FIFO_reg[2]  ( .D(n1961), .C(inClock), .Q(
        \u_inFIFO/j_FIFO [2]), .QN(\u_inFIFO/n205 ) );
  DF3 \u_inFIFO/j_FIFO_reg[1]  ( .D(n1960), .C(inClock), .Q(
        \u_inFIFO/j_FIFO [1]), .QN(\u_inFIFO/n206 ) );
  DF3 \u_inFIFO/j_FIFO_reg[0]  ( .D(n1959), .C(inClock), .Q(
        \u_inFIFO/j_FIFO [0]), .QN(\u_inFIFO/n207 ) );
  DF3 \u_inFIFO/currentState_reg[1]  ( .D(\u_inFIFO/N48 ), .C(inClock), .Q(
        \u_inFIFO/currentState [1]), .QN(\u_inFIFO/n176 ) );
  DF3 \u_inFIFO/currentState_reg[2]  ( .D(\u_inFIFO/N49 ), .C(inClock), .QN(
        \u_inFIFO/n173 ) );
  DF3 \u_inFIFO/currentState_reg[0]  ( .D(\u_inFIFO/N47 ), .C(inClock), .Q(
        \u_inFIFO/currentState [0]), .QN(\u_inFIFO/n177 ) );
  DF3 \u_inFIFO/k_FIFO_reg[1]  ( .D(\u_inFIFO/n573 ), .C(inClock), .Q(
        \u_inFIFO/N45 ), .QN(\u_inFIFO/n197 ) );
  DF3 \u_inFIFO/k_FIFO_reg[0]  ( .D(\u_inFIFO/n574 ), .C(inClock), .Q(
        \u_inFIFO/N44 ), .QN(\u_inFIFO/n198 ) );
  DF3 \u_inFIFO/currentState_reg[3]  ( .D(\u_inFIFO/N50 ), .C(inClock), .Q(
        \u_inFIFO/currentState [3]), .QN(\u_inFIFO/n154 ) );
  DF3 \u_inFIFO/sigWRCOUNT_reg[5]  ( .D(\u_inFIFO/n579 ), .C(inClock), .Q(
        \u_inFIFO/outWriteCount[5] ), .QN(\u_inFIFO/n183 ) );
  DF3 \u_inFIFO/sigWRCOUNT_reg[4]  ( .D(\u_inFIFO/n578 ), .C(inClock), .Q(
        \u_inFIFO/outWriteCount[4] ), .QN(\u_inFIFO/n184 ) );
  DF3 \u_inFIFO/sigWRCOUNT_reg[3]  ( .D(\u_inFIFO/n577 ), .C(inClock), .Q(
        \u_inFIFO/outWriteCount[3] ), .QN(\u_inFIFO/n185 ) );
  DF3 \u_inFIFO/sigWRCOUNT_reg[2]  ( .D(\u_inFIFO/n576 ), .C(inClock), .Q(
        \u_inFIFO/outWriteCount[2] ), .QN(\u_inFIFO/n186 ) );
  DF3 \u_inFIFO/sigWRCOUNT_reg[1]  ( .D(\u_inFIFO/n575 ), .C(inClock), .Q(
        \u_inFIFO/outWriteCount[1] ), .QN(\u_inFIFO/n187 ) );
  DF3 \u_inFIFO/sigWRCOUNT_reg[0]  ( .D(\u_inFIFO/n581 ), .C(inClock), .Q(
        \u_inFIFO/outWriteCount[0] ), .QN(\u_inFIFO/n188 ) );
  DF3 \u_inFIFO/sigWRCOUNT_reg[6]  ( .D(\u_inFIFO/n580 ), .C(inClock), .Q(
        \u_inFIFO/outWriteCount[6] ), .QN(\u_inFIFO/n182 ) );
  DF3 \u_inFIFO/sigRDCOUNT_reg[5]  ( .D(n1827), .C(inClock), .Q(
        \u_inFIFO/outReadCount[5] ), .QN(n219) );
  DF3 \u_inFIFO/sigRDCOUNT_reg[4]  ( .D(n1826), .C(inClock), .Q(
        \u_inFIFO/outReadCount[4] ), .QN(n162) );
  DF3 \u_inFIFO/sigRDCOUNT_reg[3]  ( .D(n1825), .C(inClock), .Q(
        \u_inFIFO/outReadCount[3] ), .QN(n168) );
  DF3 \u_inFIFO/sigRDCOUNT_reg[2]  ( .D(n1824), .C(inClock), .Q(
        \u_inFIFO/outReadCount[2] ), .QN(n166) );
  DF3 \u_inFIFO/sigRDCOUNT_reg[1]  ( .D(n1823), .C(inClock), .Q(
        \u_inFIFO/outReadCount[1] ), .QN(n126) );
  DF3 \u_inFIFO/sigRDCOUNT_reg[0]  ( .D(n1822), .C(inClock), .Q(
        \u_inFIFO/outReadCount[0] ), .QN(n129) );
  DF3 \u_inFIFO/sigRDCOUNT_reg[6]  ( .D(n1821), .C(inClock), .Q(
        \u_inFIFO/outReadCount[6] ), .QN(n217) );
  DF3 \u_inFIFO/sigWRCOUNT_reg[7]  ( .D(\u_inFIFO/n582 ), .C(inClock), .Q(
        \u_inFIFO/outWriteCount[7] ), .QN(\u_inFIFO/n179 ) );
  DF3 \u_inFIFO/i_FIFO_reg[6]  ( .D(n1820), .C(inClock), .Q(\u_inFIFO/N43 ) );
  DF3 \u_inFIFO/i_FIFO_reg[5]  ( .D(n1819), .C(inClock), .Q(n49) );
  DF3 \u_inFIFO/i_FIFO_reg[4]  ( .D(n1818), .C(inClock), .Q(\u_inFIFO/N41 ) );
  DF3 \u_inFIFO/i_FIFO_reg[3]  ( .D(n1817), .C(inClock), .Q(\u_inFIFO/N40 ) );
  DF3 \u_inFIFO/i_FIFO_reg[2]  ( .D(n1816), .C(inClock), .Q(n15) );
  DF3 \u_inFIFO/i_FIFO_reg[1]  ( .D(n1815), .C(inClock), .Q(\u_inFIFO/N38 ) );
  DF3 \u_inFIFO/i_FIFO_reg[0]  ( .D(n1814), .C(inClock), .Q(n13), .QN(n198) );
  DF3 \u_inFIFO/sigEnableCounter_reg  ( .D(\u_inFIFO/N196 ), .C(inClock), .Q(
        \u_inFIFO/sigEnableCounter ) );
  DF3 \u_coder/o_ready_reg  ( .D(\u_coder/n346 ), .C(inClock), .Q(
        \sig_MUX_inMUX3[0] ) );
  DF3 \u_coder/o_sinQ_four_reg[1]  ( .D(\u_coder/n343 ), .C(inClock), .Q(
        sig_coder_outSinQMasked[1]) );
  DF3 \u_coder/o_sinQ_four_reg[2]  ( .D(\u_coder/n342 ), .C(inClock), .Q(
        sig_coder_outSinQMasked[2]) );
  DF3 \u_coder/o_sinQ_reg[0]  ( .D(\u_coder/n339 ), .C(inClock), .Q(
        sig_coder_outSinQ[0]) );
  DF3 \u_coder/o_sinQ_reg[1]  ( .D(\u_coder/n338 ), .C(inClock), .Q(
        sig_coder_outSinQ[1]) );
  DF3 \u_coder/o_sinQ_reg[2]  ( .D(\u_coder/n337 ), .C(inClock), .Q(
        sig_coder_outSinQ[2]) );
  DF3 \u_coder/o_sinQ_reg[3]  ( .D(n1810), .C(inClock), .Q(
        sig_coder_outSinQ[3]) );
  DF3 \u_coder/o_sinQ_four_reg[3]  ( .D(\u_coder/n341 ), .C(inClock), .Q(
        sig_coder_outSinQMasked[3]) );
  DF3 \u_coder/sin_was_positiveQ_reg  ( .D(\u_coder/n345 ), .C(inClock), .Q(
        \u_coder/sin_was_positiveQ ), .QN(\u_coder/n125 ) );
  DF3 \u_coder/isPositiveQ_reg  ( .D(n1812), .C(inClock), .Q(
        \u_coder/isPositiveQ ), .QN(\u_coder/n127 ) );
  DF3 \u_coder/o_sinQ_four_reg[0]  ( .D(\u_coder/n344 ), .C(inClock), .Q(
        sig_coder_outSinQMasked[0]) );
  DF3 \u_coder/o_sinI_four_reg[0]  ( .D(\u_coder/n350 ), .C(inClock), .Q(
        sig_coder_outSinIMasked[0]) );
  DF3 \u_coder/o_sinI_four_reg[1]  ( .D(\u_coder/n349 ), .C(inClock), .Q(
        sig_coder_outSinIMasked[1]) );
  DF3 \u_coder/o_sinI_four_reg[2]  ( .D(\u_coder/n348 ), .C(inClock), .Q(
        sig_coder_outSinIMasked[2]) );
  DF3 \u_coder/o_sinI_four_reg[3]  ( .D(\u_coder/n347 ), .C(inClock), .Q(
        sig_coder_outSinIMasked[3]) );
  DF3 \u_coder/o_sinI_reg[3]  ( .D(\u_coder/n335 ), .C(inClock), .Q(
        sig_coder_outSinI[3]), .QN(\u_coder/n129 ) );
  DF3 \u_coder/o_sinI_reg[0]  ( .D(\u_coder/n336 ), .C(inClock), .Q(
        sig_coder_outSinI[0]) );
  DF3 \u_coder/o_sinI_reg[1]  ( .D(n1808), .C(inClock), .Q(
        sig_coder_outSinI[1]) );
  DF3 \u_coder/o_sinI_reg[2]  ( .D(n1807), .C(inClock), .Q(
        sig_coder_outSinI[2]) );
  DF3 \u_coder/sin_was_positiveI_reg  ( .D(\u_coder/n351 ), .C(inClock), .QN(
        \u_coder/n123 ) );
  DF3 \u_coder/isPositiveI_reg  ( .D(\u_coder/n352 ), .C(inClock), .Q(
        \u_coder/isPositiveI ), .QN(\u_coder/n126 ) );
  DF3 \u_coder/old_i_data_reg  ( .D(\u_coder/n353 ), .C(inClock), .Q(
        \u_coder/old_i_data ), .QN(n385) );
  DF3 \u_coder/i_reg[18]  ( .D(n1954), .C(inClock), .Q(\u_coder/i [18]) );
  DF3 \u_coder/i_reg[17]  ( .D(n1953), .C(inClock), .Q(\u_coder/i [17]) );
  DF3 \u_coder/i_reg[16]  ( .D(n1952), .C(inClock), .Q(\u_coder/i [16]) );
  DF3 \u_coder/i_reg[15]  ( .D(n1951), .C(inClock), .Q(\u_coder/i [15]) );
  DF3 \u_coder/i_reg[14]  ( .D(n1950), .C(inClock), .Q(\u_coder/i [14]) );
  DF3 \u_coder/i_reg[13]  ( .D(n1949), .C(inClock), .Q(\u_coder/i [13]) );
  DF3 \u_coder/i_reg[12]  ( .D(n1948), .C(inClock), .Q(\u_coder/i [12]) );
  DF3 \u_coder/i_reg[11]  ( .D(n1947), .C(inClock), .Q(\u_coder/i [11]) );
  DF3 \u_coder/i_reg[10]  ( .D(n1946), .C(inClock), .Q(\u_coder/i [10]) );
  DF3 \u_coder/i_reg[9]  ( .D(n1945), .C(inClock), .Q(\u_coder/i [9]) );
  DF3 \u_coder/i_reg[8]  ( .D(n1944), .C(inClock), .Q(\u_coder/i [8]) );
  DF3 \u_coder/i_reg[7]  ( .D(n1943), .C(inClock), .Q(\u_coder/i [7]) );
  DF3 \u_coder/i_reg[6]  ( .D(n1942), .C(inClock), .Q(\u_coder/i [6]) );
  DF3 \u_coder/i_reg[5]  ( .D(n1941), .C(inClock), .Q(\u_coder/i [5]) );
  DF3 \u_coder/i_reg[4]  ( .D(n1940), .C(inClock), .Q(\u_coder/i [4]) );
  DF3 \u_coder/i_reg[3]  ( .D(n1939), .C(inClock), .Q(\u_coder/i [3]), .QN(
        \u_coder/n101 ) );
  DF3 \u_coder/i_reg[2]  ( .D(n1938), .C(inClock), .Q(\u_coder/i [2]), .QN(
        \u_coder/n103 ) );
  DF3 \u_coder/i_reg[1]  ( .D(n1937), .C(inClock), .Q(\u_coder/i [1]), .QN(
        \u_coder/n104 ) );
  DF3 \u_coder/i_reg[0]  ( .D(n1936), .C(inClock), .Q(\u_coder/i [0]), .QN(
        \u_coder/n105 ) );
  DF3 \u_coder/is9_reg  ( .D(\u_coder/n340 ), .C(inClock), .Q(\u_coder/is9 ), 
        .QN(\u_coder/n128 ) );
  DF3 \u_coder/i_reg[19]  ( .D(n1935), .C(inClock), .Q(\u_coder/i [19]) );
  DF3 \u_coder/stateI_reg[0]  ( .D(\u_coder/N499 ), .C(inClock), .Q(
        \u_coder/stateI[0] ), .QN(\u_coder/n91 ) );
  DF3 \u_coder/next_stateI_reg[0]  ( .D(\u_coder/n354 ), .C(inClock), .QN(
        \u_coder/n130 ) );
  DF3 \u_coder/IorQ_reg  ( .D(\u_coder/n355 ), .C(inClock), .Q(\u_coder/IorQ )
         );
  DF3 \u_coder/j_reg[18]  ( .D(n1934), .C(inClock), .Q(\u_coder/j [18]) );
  DF3 \u_coder/j_reg[17]  ( .D(n1933), .C(inClock), .Q(\u_coder/j [17]) );
  DF3 \u_coder/j_reg[16]  ( .D(n1932), .C(inClock), .Q(\u_coder/j [16]) );
  DF3 \u_coder/j_reg[15]  ( .D(n1931), .C(inClock), .Q(\u_coder/j [15]) );
  DF3 \u_coder/j_reg[14]  ( .D(n1930), .C(inClock), .Q(\u_coder/j [14]) );
  DF3 \u_coder/j_reg[13]  ( .D(n1929), .C(inClock), .Q(\u_coder/j [13]) );
  DF3 \u_coder/j_reg[12]  ( .D(n1928), .C(inClock), .Q(\u_coder/j [12]) );
  DF3 \u_coder/j_reg[11]  ( .D(n1927), .C(inClock), .Q(\u_coder/j [11]) );
  DF3 \u_coder/j_reg[10]  ( .D(n1926), .C(inClock), .Q(\u_coder/j [10]) );
  DF3 \u_coder/j_reg[9]  ( .D(n1925), .C(inClock), .Q(\u_coder/j [9]) );
  DF3 \u_coder/j_reg[8]  ( .D(n1924), .C(inClock), .Q(\u_coder/j [8]) );
  DF3 \u_coder/j_reg[7]  ( .D(n1923), .C(inClock), .Q(\u_coder/j [7]) );
  DF3 \u_coder/j_reg[6]  ( .D(n1922), .C(inClock), .Q(\u_coder/j [6]) );
  DF3 \u_coder/j_reg[5]  ( .D(n1921), .C(inClock), .Q(\u_coder/j [5]) );
  DF3 \u_coder/j_reg[4]  ( .D(n1920), .C(inClock), .Q(\u_coder/j [4]) );
  DF3 \u_coder/j_reg[3]  ( .D(n1919), .C(inClock), .Q(\u_coder/j [3]), .QN(
        \u_coder/n117 ) );
  DF3 \u_coder/j_reg[2]  ( .D(n1918), .C(inClock), .Q(\u_coder/j [2]), .QN(
        \u_coder/n118 ) );
  DF3 \u_coder/j_reg[1]  ( .D(n1917), .C(inClock), .Q(\u_coder/j [1]) );
  DF3 \u_coder/j_reg[0]  ( .D(n1916), .C(inClock), .Q(\u_coder/j [0]), .QN(
        \u_coder/n120 ) );
  DF3 \u_coder/j_reg[19]  ( .D(n1915), .C(inClock), .Q(\u_coder/j [19]) );
  DF3 \u_coder/stateQ_reg[0]  ( .D(\u_coder/N501 ), .C(inClock), .Q(
        \u_coder/stateQ[0] ), .QN(\u_coder/n94 ) );
  DF3 \u_coder/next_stateQ_reg[0]  ( .D(\u_coder/n356 ), .C(inClock), .QN(
        \u_coder/n131 ) );
  DF3 \u_coder/clk_10M_reg  ( .D(n2186), .C(inClock), .Q(\u_coder/clk_10M ) );
  DF3 \u_coder/c_reg[19]  ( .D(\u_coder/N522 ), .C(inClock), .Q(
        \u_coder/c [19]) );
  DF3 \u_coder/c_reg[18]  ( .D(\u_coder/N521 ), .C(inClock), .Q(
        \u_coder/c [18]) );
  DF3 \u_coder/c_reg[17]  ( .D(\u_coder/N520 ), .C(inClock), .Q(
        \u_coder/c [17]) );
  DF3 \u_coder/c_reg[16]  ( .D(\u_coder/N519 ), .C(inClock), .Q(
        \u_coder/c [16]) );
  DF3 \u_coder/c_reg[15]  ( .D(\u_coder/N518 ), .C(inClock), .Q(
        \u_coder/c [15]) );
  DF3 \u_coder/c_reg[14]  ( .D(\u_coder/N517 ), .C(inClock), .Q(
        \u_coder/c [14]) );
  DF3 \u_coder/c_reg[13]  ( .D(\u_coder/N516 ), .C(inClock), .Q(
        \u_coder/c [13]) );
  DF3 \u_coder/c_reg[12]  ( .D(\u_coder/N515 ), .C(inClock), .Q(
        \u_coder/c [12]) );
  DF3 \u_coder/c_reg[11]  ( .D(\u_coder/N514 ), .C(inClock), .Q(
        \u_coder/c [11]) );
  DF3 \u_coder/c_reg[10]  ( .D(\u_coder/N513 ), .C(inClock), .Q(
        \u_coder/c [10]) );
  DF3 \u_coder/c_reg[9]  ( .D(\u_coder/N512 ), .C(inClock), .Q(\u_coder/c [9])
         );
  DF3 \u_coder/c_reg[8]  ( .D(\u_coder/N511 ), .C(inClock), .Q(\u_coder/c [8])
         );
  DF3 \u_coder/c_reg[7]  ( .D(\u_coder/N510 ), .C(inClock), .Q(\u_coder/c [7])
         );
  DF3 \u_coder/c_reg[6]  ( .D(\u_coder/N509 ), .C(inClock), .Q(\u_coder/c [6])
         );
  DF3 \u_coder/c_reg[5]  ( .D(\u_coder/N508 ), .C(inClock), .Q(\u_coder/c [5])
         );
  DF3 \u_coder/c_reg[4]  ( .D(\u_coder/N507 ), .C(inClock), .Q(\u_coder/c [4])
         );
  DF3 \u_coder/c_reg[3]  ( .D(\u_coder/N506 ), .C(inClock), .Q(\u_coder/c [3])
         );
  DF3 \u_coder/c_reg[2]  ( .D(\u_coder/N505 ), .C(inClock), .Q(\u_coder/c [2])
         );
  DF3 \u_coder/c_reg[1]  ( .D(\u_coder/N504 ), .C(inClock), .Q(\u_coder/c [1])
         );
  DF3 \u_coder/c_reg[0]  ( .D(\u_coder/N503 ), .C(inClock), .Q(\u_coder/c [0]), 
        .QN(\u_coder/n33 ) );
  DF3 \u_cordic/o_dir_reg  ( .D(\u_cordic/n32 ), .C(inClock), .Q(
        \sig_MUX_inMUX14[0] ), .QN(\u_cordic/n12 ) );
  DF3 \u_cordic/I_reg[0]  ( .D(n2115), .C(inClock), .Q(\u_cordic/I [0]) );
  DF3 \u_cordic/I_reg[1]  ( .D(n2113), .C(inClock), .Q(\u_cordic/I [1]) );
  DF3 \u_cordic/I_reg[2]  ( .D(n2111), .C(inClock), .Q(\u_cordic/I [2]) );
  DF3 \u_cordic/I_reg[3]  ( .D(n2109), .C(inClock), .Q(\u_cordic/I [3]) );
  DF3 \u_cordic/Q_reg[0]  ( .D(n2123), .C(inClock), .Q(\u_cordic/Q [0]) );
  DF3 \u_cordic/Q_reg[1]  ( .D(n2121), .C(inClock), .Q(\u_cordic/Q [1]) );
  DF3 \u_cordic/Q_reg[2]  ( .D(n2119), .C(inClock), .Q(\u_cordic/Q [2]) );
  DF3 \u_cordic/Q_reg[3]  ( .D(n2117), .C(inClock), .Q(\u_cordic/Q [3]) );
  DF3 \u_cordic/present_state_reg[2]  ( .D(\u_cordic/N16 ), .C(inClock), .Q(
        \u_cordic/present_state [2]), .QN(\u_cordic/n9 ) );
  DF3 \u_cordic/present_state_reg[1]  ( .D(\u_cordic/N15 ), .C(inClock), .Q(
        \u_cordic/present_state [1]), .QN(\u_cordic/n10 ) );
  DF3 \u_cordic/present_state_reg[0]  ( .D(\u_cordic/N14 ), .C(inClock), .Q(
        \u_cordic/present_state [0]), .QN(\u_cordic/n11 ) );
  DF3 \u_cdr/dir_reg  ( .D(\u_cdr/n50 ), .C(inClock), .Q(\u_cdr/dir ) );
  DF3 \u_cdr/cnt_reg[2]  ( .D(\u_cdr/n52 ), .C(inClock), .QN(\u_cdr/n16 ) );
  DF3 \u_cdr/cnt_reg[1]  ( .D(\u_cdr/n51 ), .C(inClock), .Q(\u_cdr/cnt [1]), 
        .QN(\u_cdr/n17 ) );
  JK3 \u_cdr/cnt_reg[0]  ( .J(\u_cdr/n33 ), .K(\u_cdr/n35 ), .C(inClock), .Q(
        \u_cdr/cnt [0]), .QN(\u_cdr/n18 ) );
  DF3 \u_cdr/flag_reg  ( .D(\u_cdr/n53 ), .C(inClock), .Q(\u_cdr/flag ), .QN(
        n320) );
  DF3 \u_cdr/cnt_d_reg[1]  ( .D(\u_cdr/n54 ), .C(inClock), .Q(\u_cdr/cnt_d [1]), .QN(\u_cdr/n14 ) );
  DF3 \u_cdr/cnt_d_reg[0]  ( .D(\u_cdr/n55 ), .C(inClock), .Q(\u_cdr/cnt_d [0]), .QN(\u_cdr/n15 ) );
  DF3 \u_cdr/cnt_in_reg[3]  ( .D(\u_cdr/n56 ), .C(inClock), .Q(
        \u_cdr/cnt_in [3]), .QN(n50) );
  DF3 \u_cdr/cnt_in_reg[2]  ( .D(\u_cdr/n57 ), .C(inClock), .Q(
        \u_cdr/cnt_in [2]), .QN(n290) );
  DF3 \u_cdr/cnt_in_reg[1]  ( .D(\u_cdr/n58 ), .C(inClock), .Q(
        \u_cdr/cnt_in [1]), .QN(n20) );
  DF3 \u_cdr/cnt_in_reg[0]  ( .D(\u_cdr/n59 ), .C(inClock), .Q(
        \u_cdr/cnt_in [0]), .QN(n289) );
  DF3 \u_outFIFO/sigOutData_reg[0]  ( .D(n1581), .C(inClock), .Q(
        sig_outFIFO_outData[0]) );
  DF3 \u_outFIFO/sigOutData_reg[1]  ( .D(n1582), .C(inClock), .Q(
        sig_outFIFO_outData[1]) );
  DF3 \u_outFIFO/sigOutData_reg[2]  ( .D(n1583), .C(inClock), .Q(
        sig_outFIFO_outData[2]) );
  DF3 \u_outFIFO/sigOutData_reg[3]  ( .D(n1584), .C(inClock), .Q(
        sig_outFIFO_outData[3]) );
  DF3 \u_outFIFO/FIFO_reg[75][3]  ( .D(\u_outFIFO/n1161 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[75][3] ) );
  DF3 \u_outFIFO/FIFO_reg[76][0]  ( .D(\u_outFIFO/n1162 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[76][0] ) );
  DF3 \u_outFIFO/FIFO_reg[76][1]  ( .D(\u_outFIFO/n1163 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[76][1] ) );
  DF3 \u_outFIFO/FIFO_reg[76][2]  ( .D(\u_outFIFO/n1164 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[76][2] ) );
  DF3 \u_outFIFO/FIFO_reg[76][3]  ( .D(\u_outFIFO/n1165 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[76][3] ) );
  DF3 \u_outFIFO/FIFO_reg[77][0]  ( .D(\u_outFIFO/n1166 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[77][0] ) );
  DF3 \u_outFIFO/FIFO_reg[77][1]  ( .D(\u_outFIFO/n1167 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[77][1] ) );
  DF3 \u_outFIFO/FIFO_reg[77][2]  ( .D(\u_outFIFO/n1168 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[77][2] ) );
  DF3 \u_outFIFO/FIFO_reg[77][3]  ( .D(\u_outFIFO/n1169 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[77][3] ) );
  DF3 \u_outFIFO/FIFO_reg[78][0]  ( .D(\u_outFIFO/n1170 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[78][0] ) );
  DF3 \u_outFIFO/FIFO_reg[78][1]  ( .D(\u_outFIFO/n1171 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[78][1] ) );
  DF3 \u_outFIFO/FIFO_reg[78][2]  ( .D(\u_outFIFO/n1172 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[78][2] ) );
  DF3 \u_outFIFO/FIFO_reg[78][3]  ( .D(\u_outFIFO/n1173 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[78][3] ) );
  DF3 \u_outFIFO/FIFO_reg[79][0]  ( .D(\u_outFIFO/n1174 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[79][0] ) );
  DF3 \u_outFIFO/FIFO_reg[79][1]  ( .D(\u_outFIFO/n1175 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[79][1] ) );
  DF3 \u_outFIFO/FIFO_reg[79][2]  ( .D(\u_outFIFO/n1176 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[79][2] ) );
  DF3 \u_outFIFO/FIFO_reg[79][3]  ( .D(\u_outFIFO/n1177 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[79][3] ) );
  DF3 \u_outFIFO/FIFO_reg[80][0]  ( .D(\u_outFIFO/n1178 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[80][0] ) );
  DF3 \u_outFIFO/FIFO_reg[80][1]  ( .D(\u_outFIFO/n1179 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[80][1] ) );
  DF3 \u_outFIFO/FIFO_reg[80][2]  ( .D(\u_outFIFO/n1180 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[80][2] ) );
  DF3 \u_outFIFO/FIFO_reg[80][3]  ( .D(\u_outFIFO/n1181 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[80][3] ) );
  DF3 \u_outFIFO/FIFO_reg[81][0]  ( .D(\u_outFIFO/n1182 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[81][0] ) );
  DF3 \u_outFIFO/FIFO_reg[81][1]  ( .D(\u_outFIFO/n1183 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[81][1] ) );
  DF3 \u_outFIFO/FIFO_reg[81][2]  ( .D(\u_outFIFO/n1184 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[81][2] ) );
  DF3 \u_outFIFO/FIFO_reg[81][3]  ( .D(\u_outFIFO/n1185 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[81][3] ) );
  DF3 \u_outFIFO/FIFO_reg[82][0]  ( .D(\u_outFIFO/n1186 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[82][0] ) );
  DF3 \u_outFIFO/FIFO_reg[82][1]  ( .D(\u_outFIFO/n1187 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[82][1] ) );
  DF3 \u_outFIFO/FIFO_reg[82][2]  ( .D(\u_outFIFO/n1188 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[82][2] ) );
  DF3 \u_outFIFO/FIFO_reg[82][3]  ( .D(\u_outFIFO/n1189 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[82][3] ) );
  DF3 \u_outFIFO/FIFO_reg[83][0]  ( .D(\u_outFIFO/n1190 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[83][0] ) );
  DF3 \u_outFIFO/FIFO_reg[83][1]  ( .D(\u_outFIFO/n1191 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[83][1] ) );
  DF3 \u_outFIFO/FIFO_reg[83][2]  ( .D(\u_outFIFO/n1192 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[83][2] ) );
  DF3 \u_outFIFO/FIFO_reg[83][3]  ( .D(\u_outFIFO/n1193 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[83][3] ) );
  DF3 \u_outFIFO/FIFO_reg[84][0]  ( .D(\u_outFIFO/n1194 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[84][0] ) );
  DF3 \u_outFIFO/FIFO_reg[84][1]  ( .D(\u_outFIFO/n1195 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[84][1] ) );
  DF3 \u_outFIFO/FIFO_reg[84][2]  ( .D(\u_outFIFO/n1196 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[84][2] ) );
  DF3 \u_outFIFO/FIFO_reg[84][3]  ( .D(\u_outFIFO/n1197 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[84][3] ) );
  DF3 \u_outFIFO/FIFO_reg[85][0]  ( .D(\u_outFIFO/n1198 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[85][0] ) );
  DF3 \u_outFIFO/FIFO_reg[85][1]  ( .D(\u_outFIFO/n1199 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[85][1] ) );
  DF3 \u_outFIFO/FIFO_reg[85][2]  ( .D(\u_outFIFO/n1200 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[85][2] ) );
  DF3 \u_outFIFO/FIFO_reg[85][3]  ( .D(\u_outFIFO/n1201 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[85][3] ) );
  DF3 \u_outFIFO/FIFO_reg[86][0]  ( .D(\u_outFIFO/n1202 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[86][0] ) );
  DF3 \u_outFIFO/FIFO_reg[86][1]  ( .D(\u_outFIFO/n1203 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[86][1] ) );
  DF3 \u_outFIFO/FIFO_reg[86][2]  ( .D(\u_outFIFO/n1204 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[86][2] ) );
  DF3 \u_outFIFO/FIFO_reg[86][3]  ( .D(\u_outFIFO/n1205 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[86][3] ) );
  DF3 \u_outFIFO/FIFO_reg[87][0]  ( .D(\u_outFIFO/n1206 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[87][0] ) );
  DF3 \u_outFIFO/FIFO_reg[87][1]  ( .D(\u_outFIFO/n1207 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[87][1] ) );
  DF3 \u_outFIFO/FIFO_reg[87][2]  ( .D(\u_outFIFO/n1208 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[87][2] ) );
  DF3 \u_outFIFO/FIFO_reg[87][3]  ( .D(\u_outFIFO/n1209 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[87][3] ) );
  DF3 \u_outFIFO/FIFO_reg[88][0]  ( .D(\u_outFIFO/n1210 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[88][0] ) );
  DF3 \u_outFIFO/FIFO_reg[88][1]  ( .D(\u_outFIFO/n1211 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[88][1] ) );
  DF3 \u_outFIFO/FIFO_reg[88][2]  ( .D(\u_outFIFO/n1212 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[88][2] ) );
  DF3 \u_outFIFO/FIFO_reg[88][3]  ( .D(\u_outFIFO/n1213 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[88][3] ) );
  DF3 \u_outFIFO/FIFO_reg[89][0]  ( .D(\u_outFIFO/n1214 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[89][0] ) );
  DF3 \u_outFIFO/FIFO_reg[89][1]  ( .D(\u_outFIFO/n1215 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[89][1] ) );
  DF3 \u_outFIFO/FIFO_reg[89][2]  ( .D(\u_outFIFO/n1216 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[89][2] ) );
  DF3 \u_outFIFO/FIFO_reg[89][3]  ( .D(\u_outFIFO/n1217 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[89][3] ) );
  DF3 \u_outFIFO/FIFO_reg[90][0]  ( .D(\u_outFIFO/n1218 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[90][0] ) );
  DF3 \u_outFIFO/FIFO_reg[90][1]  ( .D(\u_outFIFO/n1219 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[90][1] ) );
  DF3 \u_outFIFO/FIFO_reg[90][2]  ( .D(\u_outFIFO/n1220 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[90][2] ) );
  DF3 \u_outFIFO/FIFO_reg[90][3]  ( .D(\u_outFIFO/n1221 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[90][3] ) );
  DF3 \u_outFIFO/FIFO_reg[91][0]  ( .D(\u_outFIFO/n1222 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[91][0] ) );
  DF3 \u_outFIFO/FIFO_reg[91][1]  ( .D(\u_outFIFO/n1223 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[91][1] ) );
  DF3 \u_outFIFO/FIFO_reg[91][2]  ( .D(\u_outFIFO/n1224 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[91][2] ) );
  DF3 \u_outFIFO/FIFO_reg[91][3]  ( .D(\u_outFIFO/n1225 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[91][3] ) );
  DF3 \u_outFIFO/FIFO_reg[92][0]  ( .D(\u_outFIFO/n1226 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[92][0] ) );
  DF3 \u_outFIFO/FIFO_reg[92][1]  ( .D(\u_outFIFO/n1227 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[92][1] ) );
  DF3 \u_outFIFO/FIFO_reg[92][2]  ( .D(\u_outFIFO/n1228 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[92][2] ) );
  DF3 \u_outFIFO/FIFO_reg[92][3]  ( .D(\u_outFIFO/n1229 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[92][3] ) );
  DF3 \u_outFIFO/FIFO_reg[93][0]  ( .D(\u_outFIFO/n1230 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[93][0] ) );
  DF3 \u_outFIFO/FIFO_reg[93][1]  ( .D(\u_outFIFO/n1231 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[93][1] ) );
  DF3 \u_outFIFO/FIFO_reg[93][2]  ( .D(\u_outFIFO/n1232 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[93][2] ) );
  DF3 \u_outFIFO/FIFO_reg[93][3]  ( .D(\u_outFIFO/n1233 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[93][3] ) );
  DF3 \u_outFIFO/FIFO_reg[94][0]  ( .D(\u_outFIFO/n1234 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[94][0] ) );
  DF3 \u_outFIFO/FIFO_reg[94][1]  ( .D(\u_outFIFO/n1235 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[94][1] ) );
  DF3 \u_outFIFO/FIFO_reg[94][2]  ( .D(\u_outFIFO/n1236 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[94][2] ) );
  DF3 \u_outFIFO/FIFO_reg[94][3]  ( .D(\u_outFIFO/n1237 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[94][3] ) );
  DF3 \u_outFIFO/FIFO_reg[95][0]  ( .D(\u_outFIFO/n1238 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[95][0] ) );
  DF3 \u_outFIFO/FIFO_reg[95][1]  ( .D(\u_outFIFO/n1239 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[95][1] ) );
  DF3 \u_outFIFO/FIFO_reg[95][2]  ( .D(\u_outFIFO/n1240 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[95][2] ) );
  DF3 \u_outFIFO/FIFO_reg[95][3]  ( .D(\u_outFIFO/n1241 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[95][3] ) );
  DF3 \u_outFIFO/FIFO_reg[96][0]  ( .D(\u_outFIFO/n1242 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[96][0] ) );
  DF3 \u_outFIFO/FIFO_reg[96][1]  ( .D(\u_outFIFO/n1243 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[96][1] ) );
  DF3 \u_outFIFO/FIFO_reg[96][2]  ( .D(\u_outFIFO/n1244 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[96][2] ) );
  DF3 \u_outFIFO/FIFO_reg[96][3]  ( .D(\u_outFIFO/n1245 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[96][3] ) );
  DF3 \u_outFIFO/FIFO_reg[97][0]  ( .D(\u_outFIFO/n1246 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[97][0] ) );
  DF3 \u_outFIFO/FIFO_reg[97][1]  ( .D(\u_outFIFO/n1247 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[97][1] ) );
  DF3 \u_outFIFO/FIFO_reg[97][2]  ( .D(\u_outFIFO/n1248 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[97][2] ) );
  DF3 \u_outFIFO/FIFO_reg[97][3]  ( .D(\u_outFIFO/n1249 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[97][3] ) );
  DF3 \u_outFIFO/FIFO_reg[98][0]  ( .D(\u_outFIFO/n1250 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[98][0] ) );
  DF3 \u_outFIFO/FIFO_reg[98][1]  ( .D(\u_outFIFO/n1251 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[98][1] ) );
  DF3 \u_outFIFO/FIFO_reg[98][2]  ( .D(\u_outFIFO/n1252 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[98][2] ) );
  DF3 \u_outFIFO/FIFO_reg[98][3]  ( .D(\u_outFIFO/n1253 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[98][3] ) );
  DF3 \u_outFIFO/FIFO_reg[99][0]  ( .D(\u_outFIFO/n1254 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[99][0] ) );
  DF3 \u_outFIFO/FIFO_reg[99][1]  ( .D(\u_outFIFO/n1255 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[99][1] ) );
  DF3 \u_outFIFO/FIFO_reg[99][2]  ( .D(\u_outFIFO/n1256 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[99][2] ) );
  DF3 \u_outFIFO/FIFO_reg[99][3]  ( .D(\u_outFIFO/n1257 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[99][3] ) );
  DF3 \u_outFIFO/FIFO_reg[100][0]  ( .D(\u_outFIFO/n1258 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[100][0] ) );
  DF3 \u_outFIFO/FIFO_reg[100][1]  ( .D(\u_outFIFO/n1259 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[100][1] ) );
  DF3 \u_outFIFO/FIFO_reg[100][2]  ( .D(\u_outFIFO/n1260 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[100][2] ) );
  DF3 \u_outFIFO/FIFO_reg[100][3]  ( .D(\u_outFIFO/n1261 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[100][3] ) );
  DF3 \u_outFIFO/FIFO_reg[101][0]  ( .D(\u_outFIFO/n1262 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[101][0] ) );
  DF3 \u_outFIFO/FIFO_reg[101][1]  ( .D(\u_outFIFO/n1263 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[101][1] ) );
  DF3 \u_outFIFO/FIFO_reg[101][2]  ( .D(\u_outFIFO/n1264 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[101][2] ) );
  DF3 \u_outFIFO/FIFO_reg[101][3]  ( .D(\u_outFIFO/n1265 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[101][3] ) );
  DF3 \u_outFIFO/FIFO_reg[102][0]  ( .D(\u_outFIFO/n1266 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[102][0] ) );
  DF3 \u_outFIFO/FIFO_reg[102][1]  ( .D(\u_outFIFO/n1267 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[102][1] ) );
  DF3 \u_outFIFO/FIFO_reg[102][2]  ( .D(\u_outFIFO/n1268 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[102][2] ) );
  DF3 \u_outFIFO/FIFO_reg[102][3]  ( .D(\u_outFIFO/n1269 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[102][3] ) );
  DF3 \u_outFIFO/FIFO_reg[103][0]  ( .D(\u_outFIFO/n1270 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[103][0] ) );
  DF3 \u_outFIFO/FIFO_reg[103][1]  ( .D(\u_outFIFO/n1271 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[103][1] ) );
  DF3 \u_outFIFO/FIFO_reg[103][2]  ( .D(\u_outFIFO/n1272 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[103][2] ) );
  DF3 \u_outFIFO/FIFO_reg[103][3]  ( .D(\u_outFIFO/n1273 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[103][3] ) );
  DF3 \u_outFIFO/FIFO_reg[104][0]  ( .D(\u_outFIFO/n1274 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[104][0] ) );
  DF3 \u_outFIFO/FIFO_reg[104][1]  ( .D(\u_outFIFO/n1275 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[104][1] ) );
  DF3 \u_outFIFO/FIFO_reg[104][2]  ( .D(\u_outFIFO/n1276 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[104][2] ) );
  DF3 \u_outFIFO/FIFO_reg[104][3]  ( .D(\u_outFIFO/n1277 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[104][3] ) );
  DF3 \u_outFIFO/FIFO_reg[105][0]  ( .D(\u_outFIFO/n1278 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[105][0] ) );
  DF3 \u_outFIFO/FIFO_reg[105][1]  ( .D(\u_outFIFO/n1279 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[105][1] ) );
  DF3 \u_outFIFO/FIFO_reg[105][2]  ( .D(\u_outFIFO/n1280 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[105][2] ) );
  DF3 \u_outFIFO/FIFO_reg[105][3]  ( .D(\u_outFIFO/n1281 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[105][3] ) );
  DF3 \u_outFIFO/FIFO_reg[106][0]  ( .D(\u_outFIFO/n1282 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[106][0] ) );
  DF3 \u_outFIFO/FIFO_reg[106][1]  ( .D(\u_outFIFO/n1283 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[106][1] ) );
  DF3 \u_outFIFO/FIFO_reg[106][2]  ( .D(\u_outFIFO/n1284 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[106][2] ) );
  DF3 \u_outFIFO/FIFO_reg[106][3]  ( .D(\u_outFIFO/n1285 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[106][3] ) );
  DF3 \u_outFIFO/FIFO_reg[107][0]  ( .D(\u_outFIFO/n1286 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[107][0] ) );
  DF3 \u_outFIFO/FIFO_reg[107][1]  ( .D(\u_outFIFO/n1287 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[107][1] ) );
  DF3 \u_outFIFO/FIFO_reg[107][2]  ( .D(\u_outFIFO/n1288 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[107][2] ) );
  DF3 \u_outFIFO/FIFO_reg[107][3]  ( .D(\u_outFIFO/n1289 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[107][3] ) );
  DF3 \u_outFIFO/FIFO_reg[108][0]  ( .D(\u_outFIFO/n1290 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[108][0] ) );
  DF3 \u_outFIFO/FIFO_reg[108][1]  ( .D(\u_outFIFO/n1291 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[108][1] ) );
  DF3 \u_outFIFO/FIFO_reg[108][2]  ( .D(\u_outFIFO/n1292 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[108][2] ) );
  DF3 \u_outFIFO/FIFO_reg[108][3]  ( .D(\u_outFIFO/n1293 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[108][3] ) );
  DF3 \u_outFIFO/FIFO_reg[109][0]  ( .D(\u_outFIFO/n1294 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[109][0] ) );
  DF3 \u_outFIFO/FIFO_reg[109][1]  ( .D(\u_outFIFO/n1295 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[109][1] ) );
  DF3 \u_outFIFO/FIFO_reg[109][2]  ( .D(\u_outFIFO/n1296 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[109][2] ) );
  DF3 \u_outFIFO/FIFO_reg[109][3]  ( .D(\u_outFIFO/n1297 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[109][3] ) );
  DF3 \u_outFIFO/FIFO_reg[110][0]  ( .D(\u_outFIFO/n1298 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[110][0] ) );
  DF3 \u_outFIFO/FIFO_reg[110][1]  ( .D(\u_outFIFO/n1299 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[110][1] ) );
  DF3 \u_outFIFO/FIFO_reg[110][2]  ( .D(\u_outFIFO/n1300 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[110][2] ) );
  DF3 \u_outFIFO/FIFO_reg[110][3]  ( .D(\u_outFIFO/n1301 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[110][3] ) );
  DF3 \u_outFIFO/FIFO_reg[111][0]  ( .D(\u_outFIFO/n1302 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[111][0] ) );
  DF3 \u_outFIFO/FIFO_reg[111][1]  ( .D(\u_outFIFO/n1303 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[111][1] ) );
  DF3 \u_outFIFO/FIFO_reg[111][2]  ( .D(\u_outFIFO/n1304 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[111][2] ) );
  DF3 \u_outFIFO/FIFO_reg[111][3]  ( .D(\u_outFIFO/n1305 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[111][3] ) );
  DF3 \u_outFIFO/FIFO_reg[112][0]  ( .D(\u_outFIFO/n1306 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[112][0] ) );
  DF3 \u_outFIFO/FIFO_reg[112][1]  ( .D(\u_outFIFO/n1307 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[112][1] ) );
  DF3 \u_outFIFO/FIFO_reg[112][2]  ( .D(\u_outFIFO/n1308 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[112][2] ) );
  DF3 \u_outFIFO/FIFO_reg[112][3]  ( .D(\u_outFIFO/n1309 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[112][3] ) );
  DF3 \u_outFIFO/FIFO_reg[113][0]  ( .D(\u_outFIFO/n1310 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[113][0] ) );
  DF3 \u_outFIFO/FIFO_reg[113][1]  ( .D(\u_outFIFO/n1311 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[113][1] ) );
  DF3 \u_outFIFO/FIFO_reg[113][2]  ( .D(\u_outFIFO/n1312 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[113][2] ) );
  DF3 \u_outFIFO/FIFO_reg[113][3]  ( .D(\u_outFIFO/n1313 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[113][3] ) );
  DF3 \u_outFIFO/FIFO_reg[114][0]  ( .D(\u_outFIFO/n1314 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[114][0] ) );
  DF3 \u_outFIFO/FIFO_reg[114][1]  ( .D(\u_outFIFO/n1315 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[114][1] ) );
  DF3 \u_outFIFO/FIFO_reg[114][2]  ( .D(\u_outFIFO/n1316 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[114][2] ) );
  DF3 \u_outFIFO/FIFO_reg[114][3]  ( .D(\u_outFIFO/n1317 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[114][3] ) );
  DF3 \u_outFIFO/FIFO_reg[115][0]  ( .D(\u_outFIFO/n1318 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[115][0] ) );
  DF3 \u_outFIFO/FIFO_reg[115][1]  ( .D(\u_outFIFO/n1319 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[115][1] ) );
  DF3 \u_outFIFO/FIFO_reg[115][2]  ( .D(\u_outFIFO/n1320 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[115][2] ) );
  DF3 \u_outFIFO/FIFO_reg[115][3]  ( .D(\u_outFIFO/n1321 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[115][3] ) );
  DF3 \u_outFIFO/FIFO_reg[116][0]  ( .D(\u_outFIFO/n1322 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[116][0] ) );
  DF3 \u_outFIFO/FIFO_reg[116][1]  ( .D(\u_outFIFO/n1323 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[116][1] ) );
  DF3 \u_outFIFO/FIFO_reg[116][2]  ( .D(\u_outFIFO/n1324 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[116][2] ) );
  DF3 \u_outFIFO/FIFO_reg[116][3]  ( .D(\u_outFIFO/n1325 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[116][3] ) );
  DF3 \u_outFIFO/FIFO_reg[117][0]  ( .D(\u_outFIFO/n1326 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[117][0] ) );
  DF3 \u_outFIFO/FIFO_reg[117][1]  ( .D(\u_outFIFO/n1327 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[117][1] ) );
  DF3 \u_outFIFO/FIFO_reg[117][2]  ( .D(\u_outFIFO/n1328 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[117][2] ) );
  DF3 \u_outFIFO/FIFO_reg[117][3]  ( .D(\u_outFIFO/n1329 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[117][3] ) );
  DF3 \u_outFIFO/FIFO_reg[118][0]  ( .D(\u_outFIFO/n1330 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[118][0] ) );
  DF3 \u_outFIFO/FIFO_reg[118][1]  ( .D(\u_outFIFO/n1331 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[118][1] ) );
  DF3 \u_outFIFO/FIFO_reg[118][2]  ( .D(\u_outFIFO/n1332 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[118][2] ) );
  DF3 \u_outFIFO/FIFO_reg[118][3]  ( .D(\u_outFIFO/n1333 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[118][3] ) );
  DF3 \u_outFIFO/FIFO_reg[119][0]  ( .D(\u_outFIFO/n1334 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[119][0] ) );
  DF3 \u_outFIFO/FIFO_reg[119][1]  ( .D(\u_outFIFO/n1335 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[119][1] ) );
  DF3 \u_outFIFO/FIFO_reg[119][2]  ( .D(\u_outFIFO/n1336 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[119][2] ) );
  DF3 \u_outFIFO/FIFO_reg[119][3]  ( .D(\u_outFIFO/n1337 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[119][3] ) );
  DF3 \u_outFIFO/FIFO_reg[120][0]  ( .D(\u_outFIFO/n1338 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[120][0] ) );
  DF3 \u_outFIFO/FIFO_reg[120][1]  ( .D(\u_outFIFO/n1339 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[120][1] ) );
  DF3 \u_outFIFO/FIFO_reg[120][2]  ( .D(\u_outFIFO/n1340 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[120][2] ) );
  DF3 \u_outFIFO/FIFO_reg[120][3]  ( .D(\u_outFIFO/n1341 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[120][3] ) );
  DF3 \u_outFIFO/FIFO_reg[121][0]  ( .D(\u_outFIFO/n1342 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[121][0] ) );
  DF3 \u_outFIFO/FIFO_reg[121][1]  ( .D(\u_outFIFO/n1343 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[121][1] ) );
  DF3 \u_outFIFO/FIFO_reg[121][2]  ( .D(\u_outFIFO/n1344 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[121][2] ) );
  DF3 \u_outFIFO/FIFO_reg[121][3]  ( .D(\u_outFIFO/n1345 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[121][3] ) );
  DF3 \u_outFIFO/FIFO_reg[122][0]  ( .D(\u_outFIFO/n1346 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[122][0] ) );
  DF3 \u_outFIFO/FIFO_reg[122][1]  ( .D(\u_outFIFO/n1347 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[122][1] ) );
  DF3 \u_outFIFO/FIFO_reg[122][2]  ( .D(\u_outFIFO/n1348 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[122][2] ) );
  DF3 \u_outFIFO/FIFO_reg[122][3]  ( .D(\u_outFIFO/n1349 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[122][3] ) );
  DF3 \u_outFIFO/FIFO_reg[123][0]  ( .D(\u_outFIFO/n1350 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[123][0] ) );
  DF3 \u_outFIFO/FIFO_reg[123][1]  ( .D(\u_outFIFO/n1351 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[123][1] ) );
  DF3 \u_outFIFO/FIFO_reg[123][2]  ( .D(\u_outFIFO/n1352 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[123][2] ) );
  DF3 \u_outFIFO/FIFO_reg[123][3]  ( .D(\u_outFIFO/n1353 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[123][3] ) );
  DF3 \u_outFIFO/FIFO_reg[124][0]  ( .D(\u_outFIFO/n1354 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[124][0] ) );
  DF3 \u_outFIFO/FIFO_reg[124][1]  ( .D(\u_outFIFO/n1355 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[124][1] ) );
  DF3 \u_outFIFO/FIFO_reg[124][2]  ( .D(\u_outFIFO/n1356 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[124][2] ) );
  DF3 \u_outFIFO/FIFO_reg[124][3]  ( .D(\u_outFIFO/n1357 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[124][3] ) );
  DF3 \u_outFIFO/FIFO_reg[125][0]  ( .D(\u_outFIFO/n1358 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[125][0] ) );
  DF3 \u_outFIFO/FIFO_reg[125][1]  ( .D(\u_outFIFO/n1359 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[125][1] ) );
  DF3 \u_outFIFO/FIFO_reg[125][2]  ( .D(\u_outFIFO/n1360 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[125][2] ) );
  DF3 \u_outFIFO/FIFO_reg[125][3]  ( .D(\u_outFIFO/n1361 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[125][3] ) );
  DF3 \u_outFIFO/FIFO_reg[126][0]  ( .D(\u_outFIFO/n1362 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[126][0] ) );
  DF3 \u_outFIFO/FIFO_reg[126][1]  ( .D(\u_outFIFO/n1363 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[126][1] ) );
  DF3 \u_outFIFO/FIFO_reg[126][2]  ( .D(\u_outFIFO/n1364 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[126][2] ) );
  DF3 \u_outFIFO/FIFO_reg[126][3]  ( .D(\u_outFIFO/n1365 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[126][3] ) );
  DF3 \u_outFIFO/FIFO_reg[127][0]  ( .D(\u_outFIFO/n1366 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[127][0] ) );
  DF3 \u_outFIFO/FIFO_reg[127][1]  ( .D(\u_outFIFO/n1367 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[127][1] ) );
  DF3 \u_outFIFO/FIFO_reg[127][2]  ( .D(\u_outFIFO/n1368 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[127][2] ) );
  DF3 \u_outFIFO/FIFO_reg[127][3]  ( .D(\u_outFIFO/n1369 ), .C(inClock), .Q(
        \u_outFIFO/FIFO[127][3] ) );
  DF3 \u_outFIFO/j_FIFO_reg[6]  ( .D(\u_outFIFO/n1370 ), .C(inClock), .Q(
        \u_outFIFO/N45 ), .QN(\u_outFIFO/n295 ) );
  DF3 \u_outFIFO/j_FIFO_reg[5]  ( .D(\u_outFIFO/n1371 ), .C(inClock), .Q(
        \u_outFIFO/N44 ), .QN(\u_outFIFO/n296 ) );
  DF3 \u_outFIFO/j_FIFO_reg[4]  ( .D(\u_outFIFO/n1372 ), .C(inClock), .Q(
        \u_outFIFO/N43 ), .QN(\u_outFIFO/n297 ) );
  DF3 \u_outFIFO/j_FIFO_reg[3]  ( .D(\u_outFIFO/n1373 ), .C(inClock), .Q(
        \u_outFIFO/N42 ), .QN(\u_outFIFO/n298 ) );
  DF3 \u_outFIFO/j_FIFO_reg[2]  ( .D(\u_outFIFO/n1374 ), .C(inClock), .Q(n14), 
        .QN(\u_outFIFO/n299 ) );
  DF3 \u_outFIFO/j_FIFO_reg[1]  ( .D(\u_outFIFO/n1375 ), .C(inClock), .Q(
        \u_outFIFO/N40 ), .QN(\u_outFIFO/n300 ) );
  DF3 \u_outFIFO/j_FIFO_reg[0]  ( .D(\u_outFIFO/n1376 ), .C(inClock), .Q(
        \u_outFIFO/N39 ), .QN(\u_outFIFO/n301 ) );
  DF3 \u_outFIFO/currentState_reg[3]  ( .D(\u_outFIFO/N50 ), .C(inClock), .QN(
        \u_outFIFO/n253 ) );
  DF3 \u_outFIFO/currentState_reg[1]  ( .D(\u_outFIFO/N48 ), .C(inClock), .Q(
        \u_outFIFO/currentState [1]), .QN(\u_outFIFO/n256 ) );
  DF3 \u_outFIFO/sigRDCOUNT_reg[6]  ( .D(n1804), .C(inClock), .Q(
        \u_outFIFO/outReadCount[6] ), .QN(n218) );
  DF3 \u_outFIFO/sigRDCOUNT_reg[5]  ( .D(n1803), .C(inClock), .Q(
        \u_outFIFO/outReadCount[5] ), .QN(n220) );
  DF3 \u_outFIFO/sigRDCOUNT_reg[4]  ( .D(n1802), .C(inClock), .Q(
        \u_outFIFO/outReadCount[4] ), .QN(n196) );
  DF3 \u_outFIFO/sigRDCOUNT_reg[3]  ( .D(n1801), .C(inClock), .Q(
        \u_outFIFO/outReadCount[3] ), .QN(n169) );
  DF3 \u_outFIFO/sigRDCOUNT_reg[2]  ( .D(n1800), .C(inClock), .Q(
        \u_outFIFO/outReadCount[2] ), .QN(n167) );
  DF3 \u_outFIFO/sigRDCOUNT_reg[1]  ( .D(n1799), .C(inClock), .Q(
        \u_outFIFO/outReadCount[1] ), .QN(n161) );
  DF3 \u_outFIFO/sigRDCOUNT_reg[0]  ( .D(n1798), .C(inClock), .Q(
        \u_outFIFO/outReadCount[0] ), .QN(n130) );
  DF3 \u_outFIFO/currentState_reg[0]  ( .D(\u_outFIFO/N47 ), .C(inClock), .Q(
        \u_outFIFO/currentState [0]), .QN(\u_outFIFO/n257 ) );
  DF3 \u_outFIFO/k_FIFO_reg[1]  ( .D(\u_outFIFO/n1377 ), .C(inClock), .Q(
        \u_outFIFO/k_FIFO [1]), .QN(\u_outFIFO/n284 ) );
  JK3 \u_outFIFO/k_FIFO_reg[0]  ( .J(n926), .K(n1191), .C(inClock), .Q(
        \u_outFIFO/k_FIFO [0]), .QN(\u_outFIFO/n285 ) );
  DF3 \u_outFIFO/currentState_reg[2]  ( .D(\u_outFIFO/N49 ), .C(inClock), .Q(
        \u_outFIFO/currentState [2]), .QN(\u_outFIFO/n254 ) );
  DF3 \u_outFIFO/sigWRCOUNT_reg[5]  ( .D(\u_outFIFO/n1379 ), .C(inClock), .Q(
        \u_outFIFO/outWriteCount[5] ), .QN(\u_outFIFO/n261 ) );
  DF3 \u_outFIFO/sigWRCOUNT_reg[4]  ( .D(\u_outFIFO/n1380 ), .C(inClock), .Q(
        \u_outFIFO/outWriteCount[4] ), .QN(\u_outFIFO/n262 ) );
  DF3 \u_outFIFO/sigWRCOUNT_reg[3]  ( .D(\u_outFIFO/n1381 ), .C(inClock), .Q(
        \u_outFIFO/outWriteCount[3] ), .QN(\u_outFIFO/n263 ) );
  DF3 \u_outFIFO/sigWRCOUNT_reg[2]  ( .D(\u_outFIFO/n1382 ), .C(inClock), .Q(
        \u_outFIFO/outWriteCount[2] ), .QN(\u_outFIFO/n264 ) );
  DF3 \u_outFIFO/sigWRCOUNT_reg[1]  ( .D(\u_outFIFO/n1383 ), .C(inClock), .Q(
        \u_outFIFO/outWriteCount[1] ), .QN(\u_outFIFO/n265 ) );
  DF3 \u_outFIFO/sigWRCOUNT_reg[0]  ( .D(\u_outFIFO/n1384 ), .C(inClock), .Q(
        \u_outFIFO/outWriteCount[0] ), .QN(\u_outFIFO/n266 ) );
  DF3 \u_outFIFO/sigWRCOUNT_reg[6]  ( .D(\u_outFIFO/n1378 ), .C(inClock), .Q(
        \u_outFIFO/outWriteCount[6] ), .QN(\u_outFIFO/n260 ) );
  DF3 \u_outFIFO/sigWRCOUNT_reg[7]  ( .D(\u_outFIFO/n1385 ), .C(inClock), .Q(
        \u_outFIFO/outWriteCount[7] ), .QN(\u_outFIFO/n258 ) );
  DF3 \u_outFIFO/i_FIFO_reg[6]  ( .D(\u_outFIFO/n1386 ), .C(inClock), .Q(
        \u_outFIFO/i_FIFO [6]), .QN(\u_outFIFO/n267 ) );
  DF3 \u_outFIFO/i_FIFO_reg[5]  ( .D(\u_outFIFO/n1387 ), .C(inClock), .Q(
        \u_outFIFO/i_FIFO [5]), .QN(\u_outFIFO/n275 ) );
  DF3 \u_outFIFO/i_FIFO_reg[4]  ( .D(\u_outFIFO/n1388 ), .C(inClock), .Q(
        \u_outFIFO/i_FIFO [4]), .QN(\u_outFIFO/n276 ) );
  DF3 \u_outFIFO/i_FIFO_reg[3]  ( .D(\u_outFIFO/n1389 ), .C(inClock), .Q(
        \u_outFIFO/i_FIFO [3]), .QN(\u_outFIFO/n277 ) );
  DF3 \u_outFIFO/i_FIFO_reg[2]  ( .D(\u_outFIFO/n1390 ), .C(inClock), .Q(
        \u_outFIFO/i_FIFO [2]), .QN(\u_outFIFO/n278 ) );
  DF3 \u_outFIFO/i_FIFO_reg[1]  ( .D(\u_outFIFO/n1391 ), .C(inClock), .Q(
        \u_outFIFO/i_FIFO [1]), .QN(\u_outFIFO/n279 ) );
  DF3 \u_outFIFO/i_FIFO_reg[0]  ( .D(\u_outFIFO/n1392 ), .C(inClock), .Q(
        \u_outFIFO/i_FIFO [0]), .QN(\u_outFIFO/n280 ) );
  DF3 \u_outFIFO/sigEnableCounter_reg  ( .D(\u_outFIFO/N198 ), .C(inClock), 
        .Q(\u_outFIFO/sigEnableCounter ) );
  DF3 \u_decoder/iq_demod/o_I_prefilter_reg[0]  ( .D(n2274), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_0 [0]), .QN(n84) );
  DF3 \u_decoder/iq_demod/o_I_prefilter_reg[1]  ( .D(n2299), .C(inClock), .Q(
        n12), .QN(n74) );
  DF3 \u_decoder/iq_demod/o_I_prefilter_reg[2]  ( .D(n2301), .C(inClock), .Q(
        n4), .QN(n89) );
  DF3 \u_decoder/iq_demod/o_I_prefilter_reg[3]  ( .D(n2302), .C(inClock), .Q(
        n8), .QN(n80) );
  DF3 \u_decoder/iq_demod/o_I_prefilter_reg[4]  ( .D(n2303), .C(inClock), .Q(
        \u_decoder/I_prefilter [4]), .QN(n164) );
  DF3 \u_decoder/iq_demod/o_I_prefilter_reg[5]  ( .D(n2304), .C(inClock), .Q(
        n10), .QN(n16) );
  DF3 \u_decoder/iq_demod/o_I_prefilter_reg[6]  ( .D(n2306), .C(inClock), .Q(
        n6), .QN(n18) );
  DF3 \u_decoder/iq_demod/o_I_prefilter_reg[7]  ( .D(n2307), .C(inClock), .Q(
        \u_decoder/I_prefilter [7]), .QN(n194) );
  DF3 \u_decoder/iq_demod/o_Q_prefilter_reg[0]  ( .D(n2345), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_0 [0]), .QN(n88) );
  DF3 \u_decoder/iq_demod/o_Q_prefilter_reg[1]  ( .D(n2370), .C(inClock), .Q(
        n11), .QN(n75) );
  DF3 \u_decoder/iq_demod/o_Q_prefilter_reg[2]  ( .D(n2372), .C(inClock), .Q(
        n3), .QN(n90) );
  DF3 \u_decoder/iq_demod/o_Q_prefilter_reg[3]  ( .D(n2373), .C(inClock), .Q(
        n7), .QN(n81) );
  DF3 \u_decoder/iq_demod/o_Q_prefilter_reg[4]  ( .D(n2374), .C(inClock), .Q(
        \u_decoder/Q_prefilter [4]), .QN(n165) );
  DF3 \u_decoder/iq_demod/o_Q_prefilter_reg[5]  ( .D(n2375), .C(inClock), .Q(
        n9), .QN(n17) );
  DF3 \u_decoder/iq_demod/o_Q_prefilter_reg[6]  ( .D(n2377), .C(inClock), .Q(
        n5), .QN(n19) );
  DF3 \u_decoder/iq_demod/o_Q_prefilter_reg[7]  ( .D(n2378), .C(inClock), .Q(
        \u_decoder/Q_prefilter [7]), .QN(n195) );
  DF3 \u_decoder/iq_demod/o_sample_ready_reg  ( .D(n2379), .C(inClock), .Q(
        \u_decoder/sample_ready ), .QN(n294) );
  DF3 \u_decoder/iq_demod/Q_if_buff_reg[0]  ( .D(n1580), .C(inClock), .Q(
        \u_decoder/iq_demod/Q_if_signed [0]), .QN(n123) );
  DF3 \u_decoder/iq_demod/Q_if_buff_reg[1]  ( .D(n1579), .C(inClock), .Q(
        \u_decoder/iq_demod/Q_if_signed [1]), .QN(n120) );
  DF3 \u_decoder/iq_demod/Q_if_buff_reg[2]  ( .D(n1578), .C(inClock), .Q(
        \u_decoder/iq_demod/Q_if_signed [2]), .QN(n124) );
  DF3 \u_decoder/iq_demod/Q_if_buff_reg[3]  ( .D(n1577), .C(inClock), .Q(
        \u_decoder/iq_demod/Q_if_buff[3] ), .QN(
        \u_decoder/iq_demod/Q_if_signed [3]) );
  DF3 \u_decoder/iq_demod/I_if_buff_reg[0]  ( .D(n1576), .C(inClock), .Q(
        \u_decoder/iq_demod/I_if_signed [0]), .QN(n122) );
  DF3 \u_decoder/iq_demod/I_if_buff_reg[1]  ( .D(n1575), .C(inClock), .Q(
        \u_decoder/iq_demod/I_if_signed [1]), .QN(n121) );
  DF3 \u_decoder/iq_demod/I_if_buff_reg[2]  ( .D(n1574), .C(inClock), .Q(
        \u_decoder/iq_demod/I_if_signed [2]), .QN(n125) );
  DF3 \u_decoder/iq_demod/I_if_buff_reg[3]  ( .D(n1573), .C(inClock), .Q(
        \u_decoder/iq_demod/I_if_buff[3] ), .QN(
        \u_decoder/iq_demod/I_if_signed [3]) );
  DF3 \u_decoder/iq_demod/state_reg[1]  ( .D(n1909), .C(inClock), .Q(
        \u_decoder/iq_demod/state [1]) );
  DF3 \u_decoder/iq_demod/state_reg[0]  ( .D(\u_decoder/iq_demod/N13 ), .C(
        inClock), .Q(\u_decoder/iq_demod/state [0]), .QN(
        \u_decoder/iq_demod/n30 ) );
  DF3 \u_decoder/fir_filter/o_Q_postfilter_reg[3]  ( .D(n2399), .C(inClock), 
        .Q(sig_decod_outQ[3]) );
  DF3 \u_decoder/fir_filter/o_Q_postfilter_reg[2]  ( .D(n2400), .C(inClock), 
        .Q(sig_decod_outQ[2]) );
  DF3 \u_decoder/fir_filter/o_Q_postfilter_reg[1]  ( .D(n2401), .C(inClock), 
        .Q(sig_decod_outQ[1]) );
  DF3 \u_decoder/fir_filter/o_Q_postfilter_reg[0]  ( .D(n2402), .C(inClock), 
        .Q(sig_decod_outQ[0]) );
  DF3 \u_decoder/fir_filter/Q_data_add_1_buff_reg[14]  ( .D(n2403), .C(inClock), .Q(\u_decoder/fir_filter/Q_data_add_1_buff [14]) );
  DF3 \u_decoder/fir_filter/Q_data_add_1_buff_reg[13]  ( .D(n2404), .C(inClock), .Q(\u_decoder/fir_filter/Q_data_add_1_buff [13]) );
  DF3 \u_decoder/fir_filter/Q_data_add_1_buff_reg[12]  ( .D(n2405), .C(inClock), .Q(\u_decoder/fir_filter/Q_data_add_1_buff [12]) );
  DF3 \u_decoder/fir_filter/Q_data_add_1_buff_reg[11]  ( .D(n2406), .C(inClock), .Q(\u_decoder/fir_filter/Q_data_add_1_buff [11]) );
  DF3 \u_decoder/fir_filter/Q_data_add_1_buff_reg[10]  ( .D(n2407), .C(inClock), .Q(\u_decoder/fir_filter/Q_data_add_1_buff [10]) );
  DF3 \u_decoder/fir_filter/Q_data_add_1_buff_reg[9]  ( .D(n2410), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_1_buff [9]) );
  DF3 \u_decoder/fir_filter/Q_data_add_1_buff_reg[8]  ( .D(n2411), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_1_buff [8]) );
  DF3 \u_decoder/fir_filter/Q_data_add_1_buff_reg[7]  ( .D(n2414), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_1_buff [7]) );
  DF3 \u_decoder/fir_filter/Q_data_add_1_buff_reg[6]  ( .D(n2415), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_1_buff [6]) );
  DF3 \u_decoder/fir_filter/Q_data_add_1_buff_reg[5]  ( .D(n2417), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_1_buff [5]) );
  DF3 \u_decoder/fir_filter/Q_data_add_1_buff_reg[4]  ( .D(n2419), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_1_buff [4]) );
  DF3 \u_decoder/fir_filter/Q_data_add_1_buff_reg[3]  ( .D(n2421), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_1_buff [3]) );
  DF3 \u_decoder/fir_filter/Q_data_add_1_buff_reg[2]  ( .D(n2423), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_1_buff [2]) );
  DF3 \u_decoder/fir_filter/Q_data_add_1_buff_reg[1]  ( .D(n2425), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_1_buff [1]), .QN(n24) );
  DF3 \u_decoder/fir_filter/Q_data_add_1_buff_reg[0]  ( .D(n2426), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_1_buff [0]) );
  DF3 \u_decoder/fir_filter/Q_data_add_2_buff_reg[14]  ( .D(n2427), .C(inClock), .Q(\u_decoder/fir_filter/Q_data_add_2_buff [14]) );
  DF3 \u_decoder/fir_filter/Q_data_add_2_buff_reg[13]  ( .D(n2428), .C(inClock), .Q(\u_decoder/fir_filter/Q_data_add_2_buff [13]) );
  DF3 \u_decoder/fir_filter/Q_data_add_2_buff_reg[12]  ( .D(n2429), .C(inClock), .Q(\u_decoder/fir_filter/Q_data_add_2_buff [12]) );
  DF3 \u_decoder/fir_filter/Q_data_add_2_buff_reg[11]  ( .D(n2430), .C(inClock), .Q(\u_decoder/fir_filter/Q_data_add_2_buff [11]) );
  DF3 \u_decoder/fir_filter/Q_data_add_2_buff_reg[10]  ( .D(n2431), .C(inClock), .Q(\u_decoder/fir_filter/Q_data_add_2_buff [10]) );
  DF3 \u_decoder/fir_filter/Q_data_add_2_buff_reg[9]  ( .D(n2432), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_2_buff [9]) );
  DF3 \u_decoder/fir_filter/Q_data_add_2_buff_reg[8]  ( .D(n2433), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_2_buff [8]) );
  DF3 \u_decoder/fir_filter/Q_data_add_2_buff_reg[7]  ( .D(n2434), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_2_buff [7]) );
  DF3 \u_decoder/fir_filter/Q_data_add_2_buff_reg[6]  ( .D(n2435), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_2_buff [6]) );
  DF3 \u_decoder/fir_filter/Q_data_add_2_buff_reg[5]  ( .D(n2436), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_2_buff [5]) );
  DF3 \u_decoder/fir_filter/Q_data_add_2_buff_reg[4]  ( .D(n2437), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_2_buff [4]) );
  DF3 \u_decoder/fir_filter/Q_data_add_2_buff_reg[3]  ( .D(n2438), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_2_buff [3]) );
  DF3 \u_decoder/fir_filter/Q_data_add_2_buff_reg[2]  ( .D(n2439), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_2_buff [2]) );
  DF3 \u_decoder/fir_filter/Q_data_add_2_buff_reg[1]  ( .D(n2440), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_2_buff [1]) );
  DF3 \u_decoder/fir_filter/Q_data_add_2_buff_reg[0]  ( .D(n2441), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_2_buff [0]), .QN(n117) );
  DF3 \u_decoder/fir_filter/Q_data_add_3_buff_reg[14]  ( .D(n2442), .C(inClock), .Q(\u_decoder/fir_filter/Q_data_add_3_buff [14]) );
  DF3 \u_decoder/fir_filter/Q_data_add_3_buff_reg[13]  ( .D(n2443), .C(inClock), .Q(\u_decoder/fir_filter/Q_data_add_3_buff [13]) );
  DF3 \u_decoder/fir_filter/Q_data_add_3_buff_reg[12]  ( .D(n2444), .C(inClock), .Q(\u_decoder/fir_filter/Q_data_add_3_buff [12]) );
  DF3 \u_decoder/fir_filter/Q_data_add_3_buff_reg[11]  ( .D(n2445), .C(inClock), .Q(\u_decoder/fir_filter/Q_data_add_3_buff [11]) );
  DF3 \u_decoder/fir_filter/Q_data_add_3_buff_reg[10]  ( .D(n2446), .C(inClock), .Q(\u_decoder/fir_filter/Q_data_add_3_buff [10]) );
  DF3 \u_decoder/fir_filter/Q_data_add_3_buff_reg[9]  ( .D(n2447), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_3_buff [9]) );
  DF3 \u_decoder/fir_filter/Q_data_add_3_buff_reg[8]  ( .D(n2448), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_3_buff [8]) );
  DF3 \u_decoder/fir_filter/Q_data_add_3_buff_reg[7]  ( .D(n2449), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_3_buff [7]) );
  DF3 \u_decoder/fir_filter/Q_data_add_3_buff_reg[6]  ( .D(n2450), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_3_buff [6]) );
  DF3 \u_decoder/fir_filter/Q_data_add_3_buff_reg[5]  ( .D(n2451), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_3_buff [5]) );
  DF3 \u_decoder/fir_filter/Q_data_add_3_buff_reg[4]  ( .D(n2452), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_3_buff [4]) );
  DF3 \u_decoder/fir_filter/Q_data_add_3_buff_reg[3]  ( .D(n2453), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_3_buff [3]) );
  DF3 \u_decoder/fir_filter/Q_data_add_3_buff_reg[2]  ( .D(n2454), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_3_buff [2]) );
  DF3 \u_decoder/fir_filter/Q_data_add_3_buff_reg[1]  ( .D(n2455), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_3_buff [1]) );
  DF3 \u_decoder/fir_filter/Q_data_add_3_buff_reg[0]  ( .D(n2456), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_3_buff [0]), .QN(n116) );
  DF3 \u_decoder/fir_filter/Q_data_add_4_buff_reg[14]  ( .D(n2457), .C(inClock), .Q(\u_decoder/fir_filter/Q_data_add_4_buff [14]) );
  DF3 \u_decoder/fir_filter/Q_data_add_4_buff_reg[13]  ( .D(n2458), .C(inClock), .Q(\u_decoder/fir_filter/Q_data_add_4_buff [13]) );
  DF3 \u_decoder/fir_filter/Q_data_add_4_buff_reg[12]  ( .D(n2459), .C(inClock), .Q(\u_decoder/fir_filter/Q_data_add_4_buff [12]) );
  DF3 \u_decoder/fir_filter/Q_data_add_4_buff_reg[11]  ( .D(n2460), .C(inClock), .Q(\u_decoder/fir_filter/Q_data_add_4_buff [11]) );
  DF3 \u_decoder/fir_filter/Q_data_add_4_buff_reg[10]  ( .D(n2461), .C(inClock), .Q(\u_decoder/fir_filter/Q_data_add_4_buff [10]) );
  DF3 \u_decoder/fir_filter/Q_data_add_4_buff_reg[9]  ( .D(n2462), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_4_buff [9]) );
  DF3 \u_decoder/fir_filter/Q_data_add_4_buff_reg[8]  ( .D(n2463), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_4_buff [8]) );
  DF3 \u_decoder/fir_filter/Q_data_add_4_buff_reg[7]  ( .D(n2464), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_4_buff [7]) );
  DF3 \u_decoder/fir_filter/Q_data_add_4_buff_reg[6]  ( .D(n2465), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_4_buff [6]) );
  DF3 \u_decoder/fir_filter/Q_data_add_4_buff_reg[5]  ( .D(n2466), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_4_buff [5]) );
  DF3 \u_decoder/fir_filter/Q_data_add_4_buff_reg[4]  ( .D(n2467), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_4_buff [4]) );
  DF3 \u_decoder/fir_filter/Q_data_add_4_buff_reg[3]  ( .D(n2468), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_4_buff [3]) );
  DF3 \u_decoder/fir_filter/Q_data_add_4_buff_reg[2]  ( .D(n2469), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_4_buff [2]) );
  DF3 \u_decoder/fir_filter/Q_data_add_4_buff_reg[1]  ( .D(n2470), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_4_buff [1]) );
  DF3 \u_decoder/fir_filter/Q_data_add_4_buff_reg[0]  ( .D(n2471), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_4_buff [0]), .QN(n115) );
  DF3 \u_decoder/fir_filter/Q_data_add_5_buff_reg[14]  ( .D(n2472), .C(inClock), .Q(\u_decoder/fir_filter/Q_data_add_5_buff [14]) );
  DF3 \u_decoder/fir_filter/Q_data_add_5_buff_reg[13]  ( .D(n2473), .C(inClock), .Q(\u_decoder/fir_filter/Q_data_add_5_buff [13]) );
  DF3 \u_decoder/fir_filter/Q_data_add_5_buff_reg[12]  ( .D(n2474), .C(inClock), .Q(\u_decoder/fir_filter/Q_data_add_5_buff [12]) );
  DF3 \u_decoder/fir_filter/Q_data_add_5_buff_reg[11]  ( .D(n2475), .C(inClock), .Q(\u_decoder/fir_filter/Q_data_add_5_buff [11]) );
  DF3 \u_decoder/fir_filter/Q_data_add_5_buff_reg[10]  ( .D(n2476), .C(inClock), .Q(\u_decoder/fir_filter/Q_data_add_5_buff [10]) );
  DF3 \u_decoder/fir_filter/Q_data_add_5_buff_reg[9]  ( .D(n2477), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_5_buff [9]) );
  DF3 \u_decoder/fir_filter/Q_data_add_5_buff_reg[8]  ( .D(n2478), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_5_buff [8]) );
  DF3 \u_decoder/fir_filter/Q_data_add_5_buff_reg[7]  ( .D(n2479), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_5_buff [7]) );
  DF3 \u_decoder/fir_filter/Q_data_add_5_buff_reg[6]  ( .D(n2480), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_5_buff [6]) );
  DF3 \u_decoder/fir_filter/Q_data_add_5_buff_reg[5]  ( .D(n2481), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_5_buff [5]) );
  DF3 \u_decoder/fir_filter/Q_data_add_5_buff_reg[4]  ( .D(n2482), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_5_buff [4]) );
  DF3 \u_decoder/fir_filter/Q_data_add_5_buff_reg[3]  ( .D(n2483), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_5_buff [3]) );
  DF3 \u_decoder/fir_filter/Q_data_add_5_buff_reg[2]  ( .D(n2484), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_5_buff [2]) );
  DF3 \u_decoder/fir_filter/Q_data_add_5_buff_reg[1]  ( .D(n2485), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_5_buff [1]) );
  DF3 \u_decoder/fir_filter/Q_data_add_5_buff_reg[0]  ( .D(n2486), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_5_buff [0]), .QN(n119) );
  DF3 \u_decoder/fir_filter/Q_data_add_6_buff_reg[14]  ( .D(n2487), .C(inClock), .Q(\u_decoder/fir_filter/Q_data_add_6_buff [14]) );
  DF3 \u_decoder/fir_filter/Q_data_add_6_buff_reg[13]  ( .D(n2488), .C(inClock), .Q(\u_decoder/fir_filter/Q_data_add_6_buff [13]) );
  DF3 \u_decoder/fir_filter/Q_data_add_6_buff_reg[12]  ( .D(n2489), .C(inClock), .Q(\u_decoder/fir_filter/Q_data_add_6_buff [12]) );
  DF3 \u_decoder/fir_filter/Q_data_add_6_buff_reg[11]  ( .D(n2490), .C(inClock), .Q(\u_decoder/fir_filter/Q_data_add_6_buff [11]) );
  DF3 \u_decoder/fir_filter/Q_data_add_6_buff_reg[10]  ( .D(n2491), .C(inClock), .Q(\u_decoder/fir_filter/Q_data_add_6_buff [10]) );
  DF3 \u_decoder/fir_filter/Q_data_add_6_buff_reg[9]  ( .D(n2492), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_6_buff [9]) );
  DF3 \u_decoder/fir_filter/Q_data_add_6_buff_reg[8]  ( .D(n2493), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_6_buff [8]) );
  DF3 \u_decoder/fir_filter/Q_data_add_6_buff_reg[7]  ( .D(n2494), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_6_buff [7]) );
  DF3 \u_decoder/fir_filter/Q_data_add_6_buff_reg[6]  ( .D(n2495), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_6_buff [6]) );
  DF3 \u_decoder/fir_filter/Q_data_add_6_buff_reg[5]  ( .D(n2496), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_6_buff [5]) );
  DF3 \u_decoder/fir_filter/Q_data_add_6_buff_reg[4]  ( .D(n2497), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_6_buff [4]) );
  DF3 \u_decoder/fir_filter/Q_data_add_6_buff_reg[3]  ( .D(n2498), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_6_buff [3]) );
  DF3 \u_decoder/fir_filter/Q_data_add_6_buff_reg[2]  ( .D(n2499), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_6_buff [2]) );
  DF3 \u_decoder/fir_filter/Q_data_add_6_buff_reg[1]  ( .D(n2500), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_6_buff [1]) );
  DF3 \u_decoder/fir_filter/Q_data_add_6_buff_reg[0]  ( .D(n2501), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_6_buff [0]), .QN(n114) );
  DF3 \u_decoder/fir_filter/Q_data_add_7_buff_reg[14]  ( .D(n2502), .C(inClock), .Q(\u_decoder/fir_filter/Q_data_add_7_buff [14]) );
  DF3 \u_decoder/fir_filter/Q_data_add_7_buff_reg[13]  ( .D(n2503), .C(inClock), .Q(\u_decoder/fir_filter/Q_data_add_7_buff [13]) );
  DF3 \u_decoder/fir_filter/Q_data_add_7_buff_reg[12]  ( .D(n2504), .C(inClock), .Q(\u_decoder/fir_filter/Q_data_add_7_buff [12]) );
  DF3 \u_decoder/fir_filter/Q_data_add_7_buff_reg[11]  ( .D(n2505), .C(inClock), .Q(\u_decoder/fir_filter/Q_data_add_7_buff [11]) );
  DF3 \u_decoder/fir_filter/Q_data_add_7_buff_reg[10]  ( .D(n2506), .C(inClock), .Q(\u_decoder/fir_filter/Q_data_add_7_buff [10]) );
  DF3 \u_decoder/fir_filter/Q_data_add_7_buff_reg[9]  ( .D(n2507), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_7_buff [9]) );
  DF3 \u_decoder/fir_filter/Q_data_add_7_buff_reg[8]  ( .D(n2508), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_7_buff [8]) );
  DF3 \u_decoder/fir_filter/Q_data_add_7_buff_reg[7]  ( .D(n2509), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_7_buff [7]) );
  DF3 \u_decoder/fir_filter/Q_data_add_7_buff_reg[6]  ( .D(n2510), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_7_buff [6]) );
  DF3 \u_decoder/fir_filter/Q_data_add_7_buff_reg[5]  ( .D(n2511), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_7_buff [5]) );
  DF3 \u_decoder/fir_filter/Q_data_add_7_buff_reg[4]  ( .D(n2512), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_7_buff [4]) );
  DF3 \u_decoder/fir_filter/Q_data_add_7_buff_reg[3]  ( .D(n2513), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_7_buff [3]) );
  DF3 \u_decoder/fir_filter/Q_data_add_7_buff_reg[2]  ( .D(n2514), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_7_buff [2]) );
  DF3 \u_decoder/fir_filter/Q_data_add_7_buff_reg[1]  ( .D(n2515), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_7_buff [1]) );
  DF3 \u_decoder/fir_filter/Q_data_add_7_buff_reg[0]  ( .D(n2516), .C(inClock), 
        .Q(\u_decoder/fir_filter/Q_data_add_7_buff [0]), .QN(n113) );
  DF3 \u_decoder/fir_filter/Q_data_mult_8_buff_reg[0]  ( .D(
        \u_decoder/fir_filter/n1155 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_8_buff [0]), .QN(n107) );
  DF3 \u_decoder/fir_filter/Q_data_mult_8_buff_reg[1]  ( .D(
        \u_decoder/fir_filter/n1156 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_8_buff [1]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_8_buff_reg[2]  ( .D(
        \u_decoder/fir_filter/n1157 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_8_buff [2]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_8_buff_reg[3]  ( .D(
        \u_decoder/fir_filter/n1158 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_8_buff [3]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_8_buff_reg[4]  ( .D(
        \u_decoder/fir_filter/n1159 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_8_buff [4]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_8_buff_reg[5]  ( .D(
        \u_decoder/fir_filter/n1160 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_8_buff [5]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_8_buff_reg[6]  ( .D(
        \u_decoder/fir_filter/n1161 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_8_buff [6]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_8_buff_reg[7]  ( .D(
        \u_decoder/fir_filter/n1162 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_8_buff [7]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_8_buff_reg[8]  ( .D(
        \u_decoder/fir_filter/n1163 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_8_buff [8]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_8_buff_reg[9]  ( .D(
        \u_decoder/fir_filter/n1164 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_8_buff [9]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_8_buff_reg[10]  ( .D(
        \u_decoder/fir_filter/n1165 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_8_buff [10]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_8_buff_reg[11]  ( .D(
        \u_decoder/fir_filter/n1166 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_8_buff [11]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_8_buff_reg[12]  ( .D(
        \u_decoder/fir_filter/n1167 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_8_buff [12]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_8_buff_reg[13]  ( .D(
        \u_decoder/fir_filter/n1168 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_8_buff [13]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_8_buff_reg[14]  ( .D(
        \u_decoder/fir_filter/n1169 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_8_buff [14]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_8_delay_reg[0]  ( .D(
        \u_decoder/fir_filter/n1176 ), .C(inClock), .QN(
        \u_decoder/fir_filter/n442 ) );
  DF3 \u_decoder/fir_filter/Q_data_mult_8_delay_reg[1]  ( .D(
        \u_decoder/fir_filter/n1177 ), .C(inClock), .QN(
        \u_decoder/fir_filter/n441 ) );
  DF3 \u_decoder/fir_filter/Q_data_mult_8_delay_reg[2]  ( .D(
        \u_decoder/fir_filter/n1178 ), .C(inClock), .QN(
        \u_decoder/fir_filter/n440 ) );
  DF3 \u_decoder/fir_filter/Q_data_mult_8_delay_reg[3]  ( .D(
        \u_decoder/fir_filter/n1179 ), .C(inClock), .QN(
        \u_decoder/fir_filter/n439 ) );
  DF3 \u_decoder/fir_filter/Q_data_mult_8_delay_reg[4]  ( .D(
        \u_decoder/fir_filter/n1180 ), .C(inClock), .QN(
        \u_decoder/fir_filter/n438 ) );
  DF3 \u_decoder/fir_filter/Q_data_mult_8_delay_reg[5]  ( .D(
        \u_decoder/fir_filter/n1181 ), .C(inClock), .QN(
        \u_decoder/fir_filter/n437 ) );
  DF3 \u_decoder/fir_filter/Q_data_mult_8_delay_reg[6]  ( .D(
        \u_decoder/fir_filter/n1182 ), .C(inClock), .QN(
        \u_decoder/fir_filter/n436 ) );
  DF3 \u_decoder/fir_filter/Q_data_mult_8_delay_reg[7]  ( .D(
        \u_decoder/fir_filter/n1183 ), .C(inClock), .QN(
        \u_decoder/fir_filter/n435 ) );
  DF3 \u_decoder/fir_filter/Q_data_mult_8_delay_reg[8]  ( .D(
        \u_decoder/fir_filter/n1184 ), .C(inClock), .QN(
        \u_decoder/fir_filter/n434 ) );
  DF3 \u_decoder/fir_filter/Q_data_mult_8_delay_reg[9]  ( .D(
        \u_decoder/fir_filter/n1185 ), .C(inClock), .QN(
        \u_decoder/fir_filter/n433 ) );
  DF3 \u_decoder/fir_filter/Q_data_mult_8_delay_reg[10]  ( .D(
        \u_decoder/fir_filter/n1186 ), .C(inClock), .QN(
        \u_decoder/fir_filter/n432 ) );
  DF3 \u_decoder/fir_filter/Q_data_mult_8_delay_reg[11]  ( .D(
        \u_decoder/fir_filter/n1187 ), .C(inClock), .QN(
        \u_decoder/fir_filter/n431 ) );
  DF3 \u_decoder/fir_filter/Q_data_mult_8_delay_reg[12]  ( .D(
        \u_decoder/fir_filter/n1188 ), .C(inClock), .QN(
        \u_decoder/fir_filter/n430 ) );
  DF3 \u_decoder/fir_filter/Q_data_mult_8_delay_reg[13]  ( .D(
        \u_decoder/fir_filter/n1189 ), .C(inClock), .QN(
        \u_decoder/fir_filter/n429 ) );
  DF3 \u_decoder/fir_filter/Q_data_mult_8_delay_reg[14]  ( .D(
        \u_decoder/fir_filter/n1190 ), .C(inClock), .QN(
        \u_decoder/fir_filter/n428 ) );
  DF3 \u_decoder/fir_filter/Q_data_mult_7_buff_reg[0]  ( .D(
        \u_decoder/fir_filter/n1192 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_7_buff [0]), .QN(n32) );
  DF3 \u_decoder/fir_filter/Q_data_mult_7_buff_reg[1]  ( .D(
        \u_decoder/fir_filter/n1193 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_7_buff [1]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_7_buff_reg[2]  ( .D(
        \u_decoder/fir_filter/n1194 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_7_buff [2]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_7_buff_reg[3]  ( .D(
        \u_decoder/fir_filter/n1195 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_7_buff [3]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_7_buff_reg[4]  ( .D(
        \u_decoder/fir_filter/n1196 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_7_buff [4]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_7_buff_reg[5]  ( .D(
        \u_decoder/fir_filter/n1197 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_7_buff [5]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_7_buff_reg[6]  ( .D(
        \u_decoder/fir_filter/n1198 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_7_buff [6]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_7_buff_reg[7]  ( .D(
        \u_decoder/fir_filter/n1199 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_7_buff [7]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_7_buff_reg[8]  ( .D(
        \u_decoder/fir_filter/n1200 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_7_buff [8]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_7_buff_reg[9]  ( .D(
        \u_decoder/fir_filter/n1201 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_7_buff [9]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_7_buff_reg[10]  ( .D(
        \u_decoder/fir_filter/n1202 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_7_buff [10]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_7_buff_reg[11]  ( .D(
        \u_decoder/fir_filter/n1203 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_7_buff [11]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_7_buff_reg[12]  ( .D(
        \u_decoder/fir_filter/n1204 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_7_buff [12]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_7_buff_reg[13]  ( .D(
        \u_decoder/fir_filter/n1205 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_7_buff [13]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_7_buff_reg[14]  ( .D(
        \u_decoder/fir_filter/n1206 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_7_buff [14]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_6_buff_reg[0]  ( .D(n2517), .C(inClock), .Q(\u_decoder/fir_filter/Q_data_mult_6_buff [0]), .QN(n33) );
  DF3 \u_decoder/fir_filter/Q_data_mult_6_buff_reg[1]  ( .D(
        \u_decoder/fir_filter/n1209 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_6_buff [1]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_6_buff_reg[2]  ( .D(
        \u_decoder/fir_filter/n1210 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_6_buff [2]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_6_buff_reg[3]  ( .D(
        \u_decoder/fir_filter/n1211 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_6_buff [3]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_6_buff_reg[4]  ( .D(
        \u_decoder/fir_filter/n1212 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_6_buff [4]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_6_buff_reg[5]  ( .D(
        \u_decoder/fir_filter/n1213 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_6_buff [5]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_6_buff_reg[6]  ( .D(
        \u_decoder/fir_filter/n1214 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_6_buff [6]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_6_buff_reg[7]  ( .D(
        \u_decoder/fir_filter/n1215 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_6_buff [7]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_6_buff_reg[8]  ( .D(
        \u_decoder/fir_filter/n1216 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_6_buff [8]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_6_buff_reg[9]  ( .D(
        \u_decoder/fir_filter/n1217 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_6_buff [9]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_6_buff_reg[10]  ( .D(
        \u_decoder/fir_filter/n1218 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_6_buff [10]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_6_buff_reg[11]  ( .D(
        \u_decoder/fir_filter/n1219 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_6_buff [11]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_6_buff_reg[12]  ( .D(
        \u_decoder/fir_filter/n1220 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_6_buff [12]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_6_buff_reg[13]  ( .D(
        \u_decoder/fir_filter/n1221 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_6_buff [13]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_6_buff_reg[14]  ( .D(
        \u_decoder/fir_filter/n1222 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_6_buff [14]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_5_buff_reg[0]  ( .D(
        \u_decoder/fir_filter/n1224 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_5_buff [0]), .QN(n34) );
  DF3 \u_decoder/fir_filter/Q_data_mult_5_buff_reg[1]  ( .D(
        \u_decoder/fir_filter/n1225 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_5_buff [1]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_5_buff_reg[2]  ( .D(
        \u_decoder/fir_filter/n1226 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_5_buff [2]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_5_buff_reg[3]  ( .D(
        \u_decoder/fir_filter/n1227 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_5_buff [3]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_5_buff_reg[4]  ( .D(
        \u_decoder/fir_filter/n1228 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_5_buff [4]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_5_buff_reg[5]  ( .D(
        \u_decoder/fir_filter/n1229 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_5_buff [5]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_5_buff_reg[6]  ( .D(
        \u_decoder/fir_filter/n1230 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_5_buff [6]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_5_buff_reg[7]  ( .D(
        \u_decoder/fir_filter/n1231 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_5_buff [7]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_5_buff_reg[8]  ( .D(
        \u_decoder/fir_filter/n1232 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_5_buff [8]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_5_buff_reg[9]  ( .D(
        \u_decoder/fir_filter/n1233 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_5_buff [9]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_5_buff_reg[10]  ( .D(
        \u_decoder/fir_filter/n1234 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_5_buff [10]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_5_buff_reg[11]  ( .D(
        \u_decoder/fir_filter/n1235 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_5_buff [11]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_5_buff_reg[12]  ( .D(
        \u_decoder/fir_filter/n1236 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_5_buff [12]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_5_buff_reg[13]  ( .D(
        \u_decoder/fir_filter/n1237 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_5_buff [13]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_5_buff_reg[14]  ( .D(
        \u_decoder/fir_filter/n1238 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_5_buff [14]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_4_buff_reg[0]  ( .D(n2326), .C(inClock), .Q(\u_decoder/fir_filter/Q_data_mult_4_buff [0]), .QN(n39) );
  DF3 \u_decoder/fir_filter/Q_data_mult_4_buff_reg[1]  ( .D(n2369), .C(inClock), .Q(\u_decoder/fir_filter/Q_data_mult_4_buff [1]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_4_buff_reg[2]  ( .D(n2371), .C(inClock), .Q(\u_decoder/fir_filter/Q_data_mult_4_buff [2]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_4_buff_reg[3]  ( .D(n2344), .C(inClock), .Q(\u_decoder/fir_filter/Q_data_mult_4_buff [3]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_4_buff_reg[4]  ( .D(n2343), .C(inClock), .Q(\u_decoder/fir_filter/Q_data_mult_4_buff [4]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_4_buff_reg[5]  ( .D(n2342), .C(inClock), .Q(\u_decoder/fir_filter/Q_data_mult_4_buff [5]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_4_buff_reg[6]  ( .D(n2341), .C(inClock), .Q(\u_decoder/fir_filter/Q_data_mult_4_buff [6]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_4_buff_reg[7]  ( .D(n2340), .C(inClock), .Q(\u_decoder/fir_filter/Q_data_mult_4_buff [7]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_4_buff_reg[8]  ( .D(n2339), .C(inClock), .Q(\u_decoder/fir_filter/Q_data_mult_4_buff [8]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_4_buff_reg[9]  ( .D(n2338), .C(inClock), .Q(\u_decoder/fir_filter/Q_data_mult_4_buff [9]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_4_buff_reg[10]  ( .D(n2336), .C(
        inClock), .Q(\u_decoder/fir_filter/Q_data_mult_4_buff [10]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_4_buff_reg[11]  ( .D(n2332), .C(
        inClock), .Q(\u_decoder/fir_filter/Q_data_mult_4_buff [11]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_4_buff_reg[12]  ( .D(n2327), .C(
        inClock), .Q(\u_decoder/fir_filter/Q_data_mult_4_buff [12]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_4_buff_reg[13]  ( .D(n2329), .C(
        inClock), .Q(\u_decoder/fir_filter/Q_data_mult_4_buff [13]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_4_buff_reg[14]  ( .D(n2330), .C(
        inClock), .Q(\u_decoder/fir_filter/Q_data_mult_4_buff [14]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_3_buff_reg[0]  ( .D(
        \u_decoder/fir_filter/n1240 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_3_buff [0]), .QN(n35) );
  DF3 \u_decoder/fir_filter/Q_data_mult_3_buff_reg[1]  ( .D(
        \u_decoder/fir_filter/n1241 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_3_buff [1]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_3_buff_reg[2]  ( .D(
        \u_decoder/fir_filter/n1242 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_3_buff [2]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_3_buff_reg[3]  ( .D(
        \u_decoder/fir_filter/n1243 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_3_buff [3]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_3_buff_reg[4]  ( .D(
        \u_decoder/fir_filter/n1244 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_3_buff [4]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_3_buff_reg[5]  ( .D(
        \u_decoder/fir_filter/n1245 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_3_buff [5]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_3_buff_reg[6]  ( .D(
        \u_decoder/fir_filter/n1246 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_3_buff [6]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_3_buff_reg[7]  ( .D(
        \u_decoder/fir_filter/n1247 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_3_buff [7]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_3_buff_reg[8]  ( .D(
        \u_decoder/fir_filter/n1248 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_3_buff [8]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_3_buff_reg[9]  ( .D(
        \u_decoder/fir_filter/n1249 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_3_buff [9]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_3_buff_reg[10]  ( .D(
        \u_decoder/fir_filter/n1250 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_3_buff [10]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_3_buff_reg[11]  ( .D(
        \u_decoder/fir_filter/n1251 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_3_buff [11]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_3_buff_reg[12]  ( .D(
        \u_decoder/fir_filter/n1252 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_3_buff [12]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_3_buff_reg[13]  ( .D(
        \u_decoder/fir_filter/n1253 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_3_buff [13]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_3_buff_reg[14]  ( .D(
        \u_decoder/fir_filter/n1254 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_3_buff [14]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_2_buff_reg[0]  ( .D(n2518), .C(inClock), .Q(\u_decoder/fir_filter/Q_data_mult_2_buff [0]), .QN(n36) );
  DF3 \u_decoder/fir_filter/Q_data_mult_2_buff_reg[1]  ( .D(
        \u_decoder/fir_filter/n1257 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_2_buff [1]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_2_buff_reg[2]  ( .D(
        \u_decoder/fir_filter/n1258 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_2_buff [2]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_2_buff_reg[3]  ( .D(
        \u_decoder/fir_filter/n1259 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_2_buff [3]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_2_buff_reg[4]  ( .D(
        \u_decoder/fir_filter/n1260 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_2_buff [4]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_2_buff_reg[5]  ( .D(
        \u_decoder/fir_filter/n1261 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_2_buff [5]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_2_buff_reg[6]  ( .D(
        \u_decoder/fir_filter/n1262 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_2_buff [6]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_2_buff_reg[7]  ( .D(
        \u_decoder/fir_filter/n1263 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_2_buff [7]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_2_buff_reg[8]  ( .D(
        \u_decoder/fir_filter/n1264 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_2_buff [8]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_2_buff_reg[9]  ( .D(
        \u_decoder/fir_filter/n1265 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_2_buff [9]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_2_buff_reg[10]  ( .D(
        \u_decoder/fir_filter/n1266 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_2_buff [10]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_2_buff_reg[11]  ( .D(
        \u_decoder/fir_filter/n1267 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_2_buff [11]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_2_buff_reg[12]  ( .D(
        \u_decoder/fir_filter/n1268 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_2_buff [12]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_2_buff_reg[13]  ( .D(
        \u_decoder/fir_filter/n1269 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_2_buff [13]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_2_buff_reg[14]  ( .D(
        \u_decoder/fir_filter/n1270 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_2_buff [14]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_1_buff_reg[0]  ( .D(
        \u_decoder/fir_filter/n1272 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_1_buff [0]), .QN(n37) );
  DF3 \u_decoder/fir_filter/Q_data_mult_1_buff_reg[1]  ( .D(
        \u_decoder/fir_filter/n1273 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_1_buff [1]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_1_buff_reg[2]  ( .D(
        \u_decoder/fir_filter/n1274 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_1_buff [2]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_1_buff_reg[3]  ( .D(
        \u_decoder/fir_filter/n1275 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_1_buff [3]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_1_buff_reg[4]  ( .D(
        \u_decoder/fir_filter/n1276 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_1_buff [4]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_1_buff_reg[5]  ( .D(
        \u_decoder/fir_filter/n1277 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_1_buff [5]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_1_buff_reg[6]  ( .D(
        \u_decoder/fir_filter/n1278 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_1_buff [6]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_1_buff_reg[7]  ( .D(
        \u_decoder/fir_filter/n1279 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_1_buff [7]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_1_buff_reg[8]  ( .D(
        \u_decoder/fir_filter/n1280 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_1_buff [8]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_1_buff_reg[9]  ( .D(
        \u_decoder/fir_filter/n1281 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_1_buff [9]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_1_buff_reg[10]  ( .D(
        \u_decoder/fir_filter/n1282 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_1_buff [10]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_1_buff_reg[11]  ( .D(
        \u_decoder/fir_filter/n1283 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_1_buff [11]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_1_buff_reg[12]  ( .D(
        \u_decoder/fir_filter/n1284 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_1_buff [12]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_1_buff_reg[13]  ( .D(
        \u_decoder/fir_filter/n1285 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_1_buff [13]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_1_buff_reg[14]  ( .D(
        \u_decoder/fir_filter/n1286 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_1_buff [14]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_0_buff_reg[0]  ( .D(
        \u_decoder/fir_filter/n1288 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_0_buff [0]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_0_buff_reg[1]  ( .D(
        \u_decoder/fir_filter/n1289 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_0_buff [1]), .QN(n93) );
  DF3 \u_decoder/fir_filter/Q_data_mult_0_buff_reg[2]  ( .D(
        \u_decoder/fir_filter/n1290 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_0_buff [2]), .QN(n91) );
  DF3 \u_decoder/fir_filter/Q_data_mult_0_buff_reg[3]  ( .D(
        \u_decoder/fir_filter/n1291 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_0_buff [3]), .QN(n135) );
  DF3 \u_decoder/fir_filter/Q_data_mult_0_buff_reg[4]  ( .D(
        \u_decoder/fir_filter/n1292 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_0_buff [4]), .QN(n136) );
  DF3 \u_decoder/fir_filter/Q_data_mult_0_buff_reg[5]  ( .D(
        \u_decoder/fir_filter/n1293 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_0_buff [5]), .QN(n137) );
  DF3 \u_decoder/fir_filter/Q_data_mult_0_buff_reg[6]  ( .D(
        \u_decoder/fir_filter/n1294 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_0_buff [6]), .QN(n177) );
  DF3 \u_decoder/fir_filter/Q_data_mult_0_buff_reg[7]  ( .D(
        \u_decoder/fir_filter/n1295 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_0_buff [7]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_0_buff_reg[8]  ( .D(
        \u_decoder/fir_filter/n1296 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_0_buff [8]), .QN(n223) );
  DF3 \u_decoder/fir_filter/Q_data_mult_0_buff_reg[9]  ( .D(
        \u_decoder/fir_filter/n1297 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_0_buff [9]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_0_buff_reg[10]  ( .D(
        \u_decoder/fir_filter/n1298 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_0_buff [10]), .QN(n264) );
  DF3 \u_decoder/fir_filter/Q_data_mult_0_buff_reg[11]  ( .D(
        \u_decoder/fir_filter/n1299 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_0_buff [11]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_0_buff_reg[12]  ( .D(
        \u_decoder/fir_filter/n1300 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_0_buff [12]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_0_buff_reg[13]  ( .D(
        \u_decoder/fir_filter/n1301 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_0_buff [13]) );
  DF3 \u_decoder/fir_filter/Q_data_mult_0_buff_reg[14]  ( .D(
        \u_decoder/fir_filter/n1302 ), .C(inClock), .Q(
        \u_decoder/fir_filter/Q_data_mult_0_buff [14]) );
  DF3 \u_decoder/fir_filter/o_I_postfilter_reg[3]  ( .D(n2519), .C(inClock), 
        .Q(sig_decod_outI[3]) );
  DF3 \u_decoder/fir_filter/o_I_postfilter_reg[2]  ( .D(n2520), .C(inClock), 
        .Q(sig_decod_outI[2]) );
  DF3 \u_decoder/fir_filter/o_I_postfilter_reg[1]  ( .D(n2521), .C(inClock), 
        .Q(sig_decod_outI[1]) );
  DF3 \u_decoder/fir_filter/o_I_postfilter_reg[0]  ( .D(n2522), .C(inClock), 
        .Q(sig_decod_outI[0]) );
  DF3 \u_decoder/fir_filter/I_data_add_1_buff_reg[14]  ( .D(n2523), .C(inClock), .Q(\u_decoder/fir_filter/I_data_add_1_buff [14]) );
  DF3 \u_decoder/fir_filter/I_data_add_1_buff_reg[13]  ( .D(n2524), .C(inClock), .Q(\u_decoder/fir_filter/I_data_add_1_buff [13]) );
  DF3 \u_decoder/fir_filter/I_data_add_1_buff_reg[12]  ( .D(n2525), .C(inClock), .Q(\u_decoder/fir_filter/I_data_add_1_buff [12]) );
  DF3 \u_decoder/fir_filter/I_data_add_1_buff_reg[11]  ( .D(n2526), .C(inClock), .Q(\u_decoder/fir_filter/I_data_add_1_buff [11]) );
  DF3 \u_decoder/fir_filter/I_data_add_1_buff_reg[10]  ( .D(n2527), .C(inClock), .Q(\u_decoder/fir_filter/I_data_add_1_buff [10]) );
  DF3 \u_decoder/fir_filter/I_data_add_1_buff_reg[9]  ( .D(n2530), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_1_buff [9]) );
  DF3 \u_decoder/fir_filter/I_data_add_1_buff_reg[8]  ( .D(n2531), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_1_buff [8]) );
  DF3 \u_decoder/fir_filter/I_data_add_1_buff_reg[7]  ( .D(n2534), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_1_buff [7]) );
  DF3 \u_decoder/fir_filter/I_data_add_1_buff_reg[6]  ( .D(n2535), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_1_buff [6]) );
  DF3 \u_decoder/fir_filter/I_data_add_1_buff_reg[5]  ( .D(n2537), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_1_buff [5]) );
  DF3 \u_decoder/fir_filter/I_data_add_1_buff_reg[4]  ( .D(n2539), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_1_buff [4]) );
  DF3 \u_decoder/fir_filter/I_data_add_1_buff_reg[3]  ( .D(n2541), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_1_buff [3]) );
  DF3 \u_decoder/fir_filter/I_data_add_1_buff_reg[2]  ( .D(n2543), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_1_buff [2]) );
  DF3 \u_decoder/fir_filter/I_data_add_1_buff_reg[1]  ( .D(n2545), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_1_buff [1]), .QN(n25) );
  DF3 \u_decoder/fir_filter/I_data_add_1_buff_reg[0]  ( .D(n2546), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_1_buff [0]) );
  DF3 \u_decoder/fir_filter/I_data_add_2_buff_reg[14]  ( .D(n2547), .C(inClock), .Q(\u_decoder/fir_filter/I_data_add_2_buff [14]) );
  DF3 \u_decoder/fir_filter/I_data_add_2_buff_reg[13]  ( .D(n2548), .C(inClock), .Q(\u_decoder/fir_filter/I_data_add_2_buff [13]) );
  DF3 \u_decoder/fir_filter/I_data_add_2_buff_reg[12]  ( .D(n2549), .C(inClock), .Q(\u_decoder/fir_filter/I_data_add_2_buff [12]) );
  DF3 \u_decoder/fir_filter/I_data_add_2_buff_reg[11]  ( .D(n2550), .C(inClock), .Q(\u_decoder/fir_filter/I_data_add_2_buff [11]) );
  DF3 \u_decoder/fir_filter/I_data_add_2_buff_reg[10]  ( .D(n2551), .C(inClock), .Q(\u_decoder/fir_filter/I_data_add_2_buff [10]) );
  DF3 \u_decoder/fir_filter/I_data_add_2_buff_reg[9]  ( .D(n2552), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_2_buff [9]) );
  DF3 \u_decoder/fir_filter/I_data_add_2_buff_reg[8]  ( .D(n2553), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_2_buff [8]) );
  DF3 \u_decoder/fir_filter/I_data_add_2_buff_reg[7]  ( .D(n2554), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_2_buff [7]) );
  DF3 \u_decoder/fir_filter/I_data_add_2_buff_reg[6]  ( .D(n2555), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_2_buff [6]) );
  DF3 \u_decoder/fir_filter/I_data_add_2_buff_reg[5]  ( .D(n2556), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_2_buff [5]) );
  DF3 \u_decoder/fir_filter/I_data_add_2_buff_reg[4]  ( .D(n2557), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_2_buff [4]) );
  DF3 \u_decoder/fir_filter/I_data_add_2_buff_reg[3]  ( .D(n2558), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_2_buff [3]) );
  DF3 \u_decoder/fir_filter/I_data_add_2_buff_reg[2]  ( .D(n2559), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_2_buff [2]) );
  DF3 \u_decoder/fir_filter/I_data_add_2_buff_reg[1]  ( .D(n2560), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_2_buff [1]) );
  DF3 \u_decoder/fir_filter/I_data_add_2_buff_reg[0]  ( .D(n2561), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_2_buff [0]), .QN(n112) );
  DF3 \u_decoder/fir_filter/I_data_add_3_buff_reg[14]  ( .D(n2562), .C(inClock), .Q(\u_decoder/fir_filter/I_data_add_3_buff [14]) );
  DF3 \u_decoder/fir_filter/I_data_add_3_buff_reg[13]  ( .D(n2563), .C(inClock), .Q(\u_decoder/fir_filter/I_data_add_3_buff [13]) );
  DF3 \u_decoder/fir_filter/I_data_add_3_buff_reg[12]  ( .D(n2564), .C(inClock), .Q(\u_decoder/fir_filter/I_data_add_3_buff [12]) );
  DF3 \u_decoder/fir_filter/I_data_add_3_buff_reg[11]  ( .D(n2565), .C(inClock), .Q(\u_decoder/fir_filter/I_data_add_3_buff [11]) );
  DF3 \u_decoder/fir_filter/I_data_add_3_buff_reg[10]  ( .D(n2566), .C(inClock), .Q(\u_decoder/fir_filter/I_data_add_3_buff [10]) );
  DF3 \u_decoder/fir_filter/I_data_add_3_buff_reg[9]  ( .D(n2567), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_3_buff [9]) );
  DF3 \u_decoder/fir_filter/I_data_add_3_buff_reg[8]  ( .D(n2568), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_3_buff [8]) );
  DF3 \u_decoder/fir_filter/I_data_add_3_buff_reg[7]  ( .D(n2569), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_3_buff [7]) );
  DF3 \u_decoder/fir_filter/I_data_add_3_buff_reg[6]  ( .D(n2570), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_3_buff [6]) );
  DF3 \u_decoder/fir_filter/I_data_add_3_buff_reg[5]  ( .D(n2571), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_3_buff [5]) );
  DF3 \u_decoder/fir_filter/I_data_add_3_buff_reg[4]  ( .D(n2572), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_3_buff [4]) );
  DF3 \u_decoder/fir_filter/I_data_add_3_buff_reg[3]  ( .D(n2573), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_3_buff [3]) );
  DF3 \u_decoder/fir_filter/I_data_add_3_buff_reg[2]  ( .D(n2574), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_3_buff [2]) );
  DF3 \u_decoder/fir_filter/I_data_add_3_buff_reg[1]  ( .D(n2575), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_3_buff [1]) );
  DF3 \u_decoder/fir_filter/I_data_add_3_buff_reg[0]  ( .D(n2576), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_3_buff [0]), .QN(n111) );
  DF3 \u_decoder/fir_filter/I_data_add_4_buff_reg[14]  ( .D(n2577), .C(inClock), .Q(\u_decoder/fir_filter/I_data_add_4_buff [14]) );
  DF3 \u_decoder/fir_filter/I_data_add_4_buff_reg[13]  ( .D(n2578), .C(inClock), .Q(\u_decoder/fir_filter/I_data_add_4_buff [13]) );
  DF3 \u_decoder/fir_filter/I_data_add_4_buff_reg[12]  ( .D(n2579), .C(inClock), .Q(\u_decoder/fir_filter/I_data_add_4_buff [12]) );
  DF3 \u_decoder/fir_filter/I_data_add_4_buff_reg[11]  ( .D(n2580), .C(inClock), .Q(\u_decoder/fir_filter/I_data_add_4_buff [11]) );
  DF3 \u_decoder/fir_filter/I_data_add_4_buff_reg[10]  ( .D(n2581), .C(inClock), .Q(\u_decoder/fir_filter/I_data_add_4_buff [10]) );
  DF3 \u_decoder/fir_filter/I_data_add_4_buff_reg[9]  ( .D(n2582), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_4_buff [9]) );
  DF3 \u_decoder/fir_filter/I_data_add_4_buff_reg[8]  ( .D(n2583), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_4_buff [8]) );
  DF3 \u_decoder/fir_filter/I_data_add_4_buff_reg[7]  ( .D(n2584), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_4_buff [7]) );
  DF3 \u_decoder/fir_filter/I_data_add_4_buff_reg[6]  ( .D(n2585), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_4_buff [6]) );
  DF3 \u_decoder/fir_filter/I_data_add_4_buff_reg[5]  ( .D(n2586), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_4_buff [5]) );
  DF3 \u_decoder/fir_filter/I_data_add_4_buff_reg[4]  ( .D(n2587), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_4_buff [4]) );
  DF3 \u_decoder/fir_filter/I_data_add_4_buff_reg[3]  ( .D(n2588), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_4_buff [3]) );
  DF3 \u_decoder/fir_filter/I_data_add_4_buff_reg[2]  ( .D(n2589), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_4_buff [2]) );
  DF3 \u_decoder/fir_filter/I_data_add_4_buff_reg[1]  ( .D(n2590), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_4_buff [1]) );
  DF3 \u_decoder/fir_filter/I_data_add_4_buff_reg[0]  ( .D(n2591), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_4_buff [0]), .QN(n110) );
  DF3 \u_decoder/fir_filter/I_data_add_5_buff_reg[14]  ( .D(n2592), .C(inClock), .Q(\u_decoder/fir_filter/I_data_add_5_buff [14]) );
  DF3 \u_decoder/fir_filter/I_data_add_5_buff_reg[13]  ( .D(n2593), .C(inClock), .Q(\u_decoder/fir_filter/I_data_add_5_buff [13]) );
  DF3 \u_decoder/fir_filter/I_data_add_5_buff_reg[12]  ( .D(n2594), .C(inClock), .Q(\u_decoder/fir_filter/I_data_add_5_buff [12]) );
  DF3 \u_decoder/fir_filter/I_data_add_5_buff_reg[11]  ( .D(n2595), .C(inClock), .Q(\u_decoder/fir_filter/I_data_add_5_buff [11]) );
  DF3 \u_decoder/fir_filter/I_data_add_5_buff_reg[10]  ( .D(n2596), .C(inClock), .Q(\u_decoder/fir_filter/I_data_add_5_buff [10]) );
  DF3 \u_decoder/fir_filter/I_data_add_5_buff_reg[9]  ( .D(n2597), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_5_buff [9]) );
  DF3 \u_decoder/fir_filter/I_data_add_5_buff_reg[8]  ( .D(n2598), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_5_buff [8]) );
  DF3 \u_decoder/fir_filter/I_data_add_5_buff_reg[7]  ( .D(n2599), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_5_buff [7]) );
  DF3 \u_decoder/fir_filter/I_data_add_5_buff_reg[6]  ( .D(n2600), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_5_buff [6]) );
  DF3 \u_decoder/fir_filter/I_data_add_5_buff_reg[5]  ( .D(n2601), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_5_buff [5]) );
  DF3 \u_decoder/fir_filter/I_data_add_5_buff_reg[4]  ( .D(n2602), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_5_buff [4]) );
  DF3 \u_decoder/fir_filter/I_data_add_5_buff_reg[3]  ( .D(n2603), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_5_buff [3]) );
  DF3 \u_decoder/fir_filter/I_data_add_5_buff_reg[2]  ( .D(n2604), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_5_buff [2]) );
  DF3 \u_decoder/fir_filter/I_data_add_5_buff_reg[1]  ( .D(n2605), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_5_buff [1]) );
  DF3 \u_decoder/fir_filter/I_data_add_5_buff_reg[0]  ( .D(n2606), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_5_buff [0]), .QN(n118) );
  DF3 \u_decoder/fir_filter/I_data_add_6_buff_reg[14]  ( .D(n2607), .C(inClock), .Q(\u_decoder/fir_filter/I_data_add_6_buff [14]) );
  DF3 \u_decoder/fir_filter/I_data_add_6_buff_reg[13]  ( .D(n2608), .C(inClock), .Q(\u_decoder/fir_filter/I_data_add_6_buff [13]) );
  DF3 \u_decoder/fir_filter/I_data_add_6_buff_reg[12]  ( .D(n2609), .C(inClock), .Q(\u_decoder/fir_filter/I_data_add_6_buff [12]) );
  DF3 \u_decoder/fir_filter/I_data_add_6_buff_reg[11]  ( .D(n2610), .C(inClock), .Q(\u_decoder/fir_filter/I_data_add_6_buff [11]) );
  DF3 \u_decoder/fir_filter/I_data_add_6_buff_reg[10]  ( .D(n2611), .C(inClock), .Q(\u_decoder/fir_filter/I_data_add_6_buff [10]) );
  DF3 \u_decoder/fir_filter/I_data_add_6_buff_reg[9]  ( .D(n2612), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_6_buff [9]) );
  DF3 \u_decoder/fir_filter/I_data_add_6_buff_reg[8]  ( .D(n2613), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_6_buff [8]) );
  DF3 \u_decoder/fir_filter/I_data_add_6_buff_reg[7]  ( .D(n2614), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_6_buff [7]) );
  DF3 \u_decoder/fir_filter/I_data_add_6_buff_reg[6]  ( .D(n2615), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_6_buff [6]) );
  DF3 \u_decoder/fir_filter/I_data_add_6_buff_reg[5]  ( .D(n2616), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_6_buff [5]) );
  DF3 \u_decoder/fir_filter/I_data_add_6_buff_reg[4]  ( .D(n2617), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_6_buff [4]) );
  DF3 \u_decoder/fir_filter/I_data_add_6_buff_reg[3]  ( .D(n2618), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_6_buff [3]) );
  DF3 \u_decoder/fir_filter/I_data_add_6_buff_reg[2]  ( .D(n2619), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_6_buff [2]) );
  DF3 \u_decoder/fir_filter/I_data_add_6_buff_reg[1]  ( .D(n2620), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_6_buff [1]) );
  DF3 \u_decoder/fir_filter/I_data_add_6_buff_reg[0]  ( .D(n2621), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_6_buff [0]), .QN(n109) );
  DF3 \u_decoder/fir_filter/I_data_add_7_buff_reg[14]  ( .D(n2622), .C(inClock), .Q(\u_decoder/fir_filter/I_data_add_7_buff [14]) );
  DF3 \u_decoder/fir_filter/I_data_add_7_buff_reg[13]  ( .D(n2623), .C(inClock), .Q(\u_decoder/fir_filter/I_data_add_7_buff [13]) );
  DF3 \u_decoder/fir_filter/I_data_add_7_buff_reg[12]  ( .D(n2624), .C(inClock), .Q(\u_decoder/fir_filter/I_data_add_7_buff [12]) );
  DF3 \u_decoder/fir_filter/I_data_add_7_buff_reg[11]  ( .D(n2625), .C(inClock), .Q(\u_decoder/fir_filter/I_data_add_7_buff [11]) );
  DF3 \u_decoder/fir_filter/I_data_add_7_buff_reg[10]  ( .D(n2626), .C(inClock), .Q(\u_decoder/fir_filter/I_data_add_7_buff [10]) );
  DF3 \u_decoder/fir_filter/I_data_add_7_buff_reg[9]  ( .D(n2627), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_7_buff [9]) );
  DF3 \u_decoder/fir_filter/I_data_add_7_buff_reg[8]  ( .D(n2628), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_7_buff [8]) );
  DF3 \u_decoder/fir_filter/I_data_add_7_buff_reg[7]  ( .D(n2629), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_7_buff [7]) );
  DF3 \u_decoder/fir_filter/I_data_add_7_buff_reg[6]  ( .D(n2630), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_7_buff [6]) );
  DF3 \u_decoder/fir_filter/I_data_add_7_buff_reg[5]  ( .D(n2631), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_7_buff [5]) );
  DF3 \u_decoder/fir_filter/I_data_add_7_buff_reg[4]  ( .D(n2632), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_7_buff [4]) );
  DF3 \u_decoder/fir_filter/I_data_add_7_buff_reg[3]  ( .D(n2633), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_7_buff [3]) );
  DF3 \u_decoder/fir_filter/I_data_add_7_buff_reg[2]  ( .D(n2634), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_7_buff [2]) );
  DF3 \u_decoder/fir_filter/I_data_add_7_buff_reg[1]  ( .D(n2635), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_7_buff [1]) );
  DF3 \u_decoder/fir_filter/I_data_add_7_buff_reg[0]  ( .D(n2636), .C(inClock), 
        .Q(\u_decoder/fir_filter/I_data_add_7_buff [0]), .QN(n108) );
  DF3 \u_decoder/fir_filter/I_data_mult_8_buff_reg[0]  ( .D(
        \u_decoder/fir_filter/n1303 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_8_buff [0]), .QN(n106) );
  DF3 \u_decoder/fir_filter/I_data_mult_8_buff_reg[1]  ( .D(
        \u_decoder/fir_filter/n1304 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_8_buff [1]) );
  DF3 \u_decoder/fir_filter/I_data_mult_8_buff_reg[2]  ( .D(
        \u_decoder/fir_filter/n1305 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_8_buff [2]) );
  DF3 \u_decoder/fir_filter/I_data_mult_8_buff_reg[3]  ( .D(
        \u_decoder/fir_filter/n1306 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_8_buff [3]) );
  DF3 \u_decoder/fir_filter/I_data_mult_8_buff_reg[4]  ( .D(
        \u_decoder/fir_filter/n1307 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_8_buff [4]) );
  DF3 \u_decoder/fir_filter/I_data_mult_8_buff_reg[5]  ( .D(
        \u_decoder/fir_filter/n1308 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_8_buff [5]) );
  DF3 \u_decoder/fir_filter/I_data_mult_8_buff_reg[6]  ( .D(
        \u_decoder/fir_filter/n1309 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_8_buff [6]) );
  DF3 \u_decoder/fir_filter/I_data_mult_8_buff_reg[7]  ( .D(
        \u_decoder/fir_filter/n1310 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_8_buff [7]) );
  DF3 \u_decoder/fir_filter/I_data_mult_8_buff_reg[8]  ( .D(
        \u_decoder/fir_filter/n1311 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_8_buff [8]) );
  DF3 \u_decoder/fir_filter/I_data_mult_8_buff_reg[9]  ( .D(
        \u_decoder/fir_filter/n1312 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_8_buff [9]) );
  DF3 \u_decoder/fir_filter/I_data_mult_8_buff_reg[10]  ( .D(
        \u_decoder/fir_filter/n1313 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_8_buff [10]) );
  DF3 \u_decoder/fir_filter/I_data_mult_8_buff_reg[11]  ( .D(
        \u_decoder/fir_filter/n1314 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_8_buff [11]) );
  DF3 \u_decoder/fir_filter/I_data_mult_8_buff_reg[12]  ( .D(
        \u_decoder/fir_filter/n1315 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_8_buff [12]) );
  DF3 \u_decoder/fir_filter/I_data_mult_8_buff_reg[13]  ( .D(
        \u_decoder/fir_filter/n1316 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_8_buff [13]) );
  DF3 \u_decoder/fir_filter/I_data_mult_8_buff_reg[14]  ( .D(
        \u_decoder/fir_filter/n1317 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_8_buff [14]) );
  DF3 \u_decoder/fir_filter/I_data_mult_8_delay_reg[0]  ( .D(
        \u_decoder/fir_filter/n1324 ), .C(inClock), .QN(
        \u_decoder/fir_filter/n426 ) );
  DF3 \u_decoder/fir_filter/I_data_mult_8_delay_reg[1]  ( .D(
        \u_decoder/fir_filter/n1325 ), .C(inClock), .QN(
        \u_decoder/fir_filter/n425 ) );
  DF3 \u_decoder/fir_filter/I_data_mult_8_delay_reg[2]  ( .D(
        \u_decoder/fir_filter/n1326 ), .C(inClock), .QN(
        \u_decoder/fir_filter/n424 ) );
  DF3 \u_decoder/fir_filter/I_data_mult_8_delay_reg[3]  ( .D(
        \u_decoder/fir_filter/n1327 ), .C(inClock), .QN(
        \u_decoder/fir_filter/n423 ) );
  DF3 \u_decoder/fir_filter/I_data_mult_8_delay_reg[4]  ( .D(
        \u_decoder/fir_filter/n1328 ), .C(inClock), .QN(
        \u_decoder/fir_filter/n422 ) );
  DF3 \u_decoder/fir_filter/I_data_mult_8_delay_reg[5]  ( .D(
        \u_decoder/fir_filter/n1329 ), .C(inClock), .QN(
        \u_decoder/fir_filter/n421 ) );
  DF3 \u_decoder/fir_filter/I_data_mult_8_delay_reg[6]  ( .D(
        \u_decoder/fir_filter/n1330 ), .C(inClock), .QN(
        \u_decoder/fir_filter/n420 ) );
  DF3 \u_decoder/fir_filter/I_data_mult_8_delay_reg[7]  ( .D(
        \u_decoder/fir_filter/n1331 ), .C(inClock), .QN(
        \u_decoder/fir_filter/n419 ) );
  DF3 \u_decoder/fir_filter/I_data_mult_8_delay_reg[8]  ( .D(
        \u_decoder/fir_filter/n1332 ), .C(inClock), .QN(
        \u_decoder/fir_filter/n418 ) );
  DF3 \u_decoder/fir_filter/I_data_mult_8_delay_reg[9]  ( .D(
        \u_decoder/fir_filter/n1333 ), .C(inClock), .QN(
        \u_decoder/fir_filter/n417 ) );
  DF3 \u_decoder/fir_filter/I_data_mult_8_delay_reg[10]  ( .D(
        \u_decoder/fir_filter/n1334 ), .C(inClock), .QN(
        \u_decoder/fir_filter/n416 ) );
  DF3 \u_decoder/fir_filter/I_data_mult_8_delay_reg[11]  ( .D(
        \u_decoder/fir_filter/n1335 ), .C(inClock), .QN(
        \u_decoder/fir_filter/n415 ) );
  DF3 \u_decoder/fir_filter/I_data_mult_8_delay_reg[12]  ( .D(
        \u_decoder/fir_filter/n1336 ), .C(inClock), .QN(
        \u_decoder/fir_filter/n414 ) );
  DF3 \u_decoder/fir_filter/I_data_mult_8_delay_reg[13]  ( .D(
        \u_decoder/fir_filter/n1337 ), .C(inClock), .QN(
        \u_decoder/fir_filter/n413 ) );
  DF3 \u_decoder/fir_filter/I_data_mult_8_delay_reg[14]  ( .D(
        \u_decoder/fir_filter/n1338 ), .C(inClock), .QN(
        \u_decoder/fir_filter/n412 ) );
  DF3 \u_decoder/fir_filter/I_data_mult_7_buff_reg[0]  ( .D(
        \u_decoder/fir_filter/n1340 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_7_buff [0]), .QN(n26) );
  DF3 \u_decoder/fir_filter/I_data_mult_7_buff_reg[1]  ( .D(
        \u_decoder/fir_filter/n1341 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_7_buff [1]) );
  DF3 \u_decoder/fir_filter/I_data_mult_7_buff_reg[2]  ( .D(
        \u_decoder/fir_filter/n1342 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_7_buff [2]) );
  DF3 \u_decoder/fir_filter/I_data_mult_7_buff_reg[3]  ( .D(
        \u_decoder/fir_filter/n1343 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_7_buff [3]) );
  DF3 \u_decoder/fir_filter/I_data_mult_7_buff_reg[4]  ( .D(
        \u_decoder/fir_filter/n1344 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_7_buff [4]) );
  DF3 \u_decoder/fir_filter/I_data_mult_7_buff_reg[5]  ( .D(
        \u_decoder/fir_filter/n1345 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_7_buff [5]) );
  DF3 \u_decoder/fir_filter/I_data_mult_7_buff_reg[6]  ( .D(
        \u_decoder/fir_filter/n1346 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_7_buff [6]) );
  DF3 \u_decoder/fir_filter/I_data_mult_7_buff_reg[7]  ( .D(
        \u_decoder/fir_filter/n1347 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_7_buff [7]) );
  DF3 \u_decoder/fir_filter/I_data_mult_7_buff_reg[8]  ( .D(
        \u_decoder/fir_filter/n1348 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_7_buff [8]) );
  DF3 \u_decoder/fir_filter/I_data_mult_7_buff_reg[9]  ( .D(
        \u_decoder/fir_filter/n1349 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_7_buff [9]) );
  DF3 \u_decoder/fir_filter/I_data_mult_7_buff_reg[10]  ( .D(
        \u_decoder/fir_filter/n1350 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_7_buff [10]) );
  DF3 \u_decoder/fir_filter/I_data_mult_7_buff_reg[11]  ( .D(
        \u_decoder/fir_filter/n1351 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_7_buff [11]) );
  DF3 \u_decoder/fir_filter/I_data_mult_7_buff_reg[12]  ( .D(
        \u_decoder/fir_filter/n1352 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_7_buff [12]) );
  DF3 \u_decoder/fir_filter/I_data_mult_7_buff_reg[13]  ( .D(
        \u_decoder/fir_filter/n1353 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_7_buff [13]) );
  DF3 \u_decoder/fir_filter/I_data_mult_7_buff_reg[14]  ( .D(
        \u_decoder/fir_filter/n1354 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_7_buff [14]) );
  DF3 \u_decoder/fir_filter/I_data_mult_6_buff_reg[0]  ( .D(n2637), .C(inClock), .Q(\u_decoder/fir_filter/I_data_mult_6_buff [0]), .QN(n27) );
  DF3 \u_decoder/fir_filter/I_data_mult_6_buff_reg[1]  ( .D(
        \u_decoder/fir_filter/n1357 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_6_buff [1]) );
  DF3 \u_decoder/fir_filter/I_data_mult_6_buff_reg[2]  ( .D(
        \u_decoder/fir_filter/n1358 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_6_buff [2]) );
  DF3 \u_decoder/fir_filter/I_data_mult_6_buff_reg[3]  ( .D(
        \u_decoder/fir_filter/n1359 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_6_buff [3]) );
  DF3 \u_decoder/fir_filter/I_data_mult_6_buff_reg[4]  ( .D(
        \u_decoder/fir_filter/n1360 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_6_buff [4]) );
  DF3 \u_decoder/fir_filter/I_data_mult_6_buff_reg[5]  ( .D(
        \u_decoder/fir_filter/n1361 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_6_buff [5]) );
  DF3 \u_decoder/fir_filter/I_data_mult_6_buff_reg[6]  ( .D(
        \u_decoder/fir_filter/n1362 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_6_buff [6]) );
  DF3 \u_decoder/fir_filter/I_data_mult_6_buff_reg[7]  ( .D(
        \u_decoder/fir_filter/n1363 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_6_buff [7]) );
  DF3 \u_decoder/fir_filter/I_data_mult_6_buff_reg[8]  ( .D(
        \u_decoder/fir_filter/n1364 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_6_buff [8]) );
  DF3 \u_decoder/fir_filter/I_data_mult_6_buff_reg[9]  ( .D(
        \u_decoder/fir_filter/n1365 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_6_buff [9]) );
  DF3 \u_decoder/fir_filter/I_data_mult_6_buff_reg[10]  ( .D(
        \u_decoder/fir_filter/n1366 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_6_buff [10]) );
  DF3 \u_decoder/fir_filter/I_data_mult_6_buff_reg[11]  ( .D(
        \u_decoder/fir_filter/n1367 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_6_buff [11]) );
  DF3 \u_decoder/fir_filter/I_data_mult_6_buff_reg[12]  ( .D(
        \u_decoder/fir_filter/n1368 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_6_buff [12]) );
  DF3 \u_decoder/fir_filter/I_data_mult_6_buff_reg[13]  ( .D(
        \u_decoder/fir_filter/n1369 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_6_buff [13]) );
  DF3 \u_decoder/fir_filter/I_data_mult_6_buff_reg[14]  ( .D(
        \u_decoder/fir_filter/n1370 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_6_buff [14]) );
  DF3 \u_decoder/fir_filter/I_data_mult_5_buff_reg[0]  ( .D(
        \u_decoder/fir_filter/n1372 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_5_buff [0]), .QN(n28) );
  DF3 \u_decoder/fir_filter/I_data_mult_5_buff_reg[1]  ( .D(
        \u_decoder/fir_filter/n1373 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_5_buff [1]) );
  DF3 \u_decoder/fir_filter/I_data_mult_5_buff_reg[2]  ( .D(
        \u_decoder/fir_filter/n1374 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_5_buff [2]) );
  DF3 \u_decoder/fir_filter/I_data_mult_5_buff_reg[3]  ( .D(
        \u_decoder/fir_filter/n1375 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_5_buff [3]) );
  DF3 \u_decoder/fir_filter/I_data_mult_5_buff_reg[4]  ( .D(
        \u_decoder/fir_filter/n1376 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_5_buff [4]) );
  DF3 \u_decoder/fir_filter/I_data_mult_5_buff_reg[5]  ( .D(
        \u_decoder/fir_filter/n1377 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_5_buff [5]) );
  DF3 \u_decoder/fir_filter/I_data_mult_5_buff_reg[6]  ( .D(
        \u_decoder/fir_filter/n1378 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_5_buff [6]) );
  DF3 \u_decoder/fir_filter/I_data_mult_5_buff_reg[7]  ( .D(
        \u_decoder/fir_filter/n1379 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_5_buff [7]) );
  DF3 \u_decoder/fir_filter/I_data_mult_5_buff_reg[8]  ( .D(
        \u_decoder/fir_filter/n1380 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_5_buff [8]) );
  DF3 \u_decoder/fir_filter/I_data_mult_5_buff_reg[9]  ( .D(
        \u_decoder/fir_filter/n1381 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_5_buff [9]) );
  DF3 \u_decoder/fir_filter/I_data_mult_5_buff_reg[10]  ( .D(
        \u_decoder/fir_filter/n1382 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_5_buff [10]) );
  DF3 \u_decoder/fir_filter/I_data_mult_5_buff_reg[11]  ( .D(
        \u_decoder/fir_filter/n1383 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_5_buff [11]) );
  DF3 \u_decoder/fir_filter/I_data_mult_5_buff_reg[12]  ( .D(
        \u_decoder/fir_filter/n1384 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_5_buff [12]) );
  DF3 \u_decoder/fir_filter/I_data_mult_5_buff_reg[13]  ( .D(
        \u_decoder/fir_filter/n1385 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_5_buff [13]) );
  DF3 \u_decoder/fir_filter/I_data_mult_5_buff_reg[14]  ( .D(
        \u_decoder/fir_filter/n1386 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_5_buff [14]) );
  DF3 \u_decoder/fir_filter/I_data_mult_4_buff_reg[0]  ( .D(n2255), .C(inClock), .Q(\u_decoder/fir_filter/I_data_mult_4_buff [0]), .QN(n38) );
  DF3 \u_decoder/fir_filter/I_data_mult_4_buff_reg[1]  ( .D(n2298), .C(inClock), .Q(\u_decoder/fir_filter/I_data_mult_4_buff [1]) );
  DF3 \u_decoder/fir_filter/I_data_mult_4_buff_reg[2]  ( .D(n2300), .C(inClock), .Q(\u_decoder/fir_filter/I_data_mult_4_buff [2]) );
  DF3 \u_decoder/fir_filter/I_data_mult_4_buff_reg[3]  ( .D(n2273), .C(inClock), .Q(\u_decoder/fir_filter/I_data_mult_4_buff [3]) );
  DF3 \u_decoder/fir_filter/I_data_mult_4_buff_reg[4]  ( .D(n2272), .C(inClock), .Q(\u_decoder/fir_filter/I_data_mult_4_buff [4]) );
  DF3 \u_decoder/fir_filter/I_data_mult_4_buff_reg[5]  ( .D(n2271), .C(inClock), .Q(\u_decoder/fir_filter/I_data_mult_4_buff [5]) );
  DF3 \u_decoder/fir_filter/I_data_mult_4_buff_reg[6]  ( .D(n2270), .C(inClock), .Q(\u_decoder/fir_filter/I_data_mult_4_buff [6]) );
  DF3 \u_decoder/fir_filter/I_data_mult_4_buff_reg[7]  ( .D(n2269), .C(inClock), .Q(\u_decoder/fir_filter/I_data_mult_4_buff [7]) );
  DF3 \u_decoder/fir_filter/I_data_mult_4_buff_reg[8]  ( .D(n2268), .C(inClock), .Q(\u_decoder/fir_filter/I_data_mult_4_buff [8]) );
  DF3 \u_decoder/fir_filter/I_data_mult_4_buff_reg[9]  ( .D(n2267), .C(inClock), .Q(\u_decoder/fir_filter/I_data_mult_4_buff [9]) );
  DF3 \u_decoder/fir_filter/I_data_mult_4_buff_reg[10]  ( .D(n2265), .C(
        inClock), .Q(\u_decoder/fir_filter/I_data_mult_4_buff [10]) );
  DF3 \u_decoder/fir_filter/I_data_mult_4_buff_reg[11]  ( .D(n2261), .C(
        inClock), .Q(\u_decoder/fir_filter/I_data_mult_4_buff [11]) );
  DF3 \u_decoder/fir_filter/I_data_mult_4_buff_reg[12]  ( .D(n2256), .C(
        inClock), .Q(\u_decoder/fir_filter/I_data_mult_4_buff [12]) );
  DF3 \u_decoder/fir_filter/I_data_mult_4_buff_reg[13]  ( .D(n2258), .C(
        inClock), .Q(\u_decoder/fir_filter/I_data_mult_4_buff [13]) );
  DF3 \u_decoder/fir_filter/I_data_mult_4_buff_reg[14]  ( .D(n2259), .C(
        inClock), .Q(\u_decoder/fir_filter/I_data_mult_4_buff [14]) );
  DF3 \u_decoder/fir_filter/I_data_mult_3_buff_reg[0]  ( .D(
        \u_decoder/fir_filter/n1388 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_3_buff [0]), .QN(n29) );
  DF3 \u_decoder/fir_filter/I_data_mult_3_buff_reg[1]  ( .D(
        \u_decoder/fir_filter/n1389 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_3_buff [1]) );
  DF3 \u_decoder/fir_filter/I_data_mult_3_buff_reg[2]  ( .D(
        \u_decoder/fir_filter/n1390 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_3_buff [2]) );
  DF3 \u_decoder/fir_filter/I_data_mult_3_buff_reg[3]  ( .D(
        \u_decoder/fir_filter/n1391 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_3_buff [3]) );
  DF3 \u_decoder/fir_filter/I_data_mult_3_buff_reg[4]  ( .D(
        \u_decoder/fir_filter/n1392 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_3_buff [4]) );
  DF3 \u_decoder/fir_filter/I_data_mult_3_buff_reg[5]  ( .D(
        \u_decoder/fir_filter/n1393 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_3_buff [5]) );
  DF3 \u_decoder/fir_filter/I_data_mult_3_buff_reg[6]  ( .D(
        \u_decoder/fir_filter/n1394 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_3_buff [6]) );
  DF3 \u_decoder/fir_filter/I_data_mult_3_buff_reg[7]  ( .D(
        \u_decoder/fir_filter/n1395 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_3_buff [7]) );
  DF3 \u_decoder/fir_filter/I_data_mult_3_buff_reg[8]  ( .D(
        \u_decoder/fir_filter/n1396 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_3_buff [8]) );
  DF3 \u_decoder/fir_filter/I_data_mult_3_buff_reg[9]  ( .D(
        \u_decoder/fir_filter/n1397 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_3_buff [9]) );
  DF3 \u_decoder/fir_filter/I_data_mult_3_buff_reg[10]  ( .D(
        \u_decoder/fir_filter/n1398 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_3_buff [10]) );
  DF3 \u_decoder/fir_filter/I_data_mult_3_buff_reg[11]  ( .D(
        \u_decoder/fir_filter/n1399 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_3_buff [11]) );
  DF3 \u_decoder/fir_filter/I_data_mult_3_buff_reg[12]  ( .D(
        \u_decoder/fir_filter/n1400 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_3_buff [12]) );
  DF3 \u_decoder/fir_filter/I_data_mult_3_buff_reg[13]  ( .D(
        \u_decoder/fir_filter/n1401 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_3_buff [13]) );
  DF3 \u_decoder/fir_filter/I_data_mult_3_buff_reg[14]  ( .D(
        \u_decoder/fir_filter/n1402 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_3_buff [14]) );
  DF3 \u_decoder/fir_filter/I_data_mult_2_buff_reg[0]  ( .D(n2638), .C(inClock), .Q(\u_decoder/fir_filter/I_data_mult_2_buff [0]), .QN(n30) );
  DF3 \u_decoder/fir_filter/I_data_mult_2_buff_reg[1]  ( .D(
        \u_decoder/fir_filter/n1405 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_2_buff [1]) );
  DF3 \u_decoder/fir_filter/I_data_mult_2_buff_reg[2]  ( .D(
        \u_decoder/fir_filter/n1406 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_2_buff [2]) );
  DF3 \u_decoder/fir_filter/I_data_mult_2_buff_reg[3]  ( .D(
        \u_decoder/fir_filter/n1407 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_2_buff [3]) );
  DF3 \u_decoder/fir_filter/I_data_mult_2_buff_reg[4]  ( .D(
        \u_decoder/fir_filter/n1408 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_2_buff [4]) );
  DF3 \u_decoder/fir_filter/I_data_mult_2_buff_reg[5]  ( .D(
        \u_decoder/fir_filter/n1409 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_2_buff [5]) );
  DF3 \u_decoder/fir_filter/I_data_mult_2_buff_reg[6]  ( .D(
        \u_decoder/fir_filter/n1410 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_2_buff [6]) );
  DF3 \u_decoder/fir_filter/I_data_mult_2_buff_reg[7]  ( .D(
        \u_decoder/fir_filter/n1411 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_2_buff [7]) );
  DF3 \u_decoder/fir_filter/I_data_mult_2_buff_reg[8]  ( .D(
        \u_decoder/fir_filter/n1412 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_2_buff [8]) );
  DF3 \u_decoder/fir_filter/I_data_mult_2_buff_reg[9]  ( .D(
        \u_decoder/fir_filter/n1413 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_2_buff [9]) );
  DF3 \u_decoder/fir_filter/I_data_mult_2_buff_reg[10]  ( .D(
        \u_decoder/fir_filter/n1414 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_2_buff [10]) );
  DF3 \u_decoder/fir_filter/I_data_mult_2_buff_reg[11]  ( .D(
        \u_decoder/fir_filter/n1415 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_2_buff [11]) );
  DF3 \u_decoder/fir_filter/I_data_mult_2_buff_reg[12]  ( .D(
        \u_decoder/fir_filter/n1416 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_2_buff [12]) );
  DF3 \u_decoder/fir_filter/I_data_mult_2_buff_reg[13]  ( .D(
        \u_decoder/fir_filter/n1417 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_2_buff [13]) );
  DF3 \u_decoder/fir_filter/I_data_mult_2_buff_reg[14]  ( .D(
        \u_decoder/fir_filter/n1418 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_2_buff [14]) );
  DF3 \u_decoder/fir_filter/I_data_mult_1_buff_reg[0]  ( .D(
        \u_decoder/fir_filter/n1420 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_1_buff [0]), .QN(n31) );
  DF3 \u_decoder/fir_filter/I_data_mult_1_buff_reg[1]  ( .D(
        \u_decoder/fir_filter/n1421 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_1_buff [1]) );
  DF3 \u_decoder/fir_filter/I_data_mult_1_buff_reg[2]  ( .D(
        \u_decoder/fir_filter/n1422 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_1_buff [2]) );
  DF3 \u_decoder/fir_filter/I_data_mult_1_buff_reg[3]  ( .D(
        \u_decoder/fir_filter/n1423 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_1_buff [3]) );
  DF3 \u_decoder/fir_filter/I_data_mult_1_buff_reg[4]  ( .D(
        \u_decoder/fir_filter/n1424 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_1_buff [4]) );
  DF3 \u_decoder/fir_filter/I_data_mult_1_buff_reg[5]  ( .D(
        \u_decoder/fir_filter/n1425 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_1_buff [5]) );
  DF3 \u_decoder/fir_filter/I_data_mult_1_buff_reg[6]  ( .D(
        \u_decoder/fir_filter/n1426 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_1_buff [6]) );
  DF3 \u_decoder/fir_filter/I_data_mult_1_buff_reg[7]  ( .D(
        \u_decoder/fir_filter/n1427 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_1_buff [7]) );
  DF3 \u_decoder/fir_filter/I_data_mult_1_buff_reg[8]  ( .D(
        \u_decoder/fir_filter/n1428 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_1_buff [8]) );
  DF3 \u_decoder/fir_filter/I_data_mult_1_buff_reg[9]  ( .D(
        \u_decoder/fir_filter/n1429 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_1_buff [9]) );
  DF3 \u_decoder/fir_filter/I_data_mult_1_buff_reg[10]  ( .D(
        \u_decoder/fir_filter/n1430 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_1_buff [10]) );
  DF3 \u_decoder/fir_filter/I_data_mult_1_buff_reg[11]  ( .D(
        \u_decoder/fir_filter/n1431 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_1_buff [11]) );
  DF3 \u_decoder/fir_filter/I_data_mult_1_buff_reg[12]  ( .D(
        \u_decoder/fir_filter/n1432 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_1_buff [12]) );
  DF3 \u_decoder/fir_filter/I_data_mult_1_buff_reg[13]  ( .D(
        \u_decoder/fir_filter/n1433 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_1_buff [13]) );
  DF3 \u_decoder/fir_filter/I_data_mult_1_buff_reg[14]  ( .D(
        \u_decoder/fir_filter/n1434 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_1_buff [14]) );
  DF3 \u_decoder/fir_filter/I_data_mult_0_buff_reg[0]  ( .D(
        \u_decoder/fir_filter/n1436 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_0_buff [0]) );
  DF3 \u_decoder/fir_filter/I_data_mult_0_buff_reg[1]  ( .D(
        \u_decoder/fir_filter/n1437 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_0_buff [1]), .QN(n94) );
  DF3 \u_decoder/fir_filter/I_data_mult_0_buff_reg[2]  ( .D(
        \u_decoder/fir_filter/n1438 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_0_buff [2]), .QN(n92) );
  DF3 \u_decoder/fir_filter/I_data_mult_0_buff_reg[3]  ( .D(
        \u_decoder/fir_filter/n1439 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_0_buff [3]), .QN(n138) );
  DF3 \u_decoder/fir_filter/I_data_mult_0_buff_reg[4]  ( .D(
        \u_decoder/fir_filter/n1440 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_0_buff [4]), .QN(n139) );
  DF3 \u_decoder/fir_filter/I_data_mult_0_buff_reg[5]  ( .D(
        \u_decoder/fir_filter/n1441 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_0_buff [5]), .QN(n140) );
  DF3 \u_decoder/fir_filter/I_data_mult_0_buff_reg[6]  ( .D(
        \u_decoder/fir_filter/n1442 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_0_buff [6]), .QN(n178) );
  DF3 \u_decoder/fir_filter/I_data_mult_0_buff_reg[7]  ( .D(
        \u_decoder/fir_filter/n1443 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_0_buff [7]) );
  DF3 \u_decoder/fir_filter/I_data_mult_0_buff_reg[8]  ( .D(
        \u_decoder/fir_filter/n1444 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_0_buff [8]), .QN(n224) );
  DF3 \u_decoder/fir_filter/I_data_mult_0_buff_reg[9]  ( .D(
        \u_decoder/fir_filter/n1445 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_0_buff [9]) );
  DF3 \u_decoder/fir_filter/I_data_mult_0_buff_reg[10]  ( .D(
        \u_decoder/fir_filter/n1446 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_0_buff [10]), .QN(n265) );
  DF3 \u_decoder/fir_filter/I_data_mult_0_buff_reg[11]  ( .D(
        \u_decoder/fir_filter/n1447 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_0_buff [11]) );
  DF3 \u_decoder/fir_filter/I_data_mult_0_buff_reg[12]  ( .D(
        \u_decoder/fir_filter/n1448 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_0_buff [12]) );
  DF3 \u_decoder/fir_filter/I_data_mult_0_buff_reg[13]  ( .D(
        \u_decoder/fir_filter/n1449 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_0_buff [13]) );
  DF3 \u_decoder/fir_filter/I_data_mult_0_buff_reg[14]  ( .D(
        \u_decoder/fir_filter/n1450 ), .C(inClock), .Q(
        \u_decoder/fir_filter/I_data_mult_0_buff [14]) );
  DF3 \u_decoder/fir_filter/o_postfilter_ready_reg  ( .D(
        \u_decoder/fir_filter/n1451 ), .C(inClock), .Q(\sig_MUX_inMUX8[0] ) );
  DF3 \u_decoder/fir_filter/state_reg[0]  ( .D(\u_decoder/fir_filter/N11 ), 
        .C(inClock), .Q(\u_decoder/fir_filter/state [0]), .QN(
        \u_decoder/fir_filter/n410 ) );
  DF3 \u_decoder/fir_filter/state_reg[1]  ( .D(\u_decoder/fir_filter/N12 ), 
        .C(inClock), .Q(\u_decoder/fir_filter/state [1]) );
  DF3 \u_cordic/mycordic/o_angle_reg[15]  ( .D(n1868), .C(inClock), .Q(
        \u_cordic/cordic_to_rotation [15]) );
  DF3 \u_cordic/mycordic/o_angle_reg[14]  ( .D(n1869), .C(inClock), .Q(
        \u_cordic/cordic_to_rotation [14]) );
  DF3 \u_cordic/mycordic/o_angle_reg[13]  ( .D(n1870), .C(inClock), .Q(
        \u_cordic/cordic_to_rotation [13]) );
  DF3 \u_cordic/mycordic/o_angle_reg[12]  ( .D(n1871), .C(inClock), .Q(
        \u_cordic/cordic_to_rotation [12]) );
  DF3 \u_cordic/mycordic/o_angle_reg[11]  ( .D(n1872), .C(inClock), .Q(
        \u_cordic/cordic_to_rotation [11]) );
  DF3 \u_cordic/mycordic/o_angle_reg[10]  ( .D(n1873), .C(inClock), .Q(
        \u_cordic/cordic_to_rotation [10]) );
  DF3 \u_cordic/mycordic/o_angle_reg[9]  ( .D(n1874), .C(inClock), .Q(
        \u_cordic/cordic_to_rotation [9]) );
  DF3 \u_cordic/mycordic/o_angle_reg[8]  ( .D(n1875), .C(inClock), .Q(
        \u_cordic/cordic_to_rotation [8]) );
  DF3 \u_cordic/mycordic/o_angle_reg[7]  ( .D(n1876), .C(inClock), .Q(
        \u_cordic/cordic_to_rotation [7]) );
  DF3 \u_cordic/mycordic/o_angle_reg[6]  ( .D(n1877), .C(inClock), .Q(
        \u_cordic/cordic_to_rotation [6]) );
  DF3 \u_cordic/mycordic/o_angle_reg[5]  ( .D(n1878), .C(inClock), .Q(
        \u_cordic/cordic_to_rotation [5]) );
  DF3 \u_cordic/mycordic/o_angle_reg[4]  ( .D(n1879), .C(inClock), .Q(
        \u_cordic/cordic_to_rotation [4]) );
  DF3 \u_cordic/mycordic/o_angle_reg[3]  ( .D(n1880), .C(inClock), .Q(
        \u_cordic/cordic_to_rotation [3]) );
  DF3 \u_cordic/mycordic/o_angle_reg[2]  ( .D(n1882), .C(inClock), .Q(
        \u_cordic/cordic_to_rotation [2]) );
  DF3 \u_cordic/mycordic/o_angle_reg[1]  ( .D(n1893), .C(inClock), .Q(
        \u_cordic/cordic_to_rotation [1]) );
  DF3 \u_cordic/mycordic/o_angle_reg[0]  ( .D(n1902), .C(inClock), .Q(
        \u_cordic/cordic_to_rotation [0]) );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[6][15]  ( .D(n1452), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[6][15] ) );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[6][14]  ( .D(n1451), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[6][14] ), .QN(n268) );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[6][13]  ( .D(n1450), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[6][13] ), .QN(n267) );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[6][12]  ( .D(n1449), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[6][12] ), .QN(n266) );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[6][11]  ( .D(n1448), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[6][11] ), .QN(n229) );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[6][10]  ( .D(n1447), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[6][10] ), .QN(n228) );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[6][9]  ( .D(n1446), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[6][9] ), .QN(n181)
         );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[6][8]  ( .D(n1445), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[6][8] ), .QN(n182)
         );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[6][7]  ( .D(n1444), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[6][7] ), .QN(n389)
         );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[6][6]  ( .D(n1443), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[6][6] ), .QN(n141)
         );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[6][5]  ( .D(n1442), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[6][5] ), .QN(n391)
         );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[6][4]  ( .D(n1441), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[6][4] ), .QN(n387)
         );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[6][3]  ( .D(n1440), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[6][3] ), .QN(n305)
         );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[6][2]  ( .D(n1439), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[6][2] ), .QN(n96)
         );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[6][1]  ( .D(n1438), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[6][1] ), .QN(n314)
         );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[6][0]  ( .D(n1437), .C(
        inClock), .Q(\u_cordic/mycordic/N615 ), .QN(n313) );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[5][15]  ( .D(n1512), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[5][15] ) );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[5][14]  ( .D(n1511), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[5][14] ), .QN(n312) );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[5][13]  ( .D(n1510), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[5][13] ), .QN(n283) );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[5][12]  ( .D(n1509), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[5][12] ), .QN(n282) );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[5][11]  ( .D(n1508), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[5][11] ), .QN(n281) );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[5][10]  ( .D(n1507), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[5][10] ), .QN(n244) );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[5][9]  ( .D(n1506), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[5][9] ), .QN(n243)
         );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[5][8]  ( .D(n1505), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[5][8] ), .QN(n192)
         );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[5][7]  ( .D(n1504), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[5][7] ), .QN(n191)
         );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[5][6]  ( .D(n1503), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[5][6] ), .QN(n160)
         );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[5][5]  ( .D(n1502), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[5][5] ), .QN(n159)
         );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[5][4]  ( .D(n1501), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[5][4] ), .QN(n158)
         );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[5][3]  ( .D(n1500), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[5][3] ), .QN(n105)
         );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[5][2]  ( .D(n1499), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[5][2] ), .QN(n104)
         );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[5][1]  ( .D(n1498), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[5][1] ), .QN(n296)
         );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[5][0]  ( .D(n1497), .C(
        inClock), .Q(\u_cordic/mycordic/N550 ) );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[4][15]  ( .D(n1536), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[4][15] ) );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[4][14]  ( .D(n1535), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[4][14] ), .QN(n311) );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[4][13]  ( .D(n1534), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[4][13] ), .QN(n280) );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[4][12]  ( .D(n1533), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[4][12] ), .QN(n279) );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[4][11]  ( .D(n1532), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[4][11] ), .QN(n278) );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[4][10]  ( .D(n1531), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[4][10] ), .QN(n242) );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[4][9]  ( .D(n1530), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[4][9] ), .QN(n241)
         );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[4][8]  ( .D(n1529), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[4][8] ), .QN(n190)
         );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[4][7]  ( .D(n1528), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[4][7] ), .QN(n189)
         );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[4][6]  ( .D(n1527), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[4][6] ), .QN(n157)
         );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[4][5]  ( .D(n1526), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[4][5] ), .QN(n156)
         );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[4][4]  ( .D(n1525), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[4][4] ), .QN(n155)
         );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[4][3]  ( .D(n1524), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[4][3] ), .QN(n103)
         );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[4][2]  ( .D(n1523), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[4][2] ), .QN(n102)
         );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[4][1]  ( .D(n1522), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[4][1] ), .QN(n99)
         );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[4][0]  ( .D(n1521), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[4][0] ), .QN(n299)
         );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[3][15]  ( .D(n1561), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[3][15] ) );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[3][14]  ( .D(n1560), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[3][14] ), .QN(n310) );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[3][13]  ( .D(n1559), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[3][13] ), .QN(n277) );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[3][12]  ( .D(n1558), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[3][12] ), .QN(n276) );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[3][11]  ( .D(n1557), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[3][11] ), .QN(n275) );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[3][10]  ( .D(n1556), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[3][10] ), .QN(n240) );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[3][9]  ( .D(n1555), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[3][9] ), .QN(n239)
         );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[3][8]  ( .D(n1554), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[3][8] ), .QN(n188)
         );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[3][7]  ( .D(n1553), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[3][7] ), .QN(n187)
         );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[3][6]  ( .D(n1552), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[3][6] ), .QN(n154)
         );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[3][5]  ( .D(n1551), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[3][5] ), .QN(n153)
         );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[3][4]  ( .D(n1550), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[3][4] ), .QN(n152)
         );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[3][3]  ( .D(n1549), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[3][3] ), .QN(n101)
         );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[3][2]  ( .D(n1548), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[3][2] ), .QN(n144)
         );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[3][1]  ( .D(n1547), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[3][1] ), .QN(n100)
         );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[3][0]  ( .D(n1546), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[3][0] ), .QN(n295)
         );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[2][15]  ( .D(n1468), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[2][15] ) );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[2][14]  ( .D(n1467), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[2][14] ), .QN(n309) );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[2][13]  ( .D(n1466), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[2][13] ), .QN(n274) );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[2][12]  ( .D(n1465), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[2][12] ), .QN(n273) );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[2][11]  ( .D(n1464), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[2][11] ), .QN(n272) );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[2][10]  ( .D(n1463), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[2][10] ), .QN(n238) );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[2][9]  ( .D(n1462), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[2][9] ), .QN(n237)
         );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[2][8]  ( .D(n1461), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[2][8] ), .QN(n186)
         );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[2][7]  ( .D(n1460), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[2][7] ), .QN(n185)
         );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[2][6]  ( .D(n1459), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[2][6] ), .QN(n151)
         );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[2][5]  ( .D(n1458), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[2][5] ), .QN(n150)
         );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[2][4]  ( .D(n1457), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[2][4] ), .QN(n149)
         );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[2][3]  ( .D(n1456), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[2][3] ), .QN(n143)
         );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[2][2]  ( .D(n1455), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[2][2] ), .QN(n148)
         );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[2][1]  ( .D(n1454), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[2][1] ), .QN(n298)
         );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[2][0]  ( .D(n1453), .C(
        inClock), .Q(\u_cordic/mycordic/N428 ) );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[1][15]  ( .D(n1905), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[1][15] ) );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[1][14]  ( .D(n1905), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[1][14] ), .QN(n308) );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[1][13]  ( .D(n1905), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[1][13] ), .QN(n271) );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[1][12]  ( .D(n1905), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[1][12] ), .QN(n270) );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[1][11]  ( .D(n1905), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[1][11] ), .QN(n269) );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[1][10]  ( .D(n1905), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[1][10] ), .QN(n236) );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[1][9]  ( .D(n1905), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[1][9] ), .QN(n235)
         );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[1][8]  ( .D(n1905), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[1][8] ), .QN(n184)
         );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[1][7]  ( .D(n1905), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[1][7] ), .QN(n183)
         );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[1][6]  ( .D(n1905), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[1][6] ), .QN(n147)
         );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[1][5]  ( .D(n774), .C(inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[1][5] ), .QN(n146) );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[1][4]  ( .D(n1905), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[1][4] ), .QN(n142)
         );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[1][3]  ( .D(n774), .C(inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[1][3] ), .QN(n145) );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[1][2]  ( .D(n774), .C(inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[1][2] ), .QN(n98) );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[1][1]  ( .D(n1905), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[1][1] ), .QN(n97)
         );
  DF3 \u_cordic/mycordic/present_ANGLE_table_reg[1][0]  ( .D(n1485), .C(
        inClock), .Q(\u_cordic/mycordic/present_ANGLE_table[1][0] ), .QN(n297)
         );
  DF3 \u_cordic/mycordic/present_C_table_reg[7][0]  ( .D(n1884), .C(inClock), 
        .Q(\u_cordic/mycordic/present_C_table[7][0] ) );
  DF3 \u_cordic/mycordic/present_C_table_reg[6][0]  ( .D(n1887), .C(inClock), 
        .Q(\u_cordic/mycordic/present_C_table[6][0] ) );
  DF3 \u_cordic/mycordic/present_C_table_reg[5][0]  ( .D(n1890), .C(inClock), 
        .Q(\u_cordic/mycordic/present_C_table[5][0] ) );
  DF3 \u_cordic/mycordic/present_C_table_reg[4][0]  ( .D(n1894), .C(inClock), 
        .Q(\u_cordic/mycordic/present_C_table[4][0] ) );
  DF3 \u_cordic/mycordic/present_C_table_reg[3][0]  ( .D(n1897), .C(inClock), 
        .Q(\u_cordic/mycordic/present_C_table[3][0] ) );
  DF3 \u_cordic/mycordic/present_C_table_reg[2][0]  ( .D(n1900), .C(inClock), 
        .Q(\u_cordic/mycordic/present_C_table[2][0] ) );
  DF3 \u_cordic/mycordic/present_C_table_reg[1][0]  ( .D(n1427), .C(inClock), 
        .Q(\u_cordic/mycordic/present_C_table[1][0] ) );
  DF3 \u_cordic/mycordic/present_C_table_reg[7][1]  ( .D(n1883), .C(inClock), 
        .Q(\u_cordic/mycordic/present_C_table[7][1] ), .QN(
        \u_cordic/mycordic/n110 ) );
  DF3 \u_cordic/mycordic/present_C_table_reg[6][1]  ( .D(n1886), .C(inClock), 
        .Q(\u_cordic/mycordic/present_C_table[6][1] ) );
  DF3 \u_cordic/mycordic/present_C_table_reg[5][1]  ( .D(n1889), .C(inClock), 
        .Q(\u_cordic/mycordic/present_C_table[5][1] ) );
  DF3 \u_cordic/mycordic/present_C_table_reg[4][1]  ( .D(n1892), .C(inClock), 
        .Q(\u_cordic/mycordic/present_C_table[4][1] ) );
  DF3 \u_cordic/mycordic/present_C_table_reg[3][1]  ( .D(n1896), .C(inClock), 
        .Q(\u_cordic/mycordic/present_C_table[3][1] ) );
  DF3 \u_cordic/mycordic/present_C_table_reg[2][1]  ( .D(n1899), .C(inClock), 
        .Q(\u_cordic/mycordic/present_C_table[2][1] ) );
  DF3 \u_cordic/mycordic/present_C_table_reg[1][1]  ( .D(
        \u_cordic/mycordic/N211 ), .C(inClock), .Q(
        \u_cordic/mycordic/present_C_table[1][1] ) );
  DF3 \u_cordic/mycordic/present_C_table_reg[7][2]  ( .D(n1881), .C(inClock), 
        .QN(\u_cordic/mycordic/n108 ) );
  DF3 \u_cordic/mycordic/present_C_table_reg[6][2]  ( .D(n1885), .C(inClock), 
        .Q(\u_cordic/mycordic/present_C_table[6][2] ) );
  DF3 \u_cordic/mycordic/present_C_table_reg[5][2]  ( .D(n1888), .C(inClock), 
        .Q(\u_cordic/mycordic/present_C_table[5][2] ) );
  DF3 \u_cordic/mycordic/present_C_table_reg[4][2]  ( .D(n1891), .C(inClock), 
        .Q(\u_cordic/mycordic/present_C_table[4][2] ) );
  DF3 \u_cordic/mycordic/present_C_table_reg[3][2]  ( .D(n1895), .C(inClock), 
        .Q(\u_cordic/mycordic/present_C_table[3][2] ) );
  DF3 \u_cordic/mycordic/present_C_table_reg[2][2]  ( .D(n1898), .C(inClock), 
        .Q(\u_cordic/mycordic/present_C_table[2][2] ) );
  DF3 \u_cordic/mycordic/present_C_table_reg[1][2]  ( .D(
        \u_cordic/mycordic/N212 ), .C(inClock), .Q(
        \u_cordic/mycordic/present_C_table[1][2] ) );
  DF3 \u_cordic/mycordic/present_Q_table_reg[6][7]  ( .D(n1496), .C(inClock), 
        .Q(\u_cordic/mycordic/present_Q_table[6][7] ) );
  DF3 \u_cordic/mycordic/present_Q_table_reg[5][7]  ( .D(n1520), .C(inClock), 
        .Q(\u_cordic/mycordic/present_Q_table[5][7] ) );
  DF3 \u_cordic/mycordic/present_Q_table_reg[5][6]  ( .D(n1519), .C(inClock), 
        .Q(\u_cordic/mycordic/present_Q_table[5][6] ), .QN(n286) );
  DF3 \u_cordic/mycordic/present_Q_table_reg[5][5]  ( .D(n1518), .C(inClock), 
        .Q(\u_cordic/mycordic/present_Q_table[5][5] ) );
  DF3 \u_cordic/mycordic/present_Q_table_reg[5][4]  ( .D(n1517), .C(inClock), 
        .Q(\u_cordic/mycordic/present_Q_table[5][4] ), .QN(n247) );
  DF3 \u_cordic/mycordic/present_Q_table_reg[5][3]  ( .D(n1516), .C(inClock), 
        .Q(\u_cordic/mycordic/present_Q_table[5][3] ) );
  DF3 \u_cordic/mycordic/present_Q_table_reg[5][2]  ( .D(n1515), .C(inClock), 
        .Q(\u_cordic/mycordic/present_Q_table[5][2] ), .QN(n197) );
  DF3 \u_cordic/mycordic/present_Q_table_reg[5][1]  ( .D(n1514), .C(inClock), 
        .Q(\u_cordic/mycordic/present_Q_table[5][1] ), .QN(n225) );
  DF3 \u_cordic/mycordic/present_Q_table_reg[5][0]  ( .D(n1513), .C(inClock), 
        .Q(\u_cordic/mycordic/present_Q_table[5][0] ), .QN(n180) );
  DF3 \u_cordic/mycordic/present_I_table_reg[5][7]  ( .D(n1540), .C(inClock), 
        .Q(\u_cordic/mycordic/present_I_table[5][7] ), .QN(n199) );
  DF3 \u_cordic/mycordic/present_I_table_reg[5][6]  ( .D(n1539), .C(inClock), 
        .Q(\u_cordic/mycordic/present_I_table[5][6] ) );
  DF3 \u_cordic/mycordic/present_I_table_reg[5][5]  ( .D(n1538), .C(inClock), 
        .Q(\u_cordic/mycordic/present_I_table[5][5] ), .QN(n46) );
  DF3 \u_cordic/mycordic/present_I_table_reg[5][4]  ( .D(n1537), .C(inClock), 
        .Q(\u_cordic/mycordic/present_I_table[5][4] ) );
  DF3 \u_cordic/mycordic/present_Q_table_reg[4][3]  ( .D(n1541), .C(inClock), 
        .Q(\u_cordic/mycordic/present_Q_table[4][3] ), .QN(n179) );
  DF3 \u_cordic/mycordic/present_Q_table_reg[4][4]  ( .D(n1542), .C(inClock), 
        .Q(\u_cordic/mycordic/present_Q_table[4][4] ) );
  DF3 \u_cordic/mycordic/present_Q_table_reg[4][5]  ( .D(n1543), .C(inClock), 
        .Q(\u_cordic/mycordic/present_Q_table[4][5] ), .QN(n227) );
  DF3 \u_cordic/mycordic/present_Q_table_reg[4][6]  ( .D(n1544), .C(inClock), 
        .Q(\u_cordic/mycordic/present_Q_table[4][6] ) );
  DF3 \u_cordic/mycordic/present_Q_table_reg[4][7]  ( .D(n1545), .C(inClock), 
        .Q(\u_cordic/mycordic/present_Q_table[4][7] ), .QN(n48) );
  DF3 \u_cordic/mycordic/present_I_table_reg[4][0]  ( .D(n1562), .C(inClock), 
        .Q(\u_cordic/mycordic/present_I_table[4][0] ) );
  DF3 \u_cordic/mycordic/present_I_table_reg[4][1]  ( .D(n1563), .C(inClock), 
        .Q(\u_cordic/mycordic/present_I_table[4][1] ), .QN(n226) );
  DF3 \u_cordic/mycordic/present_I_table_reg[4][2]  ( .D(n1564), .C(inClock), 
        .Q(\u_cordic/mycordic/present_I_table[4][2] ), .QN(n222) );
  DF3 \u_cordic/mycordic/present_I_table_reg[4][3]  ( .D(n1565), .C(inClock), 
        .Q(\u_cordic/mycordic/present_I_table[4][3] ), .QN(n163) );
  DF3 \u_cordic/mycordic/present_I_table_reg[4][4]  ( .D(n1566), .C(inClock), 
        .Q(\u_cordic/mycordic/present_I_table[4][4] ), .QN(n202) );
  DF3 \u_cordic/mycordic/present_I_table_reg[4][5]  ( .D(n1567), .C(inClock), 
        .Q(\u_cordic/mycordic/present_I_table[4][5] ), .QN(n201) );
  DF3 \u_cordic/mycordic/present_I_table_reg[4][6]  ( .D(n1568), .C(inClock), 
        .Q(\u_cordic/mycordic/present_I_table[4][6] ), .QN(n200) );
  DF3 \u_cordic/mycordic/present_I_table_reg[4][7]  ( .D(n1569), .C(inClock), 
        .Q(\u_cordic/mycordic/present_I_table[4][7] ), .QN(n47) );
  DF3 \u_cordic/mycordic/present_Q_table_reg[4][0]  ( .D(n1570), .C(inClock), 
        .Q(\u_cordic/mycordic/present_Q_table[4][0] ), .QN(n234) );
  DF3 \u_cordic/mycordic/present_Q_table_reg[4][1]  ( .D(n1571), .C(inClock), 
        .Q(\u_cordic/mycordic/present_Q_table[4][1] ) );
  DF3 \u_cordic/mycordic/present_Q_table_reg[4][2]  ( .D(n1572), .C(inClock), 
        .Q(\u_cordic/mycordic/present_Q_table[4][2] ) );
  DF3 \u_cordic/mycordic/present_Q_table_reg[3][7]  ( .D(n1484), .C(inClock), 
        .Q(\u_cordic/mycordic/present_Q_table[3][7] ), .QN(n245) );
  DF3 \u_cordic/mycordic/present_Q_table_reg[3][6]  ( .D(n1483), .C(inClock), 
        .Q(\u_cordic/mycordic/present_Q_table[3][6] ), .QN(n249) );
  DF3 \u_cordic/mycordic/present_Q_table_reg[3][5]  ( .D(n1482), .C(inClock), 
        .Q(\u_cordic/mycordic/present_Q_table[3][5] ), .QN(n203) );
  DF3 \u_cordic/mycordic/present_Q_table_reg[3][4]  ( .D(n1481), .C(inClock), 
        .Q(\u_cordic/mycordic/present_Q_table[3][4] ), .QN(n204) );
  DF3 \u_cordic/mycordic/present_Q_table_reg[3][3]  ( .D(n1480), .C(inClock), 
        .Q(\u_cordic/mycordic/present_Q_table[3][3] ), .QN(n205) );
  DF3 \u_cordic/mycordic/present_Q_table_reg[3][2]  ( .D(n1479), .C(inClock), 
        .Q(\u_cordic/mycordic/present_Q_table[3][2] ), .QN(n174) );
  DF3 \u_cordic/mycordic/present_Q_table_reg[3][1]  ( .D(n1478), .C(inClock), 
        .Q(\u_cordic/mycordic/present_Q_table[3][1] ) );
  DF3 \u_cordic/mycordic/present_Q_table_reg[3][0]  ( .D(n1477), .C(inClock), 
        .Q(\u_cordic/mycordic/present_Q_table[3][0] ), .QN(n231) );
  DF3 \u_cordic/mycordic/present_I_table_reg[3][7]  ( .D(n1476), .C(inClock), 
        .Q(\u_cordic/mycordic/present_I_table[3][7] ), .QN(n246) );
  DF3 \u_cordic/mycordic/present_I_table_reg[3][6]  ( .D(n1475), .C(inClock), 
        .Q(\u_cordic/mycordic/present_I_table[3][6] ), .QN(n250) );
  DF3 \u_cordic/mycordic/present_I_table_reg[3][5]  ( .D(n1474), .C(inClock), 
        .Q(\u_cordic/mycordic/present_I_table[3][5] ), .QN(n206) );
  DF3 \u_cordic/mycordic/present_I_table_reg[3][4]  ( .D(n1473), .C(inClock), 
        .Q(\u_cordic/mycordic/present_I_table[3][4] ), .QN(n207) );
  DF3 \u_cordic/mycordic/present_I_table_reg[3][3]  ( .D(n1472), .C(inClock), 
        .Q(\u_cordic/mycordic/present_I_table[3][3] ), .QN(n208) );
  DF3 \u_cordic/mycordic/present_I_table_reg[3][2]  ( .D(n1471), .C(inClock), 
        .Q(\u_cordic/mycordic/present_I_table[3][2] ), .QN(n176) );
  DF3 \u_cordic/mycordic/present_I_table_reg[3][1]  ( .D(n1470), .C(inClock), 
        .Q(\u_cordic/mycordic/present_I_table[3][1] ) );
  DF3 \u_cordic/mycordic/present_I_table_reg[3][0]  ( .D(n1469), .C(inClock), 
        .Q(\u_cordic/mycordic/present_I_table[3][0] ), .QN(n230) );
  DF3 \u_cordic/mycordic/present_I_table_reg[2][7]  ( .D(n1490), .C(inClock), 
        .Q(\u_cordic/mycordic/present_I_table[2][7] ), .QN(n288) );
  DF3 \u_cordic/mycordic/present_I_table_reg[2][6]  ( .D(n1489), .C(inClock), 
        .Q(\u_cordic/mycordic/present_I_table[2][6] ), .QN(n253) );
  DF3 \u_cordic/mycordic/present_I_table_reg[2][5]  ( .D(n1488), .C(inClock), 
        .Q(\u_cordic/mycordic/present_I_table[2][5] ), .QN(n254) );
  DF3 \u_cordic/mycordic/present_I_table_reg[2][4]  ( .D(n1487), .C(inClock), 
        .Q(\u_cordic/mycordic/present_I_table[2][4] ), .QN(n212) );
  DF3 \u_cordic/mycordic/present_I_table_reg[2][3]  ( .D(n1486), .C(inClock), 
        .Q(\u_cordic/mycordic/present_I_table[2][3] ), .QN(n213) );
  DF3 \u_cordic/mycordic/present_I_table_reg[2][2]  ( .D(n2), .C(inClock), .Q(
        \u_cordic/mycordic/present_I_table[2][2] ), .QN(n214) );
  DF3 \u_cordic/mycordic/present_I_table_reg[2][1]  ( .D(n2), .C(inClock), .Q(
        \u_cordic/mycordic/present_I_table[2][1] ), .QN(n175) );
  DF3 \u_cordic/mycordic/present_I_table_reg[2][0]  ( .D(n2), .C(inClock), .Q(
        \u_cordic/mycordic/present_I_table[2][0] ), .QN(n232) );
  DF3 \u_cordic/mycordic/present_Q_table_reg[2][7]  ( .D(n1495), .C(inClock), 
        .Q(\u_cordic/mycordic/present_Q_table[2][7] ), .QN(n287) );
  DF3 \u_cordic/mycordic/present_Q_table_reg[2][6]  ( .D(n1494), .C(inClock), 
        .Q(\u_cordic/mycordic/present_Q_table[2][6] ), .QN(n251) );
  DF3 \u_cordic/mycordic/present_Q_table_reg[2][5]  ( .D(n1493), .C(inClock), 
        .Q(\u_cordic/mycordic/present_Q_table[2][5] ), .QN(n252) );
  DF3 \u_cordic/mycordic/present_Q_table_reg[2][4]  ( .D(n1492), .C(inClock), 
        .Q(\u_cordic/mycordic/present_Q_table[2][4] ), .QN(n209) );
  DF3 \u_cordic/mycordic/present_Q_table_reg[2][3]  ( .D(n1491), .C(inClock), 
        .Q(\u_cordic/mycordic/present_Q_table[2][3] ), .QN(n210) );
  DF3 \u_cordic/mycordic/present_Q_table_reg[2][2]  ( .D(n2), .C(inClock), .Q(
        \u_cordic/mycordic/present_Q_table[2][2] ), .QN(n211) );
  DF3 \u_cordic/mycordic/present_Q_table_reg[2][1]  ( .D(n2), .C(inClock), .Q(
        \u_cordic/mycordic/present_Q_table[2][1] ), .QN(n173) );
  DF3 \u_cordic/mycordic/present_Q_table_reg[2][0]  ( .D(n2), .C(inClock), .Q(
        \u_cordic/mycordic/present_Q_table[2][0] ), .QN(n233) );
  DF3 \u_cordic/mycordic/present_Q_table_reg[1][7]  ( .D(n1436), .C(inClock), 
        .Q(\u_cordic/mycordic/present_Q_table[1][7] ), .QN(n304) );
  DF3 \u_cordic/mycordic/present_Q_table_reg[1][6]  ( .D(n1435), .C(inClock), 
        .Q(\u_cordic/mycordic/present_Q_table[1][6] ), .QN(n292) );
  DF3 \u_cordic/mycordic/present_Q_table_reg[1][5]  ( .D(n1434), .C(inClock), 
        .Q(\u_cordic/mycordic/present_Q_table[1][5] ), .QN(n258) );
  DF3 \u_cordic/mycordic/present_Q_table_reg[1][4]  ( .D(n1433), .C(inClock), 
        .Q(\u_cordic/mycordic/present_Q_table[1][4] ), .QN(n259) );
  DF3 \u_cordic/mycordic/present_Q_table_reg[1][3]  ( .D(n1432), .C(inClock), 
        .Q(\u_cordic/mycordic/present_Q_table[1][3] ), .QN(n216) );
  DF3 \u_cordic/mycordic/present_Q_table_reg[0][3]  ( .D(\u_cordic/Q [0]), .C(
        inClock), .Q(\u_cordic/mycordic/present_Q_table[0][3] ), .QN(n260) );
  DF3 \u_cordic/mycordic/present_Q_table_reg[0][4]  ( .D(\u_cordic/Q [1]), .C(
        inClock), .Q(\u_cordic/mycordic/present_Q_table[0][4] ), .QN(n55) );
  DF3 \u_cordic/mycordic/present_Q_table_reg[0][5]  ( .D(\u_cordic/Q [2]), .C(
        inClock), .Q(\u_cordic/mycordic/present_Q_table[0][5] ), .QN(n54) );
  DF3 \u_cordic/mycordic/present_Q_table_reg[0][6]  ( .D(\u_cordic/Q [3]), .C(
        inClock), .Q(\u_cordic/mycordic/present_Q_table[0][6] ), .QN(n53) );
  DF3 \u_cordic/mycordic/present_Q_table_reg[0][7]  ( .D(\u_cordic/Q [3]), .C(
        inClock), .Q(\u_cordic/mycordic/present_Q_table[0][7] ) );
  DF3 \u_cordic/mycordic/present_I_table_reg[1][7]  ( .D(
        \u_cordic/mycordic/N44 ), .C(inClock), .Q(
        \u_cordic/mycordic/present_I_table[1][7] ), .QN(n307) );
  DF3 \u_cordic/mycordic/present_I_table_reg[1][6]  ( .D(n1431), .C(inClock), 
        .Q(\u_cordic/mycordic/present_I_table[1][6] ), .QN(n291) );
  DF3 \u_cordic/mycordic/present_I_table_reg[1][5]  ( .D(n1430), .C(inClock), 
        .Q(\u_cordic/mycordic/present_I_table[1][5] ), .QN(n256) );
  DF3 \u_cordic/mycordic/present_I_table_reg[1][4]  ( .D(n1429), .C(inClock), 
        .Q(\u_cordic/mycordic/present_I_table[1][4] ), .QN(n257) );
  DF3 \u_cordic/mycordic/present_I_table_reg[1][3]  ( .D(n1428), .C(inClock), 
        .Q(\u_cordic/mycordic/present_I_table[1][3] ), .QN(n215) );
  DF3 \u_cordic/mycordic/present_I_table_reg[0][3]  ( .D(\u_cordic/I [0]), .C(
        inClock), .Q(\u_cordic/mycordic/present_I_table[0][3] ), .QN(n261) );
  DF3 \u_cordic/mycordic/present_I_table_reg[0][4]  ( .D(\u_cordic/I [1]), .C(
        inClock), .Q(\u_cordic/mycordic/present_I_table[0][4] ), .QN(n58) );
  DF3 \u_cordic/mycordic/present_I_table_reg[0][5]  ( .D(\u_cordic/I [2]), .C(
        inClock), .Q(\u_cordic/mycordic/present_I_table[0][5] ), .QN(n56) );
  DF3 \u_cordic/mycordic/present_I_table_reg[0][6]  ( .D(\u_cordic/I [3]), .C(
        inClock), .Q(\u_cordic/mycordic/present_I_table[0][6] ), .QN(n57) );
  DF3 \u_cordic/mycordic/present_I_table_reg[0][7]  ( .D(\u_cordic/I [3]), .C(
        inClock), .Q(\u_cordic/mycordic/present_I_table[0][7] ), .QN(n303) );
  DF3 \u_cordic/my_rotation/present_direction_reg  ( .D(n1855), .C(inClock), 
        .Q(\u_cordic/dir ) );
  DF3 \u_cordic/my_rotation/present_angle_reg[0][0]  ( .D(n1854), .C(inClock), 
        .Q(\u_cordic/my_rotation/present_angle[0][0] ) );
  DF3 \u_cordic/my_rotation/present_angle_reg[0][1]  ( .D(n1853), .C(inClock), 
        .Q(\u_cordic/my_rotation/present_angle[0][1] ) );
  DF3 \u_cordic/my_rotation/present_angle_reg[0][2]  ( .D(n1852), .C(inClock), 
        .Q(\u_cordic/my_rotation/present_angle[0][2] ) );
  DF3 \u_cordic/my_rotation/present_angle_reg[0][3]  ( .D(n1851), .C(inClock), 
        .Q(\u_cordic/my_rotation/present_angle[0][3] ) );
  DF3 \u_cordic/my_rotation/present_angle_reg[0][4]  ( .D(n1867), .C(inClock), 
        .Q(\u_cordic/my_rotation/present_angle[0][4] ) );
  DF3 \u_cordic/my_rotation/present_angle_reg[0][5]  ( .D(n1866), .C(inClock), 
        .Q(\u_cordic/my_rotation/present_angle[0][5] ) );
  DF3 \u_cordic/my_rotation/present_angle_reg[0][6]  ( .D(n1865), .C(inClock), 
        .Q(\u_cordic/my_rotation/present_angle[0][6] ) );
  DF3 \u_cordic/my_rotation/present_angle_reg[0][7]  ( .D(n1864), .C(inClock), 
        .Q(\u_cordic/my_rotation/present_angle[0][7] ) );
  DF3 \u_cordic/my_rotation/present_angle_reg[0][8]  ( .D(n1863), .C(inClock), 
        .Q(\u_cordic/my_rotation/present_angle[0][8] ) );
  DF3 \u_cordic/my_rotation/present_angle_reg[0][9]  ( .D(n1862), .C(inClock), 
        .Q(\u_cordic/my_rotation/present_angle[0][9] ) );
  DF3 \u_cordic/my_rotation/present_angle_reg[0][10]  ( .D(n1861), .C(inClock), 
        .Q(\u_cordic/my_rotation/present_angle[0][10] ) );
  DF3 \u_cordic/my_rotation/present_angle_reg[0][11]  ( .D(n1860), .C(inClock), 
        .Q(\u_cordic/my_rotation/present_angle[0][11] ) );
  DF3 \u_cordic/my_rotation/present_angle_reg[0][12]  ( .D(n1859), .C(inClock), 
        .Q(\u_cordic/my_rotation/present_angle[0][12] ) );
  DF3 \u_cordic/my_rotation/present_angle_reg[0][13]  ( .D(n1858), .C(inClock), 
        .Q(\u_cordic/my_rotation/present_angle[0][13] ) );
  DF3 \u_cordic/my_rotation/present_angle_reg[0][14]  ( .D(n1857), .C(inClock), 
        .Q(\u_cordic/my_rotation/present_angle[0][14] ) );
  DF3 \u_cordic/my_rotation/present_angle_reg[0][15]  ( .D(n1856), .C(inClock), 
        .Q(\u_cordic/my_rotation/present_angle[0][15] ) );
  DF3 \u_cdr/div1/o_nb_P_reg[2]  ( .D(\u_cdr/div1/n37 ), .C(n1401), .Q(
        \u_cdr/w_nb_P [2]), .QN(\u_cdr/div1/n9 ) );
  DF3 \u_cdr/div1/o_nb_P_reg[1]  ( .D(\u_cdr/div1/n38 ), .C(n1401), .Q(
        \u_cdr/w_nb_P [1]), .QN(\u_cdr/div1/n10 ) );
  DF3 \u_cdr/div1/o_nb_P_reg[3]  ( .D(\u_cdr/div1/n36 ), .C(n1401), .Q(
        \u_cdr/w_nb_P [3]), .QN(\u_cdr/div1/n8 ) );
  DF3 \u_cdr/div1/o_nb_P_reg[4]  ( .D(\u_cdr/div1/n35 ), .C(n1401), .Q(
        \u_cdr/w_nb_P [4]), .QN(n60) );
  DF3 \u_cdr/div1/o_nb_P_reg[5]  ( .D(\u_cdr/div1/n39 ), .C(n1401), .Q(
        \u_cdr/w_nb_P [5]), .QN(\u_cdr/div1/n7 ) );
  DF3 \u_cdr/div1/o_nb_P_reg[0]  ( .D(\u_cdr/div1/n40 ), .C(n1401), .Q(
        \u_cdr/div1/N35 ), .QN(n59) );
  DF3 \u_cdr/phd1/o_T_reg  ( .D(\u_cdr/phd1/n22 ), .C(n1401), .Q(\u_cdr/w_sT )
         );
  DF3 \u_cdr/phd1/o_E_reg  ( .D(\u_cdr/phd1/n23 ), .C(n1401), .Q(\u_cdr/w_sE ), 
        .QN(n221) );
  DF3 \u_cdr/dec1/o_data_reg  ( .D(n1849), .C(inClock), .Q(
        \sig_MUX_inMUX13[0] ), .QN(\u_cdr/dec1/n20 ) );
  DF3 \u_cdr/dec1/o_flag_reg  ( .D(\u_cdr/dec1/N73 ), .C(inClock), .Q(
        \sig_MUX_inMUX12[0] ), .QN(n52) );
  DF3 \u_cdr/dec1/cnt_r_reg[1]  ( .D(n1422), .C(inClock), .Q(
        \u_cdr/dec1/cnt_r [1]) );
  DF3 \u_cdr/dec1/cnt_r_reg[2]  ( .D(n1423), .C(inClock), .Q(
        \u_cdr/dec1/cnt_r [2]) );
  DF3 \u_cdr/dec1/cnt_r_reg[3]  ( .D(n1424), .C(inClock), .Q(
        \u_cdr/dec1/cnt_r [3]) );
  DF3 \u_cdr/dec1/cnt_r_reg[4]  ( .D(n1425), .C(inClock), .Q(
        \u_cdr/dec1/cnt_r [4]) );
  DF3 \u_cdr/dec1/cnt_r_reg[5]  ( .D(n1421), .C(inClock), .Q(
        \u_cdr/dec1/cnt_r [5]), .QN(n301) );
  DF3 \u_cdr/dec1/cnt_r_reg[0]  ( .D(n1420), .C(inClock), .Q(
        \u_cdr/dec1/cnt_r [0]), .QN(n248) );
  DF3 \u_inFIFO/os1/dff1/s_qout_reg  ( .D(n1848), .C(inClock), .Q(
        \u_inFIFO/os1/sigQout1 ), .QN(n318) );
  DF3 \u_decoder/iq_demod/cossin_dig/o_cos_reg[0]  ( .D(n2680), .C(inClock), 
        .Q(\u_decoder/iq_demod/cos_out [0]), .QN(n40) );
  DF3 \u_decoder/iq_demod/cossin_dig/o_cos_reg[1]  ( .D(
        \u_decoder/iq_demod/cossin_dig/n49 ), .C(inClock), .Q(
        \u_decoder/iq_demod/cos_out [1]), .QN(n41) );
  DF3 \u_decoder/iq_demod/cossin_dig/o_cos_reg[2]  ( .D(
        \u_decoder/iq_demod/cossin_dig/n50 ), .C(inClock), .Q(
        \u_decoder/iq_demod/cos_out [2]), .QN(n43) );
  DF3 \u_decoder/iq_demod/cossin_dig/o_cos_reg[3]  ( .D(n2681), .C(inClock), 
        .Q(\u_decoder/iq_demod/cos_out [3]), .QN(n22) );
  DF3 \u_decoder/iq_demod/cossin_dig/o_sin_reg[0]  ( .D(
        \u_decoder/iq_demod/cossin_dig/n51 ), .C(inClock), .Q(
        \u_decoder/iq_demod/sin_out [0]), .QN(n42) );
  DF3 \u_decoder/iq_demod/cossin_dig/o_sin_reg[1]  ( .D(n2682), .C(inClock), 
        .Q(\u_decoder/iq_demod/sin_out [1]), .QN(n44) );
  DF3 \u_decoder/iq_demod/cossin_dig/o_sin_reg[2]  ( .D(n2683), .C(inClock), 
        .Q(\u_decoder/iq_demod/sin_out [2]), .QN(n45) );
  DF3 \u_decoder/iq_demod/cossin_dig/o_sin_reg[3]  ( .D(n2684), .C(inClock), 
        .Q(\u_decoder/iq_demod/sin_out [3]), .QN(n23) );
  DF3 \u_decoder/iq_demod/cossin_dig/val_counter_reg[2]  ( .D(n1846), .C(
        inClock), .Q(\u_decoder/iq_demod/cossin_dig/val_counter [2]) );
  DF3 \u_decoder/iq_demod/cossin_dig/val_counter_reg[1]  ( .D(
        \u_decoder/iq_demod/cossin_dig/n52 ), .C(inClock), .Q(
        \u_decoder/iq_demod/cossin_dig/val_counter [1]), .QN(
        \u_decoder/iq_demod/cossin_dig/n19 ) );
  DF3 \u_decoder/iq_demod/cossin_dig/val_counter_reg[0]  ( .D(
        \u_decoder/iq_demod/cossin_dig/n53 ), .C(inClock), .Q(
        \u_decoder/iq_demod/cossin_dig/N55 ), .QN(
        \u_decoder/iq_demod/cossin_dig/n21 ) );
  DF3 \u_decoder/iq_demod/cossin_dig/state_reg[1]  ( .D(
        \u_decoder/iq_demod/cossin_dig/N42 ), .C(inClock), .QN(
        \u_decoder/iq_demod/cossin_dig/n23 ) );
  DF3 \u_decoder/iq_demod/cossin_dig/counter_reg[2]  ( .D(
        \u_decoder/iq_demod/cossin_dig/N22 ), .C(inClock), .Q(
        \u_decoder/iq_demod/cossin_dig/counter [2]), .QN(
        \u_decoder/iq_demod/cossin_dig/n10 ) );
  DF3 \u_decoder/iq_demod/cossin_dig/counter_reg[1]  ( .D(
        \u_decoder/iq_demod/cossin_dig/N21 ), .C(inClock), .Q(
        \u_decoder/iq_demod/cossin_dig/counter [1]) );
  DF3 \u_decoder/iq_demod/cossin_dig/counter_reg[0]  ( .D(
        \u_decoder/iq_demod/cossin_dig/N20 ), .C(inClock), .Q(
        \u_decoder/iq_demod/cossin_dig/counter [0]) );
  DF3 \u_decoder/iq_demod/cossin_dig/state_reg[0]  ( .D(
        \u_decoder/iq_demod/cossin_dig/N41 ), .C(inClock), .Q(
        \u_decoder/iq_demod/cossin_dig/state[0] ) );
  DF3 \u_cdr/div1/cnt_div/o_en_freq_synch_reg  ( .D(\u_cdr/div1/cnt_div/N88 ), 
        .C(inClock), .Q(\u_cdr/div1/w_en_freq_synch ) );
  DF3 \u_cdr/div1/cnt_div/cnt_reg[1]  ( .D(n1416), .C(inClock), .Q(
        \u_cdr/div1/cnt_div/cnt [1]) );
  DF3 \u_cdr/div1/cnt_div/cnt_reg[2]  ( .D(n1417), .C(inClock), .Q(
        \u_cdr/div1/cnt_div/cnt [2]) );
  DF3 \u_cdr/div1/cnt_div/cnt_reg[3]  ( .D(n1418), .C(inClock), .Q(
        \u_cdr/div1/cnt_div/cnt [3]) );
  DF3 \u_cdr/div1/cnt_div/cnt_reg[4]  ( .D(n1419), .C(inClock), .Q(
        \u_cdr/div1/cnt_div/cnt [4]) );
  DF3 \u_cdr/div1/cnt_div/cnt_reg[5]  ( .D(n1415), .C(inClock), .Q(
        \u_cdr/div1/cnt_div/cnt [5]) );
  DF3 \u_cdr/div1/cnt_div/cnt_reg[0]  ( .D(n1414), .C(inClock), .Q(
        \u_cdr/div1/cnt_div/cnt [0]), .QN(n262) );
  DF3 \u_cdr/phd1/f1/o_Q_reg  ( .D(n1844), .C(inClock), .Q(\u_cdr/phd1/w_s1 )
         );
  DF3 \u_cdr/dec1/cnt_dec/o_en_dec_reg  ( .D(\u_cdr/dec1/cnt_dec/N33 ), .C(
        inClock), .Q(\u_cdr/dec1/w_en_dec ), .QN(n306) );
  DF3 \u_cdr/dec1/cnt_dec/cnt_dec_reg[5]  ( .D(n1413), .C(inClock), .Q(
        \u_cdr/dec1/cnt_dec/cnt_dec [5]), .QN(n315) );
  DF3 \u_cdr/dec1/cnt_dec/cnt_dec_reg[4]  ( .D(n1412), .C(inClock), .Q(
        \u_cdr/dec1/cnt_dec/cnt_dec [4]) );
  DF3 \u_cdr/dec1/cnt_dec/cnt_dec_reg[3]  ( .D(n1411), .C(inClock), .Q(
        \u_cdr/dec1/cnt_dec/cnt_dec [3]) );
  DF3 \u_cdr/dec1/cnt_dec/cnt_dec_reg[2]  ( .D(n1410), .C(inClock), .Q(
        \u_cdr/dec1/cnt_dec/cnt_dec [2]) );
  DF3 \u_cdr/dec1/cnt_dec/cnt_dec_reg[1]  ( .D(n1409), .C(inClock), .Q(
        \u_cdr/dec1/cnt_dec/cnt_dec [1]), .QN(n302) );
  DF3 \u_cdr/dec1/cnt_dec/cnt_dec_reg[0]  ( .D(n1408), .C(inClock), .Q(
        \u_cdr/dec1/cnt_dec/cnt_dec [0]), .QN(n263) );
  DF3 \u_outFIFO/os2/dff2/s_qout_reg  ( .D(n1843), .C(inClock), .Q(
        \u_outFIFO/os2/sigQout2 ) );
  DF3 \u_outFIFO/os2/dff1/s_qout_reg  ( .D(n1842), .C(inClock), .Q(
        \u_outFIFO/os2/sigQout1 ), .QN(n285) );
  DF3 \u_outFIFO/os1/dff2/s_qout_reg  ( .D(n1841), .C(inClock), .Q(
        \u_outFIFO/os1/sigQout2 ) );
  DF3 \u_outFIFO/os1/dff1/s_qout_reg  ( .D(n1840), .C(inClock), .Q(
        \u_outFIFO/os1/sigQout1 ), .QN(n284) );
  DF3 \u_inFIFO/os2/dff2/s_qout_reg  ( .D(n1839), .C(inClock), .Q(
        \u_inFIFO/os2/sigQout2 ) );
  DF3 \u_inFIFO/os2/dff1/s_qout_reg  ( .D(n1838), .C(inClock), .Q(
        \u_inFIFO/os2/sigQout1 ), .QN(n317) );
  DF3 \u_inFIFO/os1/dff2/s_qout_reg  ( .D(n1837), .C(inClock), .Q(
        \u_inFIFO/os1/sigQout2 ) );
  DF3 \u_cdr/phd1/cnt_phd/o_en_reg  ( .D(n1834), .C(inClock), .QN(n62) );
  DF3 \u_cdr/phd1/cnt_phd/o_en_f_reg  ( .D(n1835), .C(inClock), .Q(
        \u_cdr/phd1/w_en_f ), .QN(n300) );
  DF3 \u_cdr/phd1/cnt_phd/o_en_m_reg  ( .D(n1836), .C(inClock), .Q(
        \u_cdr/phd1/w_en_m ), .QN(n319) );
  DF3 \u_cdr/phd1/cnt_phd/o_en_d_reg  ( .D(\u_cdr/phd1/cnt_phd/N84 ), .C(
        inClock), .Q(\u_cdr/phd1/w_en_d ) );
  DF3 \u_cdr/phd1/cnt_phd/cnt_reg[1]  ( .D(n1404), .C(inClock), .Q(
        \u_cdr/phd1/cnt_phd/cnt [1]), .QN(n293) );
  DF3 \u_cdr/phd1/cnt_phd/cnt_reg[2]  ( .D(n1405), .C(inClock), .Q(
        \u_cdr/phd1/cnt_phd/cnt [2]) );
  DF3 \u_cdr/phd1/cnt_phd/cnt_reg[3]  ( .D(n1406), .C(inClock), .Q(
        \u_cdr/phd1/cnt_phd/cnt [3]) );
  DF3 \u_cdr/phd1/cnt_phd/cnt_reg[4]  ( .D(n1407), .C(inClock), .Q(
        \u_cdr/phd1/cnt_phd/cnt [4]) );
  DF3 \u_cdr/phd1/cnt_phd/cnt_reg[5]  ( .D(n1403), .C(inClock), .Q(
        \u_cdr/phd1/cnt_phd/cnt [5]), .QN(n255) );
  DF3 \u_cdr/phd1/cnt_phd/cnt_reg[0]  ( .D(n1402), .C(inClock), .Q(
        \u_cdr/phd1/cnt_phd/cnt [0]), .QN(n3055) );
  DF3 \u_cdr/dec1/ffd_retard/o_Q_reg  ( .D(n1833), .C(inClock), .Q(
        \u_cdr/dec1/w_s_r ), .QN(n316) );
  DF3 \u_cdr/phd1/f4/o_Q_reg  ( .D(n1832), .C(inClock), .Q(\u_cdr/phd1/w_s4 )
         );
  DF3 \u_cdr/phd1/f3/o_Q_reg  ( .D(n1831), .C(inClock), .Q(\u_cdr/phd1/w_s3 )
         );
  DF3 \u_cdr/phd1/f2/o_Q_reg  ( .D(n1830), .C(inClock), .Q(\u_cdr/phd1/w_s2 )
         );
  DFE1 \u_cdr/dir_f_reg  ( .D(n1914), .E(\u_cdr/n45 ), .C(inClock), .QN(
        \u_cdr/n3 ) );
  DFE1 \u_cdr/dir_d_reg  ( .D(n1914), .E(\u_cdr/n31 ), .C(inClock), .QN(
        \u_cdr/n19 ) );
  DFE1 \u_outFIFO/FIFO_reg[2][0]  ( .D(n982), .E(\u_outFIFO/n330 ), .C(inClock), .Q(\u_outFIFO/FIFO[2][0] ) );
  DFE1 \u_outFIFO/FIFO_reg[2][1]  ( .D(n982), .E(\u_outFIFO/n332 ), .C(inClock), .Q(\u_outFIFO/FIFO[2][1] ) );
  DFE1 \u_outFIFO/FIFO_reg[2][2]  ( .D(n982), .E(\u_outFIFO/n333 ), .C(inClock), .Q(\u_outFIFO/FIFO[2][2] ) );
  DFE1 \u_outFIFO/FIFO_reg[2][3]  ( .D(n982), .E(\u_outFIFO/n334 ), .C(inClock), .Q(\u_outFIFO/FIFO[2][3] ) );
  DFE1 \u_outFIFO/FIFO_reg[6][0]  ( .D(n984), .E(\u_outFIFO/n350 ), .C(inClock), .Q(\u_outFIFO/FIFO[6][0] ) );
  DFE1 \u_outFIFO/FIFO_reg[6][1]  ( .D(n984), .E(\u_outFIFO/n352 ), .C(inClock), .Q(\u_outFIFO/FIFO[6][1] ) );
  DFE1 \u_outFIFO/FIFO_reg[6][2]  ( .D(n984), .E(\u_outFIFO/n353 ), .C(inClock), .Q(\u_outFIFO/FIFO[6][2] ) );
  DFE1 \u_outFIFO/FIFO_reg[6][3]  ( .D(n984), .E(\u_outFIFO/n354 ), .C(inClock), .Q(\u_outFIFO/FIFO[6][3] ) );
  DFE1 \u_outFIFO/FIFO_reg[10][0]  ( .D(n986), .E(\u_outFIFO/n370 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[10][0] ) );
  DFE1 \u_outFIFO/FIFO_reg[10][1]  ( .D(n986), .E(\u_outFIFO/n372 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[10][1] ) );
  DFE1 \u_outFIFO/FIFO_reg[10][2]  ( .D(n986), .E(\u_outFIFO/n373 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[10][2] ) );
  DFE1 \u_outFIFO/FIFO_reg[10][3]  ( .D(n986), .E(\u_outFIFO/n374 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[10][3] ) );
  DFE1 \u_outFIFO/FIFO_reg[14][0]  ( .D(n988), .E(\u_outFIFO/n390 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[14][0] ) );
  DFE1 \u_outFIFO/FIFO_reg[14][1]  ( .D(n988), .E(\u_outFIFO/n392 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[14][1] ) );
  DFE1 \u_outFIFO/FIFO_reg[14][2]  ( .D(n988), .E(\u_outFIFO/n393 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[14][2] ) );
  DFE1 \u_outFIFO/FIFO_reg[14][3]  ( .D(n988), .E(\u_outFIFO/n394 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[14][3] ) );
  DFE1 \u_outFIFO/FIFO_reg[18][0]  ( .D(n990), .E(\u_outFIFO/n416 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[18][0] ) );
  DFE1 \u_outFIFO/FIFO_reg[18][1]  ( .D(n990), .E(\u_outFIFO/n417 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[18][1] ) );
  DFE1 \u_outFIFO/FIFO_reg[18][2]  ( .D(n990), .E(\u_outFIFO/n418 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[18][2] ) );
  DFE1 \u_outFIFO/FIFO_reg[18][3]  ( .D(n990), .E(\u_outFIFO/n419 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[18][3] ) );
  DFE1 \u_outFIFO/FIFO_reg[22][0]  ( .D(n992), .E(\u_outFIFO/n432 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[22][0] ) );
  DFE1 \u_outFIFO/FIFO_reg[22][1]  ( .D(n992), .E(\u_outFIFO/n433 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[22][1] ) );
  DFE1 \u_outFIFO/FIFO_reg[22][2]  ( .D(n992), .E(\u_outFIFO/n434 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[22][2] ) );
  DFE1 \u_outFIFO/FIFO_reg[22][3]  ( .D(n992), .E(\u_outFIFO/n435 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[22][3] ) );
  DFE1 \u_outFIFO/FIFO_reg[26][0]  ( .D(n994), .E(\u_outFIFO/n448 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[26][0] ) );
  DFE1 \u_outFIFO/FIFO_reg[26][1]  ( .D(n994), .E(\u_outFIFO/n449 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[26][1] ) );
  DFE1 \u_outFIFO/FIFO_reg[26][2]  ( .D(n994), .E(\u_outFIFO/n450 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[26][2] ) );
  DFE1 \u_outFIFO/FIFO_reg[26][3]  ( .D(n994), .E(\u_outFIFO/n451 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[26][3] ) );
  DFE1 \u_outFIFO/FIFO_reg[30][0]  ( .D(n996), .E(\u_outFIFO/n464 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[30][0] ) );
  DFE1 \u_outFIFO/FIFO_reg[30][1]  ( .D(n996), .E(\u_outFIFO/n465 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[30][1] ) );
  DFE1 \u_outFIFO/FIFO_reg[30][2]  ( .D(n996), .E(\u_outFIFO/n466 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[30][2] ) );
  DFE1 \u_outFIFO/FIFO_reg[30][3]  ( .D(n996), .E(\u_outFIFO/n467 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[30][3] ) );
  DFE1 \u_outFIFO/FIFO_reg[34][0]  ( .D(n998), .E(\u_outFIFO/n485 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[34][0] ) );
  DFE1 \u_outFIFO/FIFO_reg[34][1]  ( .D(n998), .E(\u_outFIFO/n486 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[34][1] ) );
  DFE1 \u_outFIFO/FIFO_reg[34][2]  ( .D(n998), .E(\u_outFIFO/n487 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[34][2] ) );
  DFE1 \u_outFIFO/FIFO_reg[34][3]  ( .D(n998), .E(\u_outFIFO/n488 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[34][3] ) );
  DFE1 \u_outFIFO/FIFO_reg[38][0]  ( .D(n1000), .E(\u_outFIFO/n501 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[38][0] ) );
  DFE1 \u_outFIFO/FIFO_reg[38][1]  ( .D(n1000), .E(\u_outFIFO/n502 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[38][1] ) );
  DFE1 \u_outFIFO/FIFO_reg[38][2]  ( .D(n1000), .E(\u_outFIFO/n503 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[38][2] ) );
  DFE1 \u_outFIFO/FIFO_reg[38][3]  ( .D(n1000), .E(\u_outFIFO/n504 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[38][3] ) );
  DFE1 \u_outFIFO/FIFO_reg[42][0]  ( .D(n1002), .E(\u_outFIFO/n517 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[42][0] ) );
  DFE1 \u_outFIFO/FIFO_reg[42][1]  ( .D(n1002), .E(\u_outFIFO/n518 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[42][1] ) );
  DFE1 \u_outFIFO/FIFO_reg[42][2]  ( .D(n1002), .E(\u_outFIFO/n519 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[42][2] ) );
  DFE1 \u_outFIFO/FIFO_reg[42][3]  ( .D(n1002), .E(\u_outFIFO/n520 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[42][3] ) );
  DFE1 \u_outFIFO/FIFO_reg[46][0]  ( .D(n1004), .E(\u_outFIFO/n533 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[46][0] ) );
  DFE1 \u_outFIFO/FIFO_reg[46][1]  ( .D(n1004), .E(\u_outFIFO/n534 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[46][1] ) );
  DFE1 \u_outFIFO/FIFO_reg[46][2]  ( .D(n1004), .E(\u_outFIFO/n535 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[46][2] ) );
  DFE1 \u_outFIFO/FIFO_reg[46][3]  ( .D(n1004), .E(\u_outFIFO/n536 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[46][3] ) );
  DFE1 \u_outFIFO/FIFO_reg[50][0]  ( .D(n1006), .E(\u_outFIFO/n554 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[50][0] ) );
  DFE1 \u_outFIFO/FIFO_reg[50][1]  ( .D(n1006), .E(\u_outFIFO/n555 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[50][1] ) );
  DFE1 \u_outFIFO/FIFO_reg[50][2]  ( .D(n1006), .E(\u_outFIFO/n556 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[50][2] ) );
  DFE1 \u_outFIFO/FIFO_reg[50][3]  ( .D(n1006), .E(\u_outFIFO/n557 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[50][3] ) );
  DFE1 \u_outFIFO/FIFO_reg[54][0]  ( .D(n1008), .E(\u_outFIFO/n570 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[54][0] ) );
  DFE1 \u_outFIFO/FIFO_reg[54][1]  ( .D(n1008), .E(\u_outFIFO/n571 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[54][1] ) );
  DFE1 \u_outFIFO/FIFO_reg[54][2]  ( .D(n1008), .E(\u_outFIFO/n572 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[54][2] ) );
  DFE1 \u_outFIFO/FIFO_reg[54][3]  ( .D(n1008), .E(\u_outFIFO/n573 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[54][3] ) );
  DFE1 \u_outFIFO/FIFO_reg[58][0]  ( .D(n1010), .E(\u_outFIFO/n586 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[58][0] ) );
  DFE1 \u_outFIFO/FIFO_reg[58][1]  ( .D(n1010), .E(\u_outFIFO/n587 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[58][1] ) );
  DFE1 \u_outFIFO/FIFO_reg[58][2]  ( .D(n1010), .E(\u_outFIFO/n588 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[58][2] ) );
  DFE1 \u_outFIFO/FIFO_reg[58][3]  ( .D(n1010), .E(\u_outFIFO/n589 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[58][3] ) );
  DFE1 \u_outFIFO/FIFO_reg[62][0]  ( .D(n1012), .E(\u_outFIFO/n602 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[62][0] ) );
  DFE1 \u_outFIFO/FIFO_reg[62][1]  ( .D(n1012), .E(\u_outFIFO/n603 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[62][1] ) );
  DFE1 \u_outFIFO/FIFO_reg[62][2]  ( .D(n1012), .E(\u_outFIFO/n604 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[62][2] ) );
  DFE1 \u_outFIFO/FIFO_reg[62][3]  ( .D(n1012), .E(\u_outFIFO/n605 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[62][3] ) );
  DFE1 \u_outFIFO/FIFO_reg[66][0]  ( .D(n1014), .E(\u_outFIFO/n623 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[66][0] ) );
  DFE1 \u_outFIFO/FIFO_reg[66][1]  ( .D(n1014), .E(\u_outFIFO/n624 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[66][1] ) );
  DFE1 \u_outFIFO/FIFO_reg[66][2]  ( .D(n1014), .E(\u_outFIFO/n625 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[66][2] ) );
  DFE1 \u_outFIFO/FIFO_reg[66][3]  ( .D(n1014), .E(\u_outFIFO/n626 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[66][3] ) );
  DFE1 \u_outFIFO/FIFO_reg[70][0]  ( .D(n1016), .E(\u_outFIFO/n639 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[70][0] ) );
  DFE1 \u_outFIFO/FIFO_reg[70][1]  ( .D(n1016), .E(\u_outFIFO/n640 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[70][1] ) );
  DFE1 \u_outFIFO/FIFO_reg[70][2]  ( .D(n1016), .E(\u_outFIFO/n641 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[70][2] ) );
  DFE1 \u_outFIFO/FIFO_reg[70][3]  ( .D(n1016), .E(\u_outFIFO/n642 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[70][3] ) );
  DFE1 \u_outFIFO/FIFO_reg[74][0]  ( .D(n1018), .E(\u_outFIFO/n655 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[74][0] ) );
  DFE1 \u_outFIFO/FIFO_reg[74][1]  ( .D(n1018), .E(\u_outFIFO/n656 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[74][1] ) );
  DFE1 \u_outFIFO/FIFO_reg[74][2]  ( .D(n1018), .E(\u_outFIFO/n657 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[74][2] ) );
  DFE1 \u_outFIFO/FIFO_reg[74][3]  ( .D(n1018), .E(\u_outFIFO/n658 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[74][3] ) );
  DFE1 \u_cdr/dir_m_reg  ( .D(n1914), .E(\u_cdr/n28 ), .C(inClock), .QN(
        \u_cdr/n20 ) );
  DFE1 \u_outFIFO/FIFO_reg[0][0]  ( .D(n981), .E(\u_outFIFO/n316 ), .C(inClock), .Q(\u_outFIFO/FIFO[0][0] ) );
  DFE1 \u_outFIFO/FIFO_reg[0][1]  ( .D(n981), .E(\u_outFIFO/n319 ), .C(inClock), .Q(\u_outFIFO/FIFO[0][1] ) );
  DFE1 \u_outFIFO/FIFO_reg[0][2]  ( .D(n981), .E(\u_outFIFO/n321 ), .C(inClock), .Q(\u_outFIFO/FIFO[0][2] ) );
  DFE1 \u_outFIFO/FIFO_reg[0][3]  ( .D(n981), .E(\u_outFIFO/n323 ), .C(inClock), .Q(\u_outFIFO/FIFO[0][3] ) );
  DFE1 \u_outFIFO/FIFO_reg[1][0]  ( .D(n981), .E(\u_outFIFO/n325 ), .C(inClock), .Q(\u_outFIFO/FIFO[1][0] ) );
  DFE1 \u_outFIFO/FIFO_reg[1][1]  ( .D(n981), .E(\u_outFIFO/n327 ), .C(inClock), .Q(\u_outFIFO/FIFO[1][1] ) );
  DFE1 \u_outFIFO/FIFO_reg[1][2]  ( .D(n981), .E(\u_outFIFO/n328 ), .C(inClock), .Q(\u_outFIFO/FIFO[1][2] ) );
  DFE1 \u_outFIFO/FIFO_reg[1][3]  ( .D(n981), .E(\u_outFIFO/n329 ), .C(inClock), .Q(\u_outFIFO/FIFO[1][3] ) );
  DFE1 \u_outFIFO/FIFO_reg[3][0]  ( .D(n982), .E(\u_outFIFO/n335 ), .C(inClock), .Q(\u_outFIFO/FIFO[3][0] ) );
  DFE1 \u_outFIFO/FIFO_reg[3][1]  ( .D(n982), .E(\u_outFIFO/n337 ), .C(inClock), .Q(\u_outFIFO/FIFO[3][1] ) );
  DFE1 \u_outFIFO/FIFO_reg[3][2]  ( .D(n982), .E(\u_outFIFO/n338 ), .C(inClock), .Q(\u_outFIFO/FIFO[3][2] ) );
  DFE1 \u_outFIFO/FIFO_reg[3][3]  ( .D(n982), .E(\u_outFIFO/n339 ), .C(inClock), .Q(\u_outFIFO/FIFO[3][3] ) );
  DFE1 \u_outFIFO/FIFO_reg[4][0]  ( .D(n983), .E(\u_outFIFO/n340 ), .C(inClock), .Q(\u_outFIFO/FIFO[4][0] ) );
  DFE1 \u_outFIFO/FIFO_reg[4][1]  ( .D(n983), .E(\u_outFIFO/n342 ), .C(inClock), .Q(\u_outFIFO/FIFO[4][1] ) );
  DFE1 \u_outFIFO/FIFO_reg[4][2]  ( .D(n983), .E(\u_outFIFO/n343 ), .C(inClock), .Q(\u_outFIFO/FIFO[4][2] ) );
  DFE1 \u_outFIFO/FIFO_reg[4][3]  ( .D(n983), .E(\u_outFIFO/n344 ), .C(inClock), .Q(\u_outFIFO/FIFO[4][3] ) );
  DFE1 \u_outFIFO/FIFO_reg[5][0]  ( .D(n983), .E(\u_outFIFO/n345 ), .C(inClock), .Q(\u_outFIFO/FIFO[5][0] ) );
  DFE1 \u_outFIFO/FIFO_reg[5][1]  ( .D(n983), .E(\u_outFIFO/n347 ), .C(inClock), .Q(\u_outFIFO/FIFO[5][1] ) );
  DFE1 \u_outFIFO/FIFO_reg[5][2]  ( .D(n983), .E(\u_outFIFO/n348 ), .C(inClock), .Q(\u_outFIFO/FIFO[5][2] ) );
  DFE1 \u_outFIFO/FIFO_reg[5][3]  ( .D(n983), .E(\u_outFIFO/n349 ), .C(inClock), .Q(\u_outFIFO/FIFO[5][3] ) );
  DFE1 \u_outFIFO/FIFO_reg[7][0]  ( .D(n984), .E(\u_outFIFO/n355 ), .C(inClock), .Q(\u_outFIFO/FIFO[7][0] ) );
  DFE1 \u_outFIFO/FIFO_reg[7][1]  ( .D(n984), .E(\u_outFIFO/n357 ), .C(inClock), .Q(\u_outFIFO/FIFO[7][1] ) );
  DFE1 \u_outFIFO/FIFO_reg[7][2]  ( .D(n984), .E(\u_outFIFO/n358 ), .C(inClock), .Q(\u_outFIFO/FIFO[7][2] ) );
  DFE1 \u_outFIFO/FIFO_reg[7][3]  ( .D(n984), .E(\u_outFIFO/n359 ), .C(inClock), .Q(\u_outFIFO/FIFO[7][3] ) );
  DFE1 \u_outFIFO/FIFO_reg[8][0]  ( .D(n985), .E(\u_outFIFO/n360 ), .C(inClock), .Q(\u_outFIFO/FIFO[8][0] ) );
  DFE1 \u_outFIFO/FIFO_reg[8][1]  ( .D(n985), .E(\u_outFIFO/n362 ), .C(inClock), .Q(\u_outFIFO/FIFO[8][1] ) );
  DFE1 \u_outFIFO/FIFO_reg[8][2]  ( .D(n985), .E(\u_outFIFO/n363 ), .C(inClock), .Q(\u_outFIFO/FIFO[8][2] ) );
  DFE1 \u_outFIFO/FIFO_reg[8][3]  ( .D(n985), .E(\u_outFIFO/n364 ), .C(inClock), .Q(\u_outFIFO/FIFO[8][3] ) );
  DFE1 \u_outFIFO/FIFO_reg[9][0]  ( .D(n985), .E(\u_outFIFO/n365 ), .C(inClock), .Q(\u_outFIFO/FIFO[9][0] ) );
  DFE1 \u_outFIFO/FIFO_reg[9][1]  ( .D(n985), .E(\u_outFIFO/n367 ), .C(inClock), .Q(\u_outFIFO/FIFO[9][1] ) );
  DFE1 \u_outFIFO/FIFO_reg[9][2]  ( .D(n985), .E(\u_outFIFO/n368 ), .C(inClock), .Q(\u_outFIFO/FIFO[9][2] ) );
  DFE1 \u_outFIFO/FIFO_reg[9][3]  ( .D(n985), .E(\u_outFIFO/n369 ), .C(inClock), .Q(\u_outFIFO/FIFO[9][3] ) );
  DFE1 \u_outFIFO/FIFO_reg[11][0]  ( .D(n986), .E(\u_outFIFO/n375 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[11][0] ) );
  DFE1 \u_outFIFO/FIFO_reg[11][1]  ( .D(n986), .E(\u_outFIFO/n377 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[11][1] ) );
  DFE1 \u_outFIFO/FIFO_reg[11][2]  ( .D(n986), .E(\u_outFIFO/n378 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[11][2] ) );
  DFE1 \u_outFIFO/FIFO_reg[11][3]  ( .D(n986), .E(\u_outFIFO/n379 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[11][3] ) );
  DFE1 \u_outFIFO/FIFO_reg[12][0]  ( .D(n987), .E(\u_outFIFO/n380 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[12][0] ) );
  DFE1 \u_outFIFO/FIFO_reg[12][1]  ( .D(n987), .E(\u_outFIFO/n382 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[12][1] ) );
  DFE1 \u_outFIFO/FIFO_reg[12][2]  ( .D(n987), .E(\u_outFIFO/n383 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[12][2] ) );
  DFE1 \u_outFIFO/FIFO_reg[12][3]  ( .D(n987), .E(\u_outFIFO/n384 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[12][3] ) );
  DFE1 \u_outFIFO/FIFO_reg[13][0]  ( .D(n987), .E(\u_outFIFO/n385 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[13][0] ) );
  DFE1 \u_outFIFO/FIFO_reg[13][1]  ( .D(n987), .E(\u_outFIFO/n387 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[13][1] ) );
  DFE1 \u_outFIFO/FIFO_reg[13][2]  ( .D(n987), .E(\u_outFIFO/n388 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[13][2] ) );
  DFE1 \u_outFIFO/FIFO_reg[13][3]  ( .D(n987), .E(\u_outFIFO/n389 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[13][3] ) );
  DFE1 \u_outFIFO/FIFO_reg[15][0]  ( .D(n988), .E(\u_outFIFO/n395 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[15][0] ) );
  DFE1 \u_outFIFO/FIFO_reg[15][1]  ( .D(n988), .E(\u_outFIFO/n398 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[15][1] ) );
  DFE1 \u_outFIFO/FIFO_reg[15][2]  ( .D(n988), .E(\u_outFIFO/n400 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[15][2] ) );
  DFE1 \u_outFIFO/FIFO_reg[15][3]  ( .D(n988), .E(\u_outFIFO/n402 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[15][3] ) );
  DFE1 \u_outFIFO/FIFO_reg[16][0]  ( .D(n989), .E(\u_outFIFO/n404 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[16][0] ) );
  DFE1 \u_outFIFO/FIFO_reg[16][1]  ( .D(n989), .E(\u_outFIFO/n406 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[16][1] ) );
  DFE1 \u_outFIFO/FIFO_reg[16][2]  ( .D(n989), .E(\u_outFIFO/n408 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[16][2] ) );
  DFE1 \u_outFIFO/FIFO_reg[16][3]  ( .D(n989), .E(\u_outFIFO/n410 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[16][3] ) );
  DFE1 \u_outFIFO/FIFO_reg[17][0]  ( .D(n989), .E(\u_outFIFO/n412 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[17][0] ) );
  DFE1 \u_outFIFO/FIFO_reg[17][1]  ( .D(n989), .E(\u_outFIFO/n413 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[17][1] ) );
  DFE1 \u_outFIFO/FIFO_reg[17][2]  ( .D(n989), .E(\u_outFIFO/n414 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[17][2] ) );
  DFE1 \u_outFIFO/FIFO_reg[17][3]  ( .D(n989), .E(\u_outFIFO/n415 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[17][3] ) );
  DFE1 \u_outFIFO/FIFO_reg[19][0]  ( .D(n990), .E(\u_outFIFO/n420 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[19][0] ) );
  DFE1 \u_outFIFO/FIFO_reg[19][1]  ( .D(n990), .E(\u_outFIFO/n421 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[19][1] ) );
  DFE1 \u_outFIFO/FIFO_reg[19][2]  ( .D(n990), .E(\u_outFIFO/n422 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[19][2] ) );
  DFE1 \u_outFIFO/FIFO_reg[19][3]  ( .D(n990), .E(\u_outFIFO/n423 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[19][3] ) );
  DFE1 \u_outFIFO/FIFO_reg[20][0]  ( .D(n991), .E(\u_outFIFO/n424 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[20][0] ) );
  DFE1 \u_outFIFO/FIFO_reg[20][1]  ( .D(n991), .E(\u_outFIFO/n425 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[20][1] ) );
  DFE1 \u_outFIFO/FIFO_reg[20][2]  ( .D(n991), .E(\u_outFIFO/n426 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[20][2] ) );
  DFE1 \u_outFIFO/FIFO_reg[20][3]  ( .D(n991), .E(\u_outFIFO/n427 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[20][3] ) );
  DFE1 \u_outFIFO/FIFO_reg[21][0]  ( .D(n991), .E(\u_outFIFO/n428 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[21][0] ) );
  DFE1 \u_outFIFO/FIFO_reg[21][1]  ( .D(n991), .E(\u_outFIFO/n429 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[21][1] ) );
  DFE1 \u_outFIFO/FIFO_reg[21][2]  ( .D(n991), .E(\u_outFIFO/n430 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[21][2] ) );
  DFE1 \u_outFIFO/FIFO_reg[21][3]  ( .D(n991), .E(\u_outFIFO/n431 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[21][3] ) );
  DFE1 \u_outFIFO/FIFO_reg[23][0]  ( .D(n992), .E(\u_outFIFO/n436 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[23][0] ) );
  DFE1 \u_outFIFO/FIFO_reg[23][1]  ( .D(n992), .E(\u_outFIFO/n437 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[23][1] ) );
  DFE1 \u_outFIFO/FIFO_reg[23][2]  ( .D(n992), .E(\u_outFIFO/n438 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[23][2] ) );
  DFE1 \u_outFIFO/FIFO_reg[23][3]  ( .D(n992), .E(\u_outFIFO/n439 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[23][3] ) );
  DFE1 \u_outFIFO/FIFO_reg[24][0]  ( .D(n993), .E(\u_outFIFO/n440 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[24][0] ) );
  DFE1 \u_outFIFO/FIFO_reg[24][1]  ( .D(n993), .E(\u_outFIFO/n441 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[24][1] ) );
  DFE1 \u_outFIFO/FIFO_reg[24][2]  ( .D(n993), .E(\u_outFIFO/n442 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[24][2] ) );
  DFE1 \u_outFIFO/FIFO_reg[24][3]  ( .D(n993), .E(\u_outFIFO/n443 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[24][3] ) );
  DFE1 \u_outFIFO/FIFO_reg[25][0]  ( .D(n993), .E(\u_outFIFO/n444 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[25][0] ) );
  DFE1 \u_outFIFO/FIFO_reg[25][1]  ( .D(n993), .E(\u_outFIFO/n445 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[25][1] ) );
  DFE1 \u_outFIFO/FIFO_reg[25][2]  ( .D(n993), .E(\u_outFIFO/n446 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[25][2] ) );
  DFE1 \u_outFIFO/FIFO_reg[25][3]  ( .D(n993), .E(\u_outFIFO/n447 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[25][3] ) );
  DFE1 \u_outFIFO/FIFO_reg[27][0]  ( .D(n994), .E(\u_outFIFO/n452 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[27][0] ) );
  DFE1 \u_outFIFO/FIFO_reg[27][1]  ( .D(n994), .E(\u_outFIFO/n453 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[27][1] ) );
  DFE1 \u_outFIFO/FIFO_reg[27][2]  ( .D(n994), .E(\u_outFIFO/n454 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[27][2] ) );
  DFE1 \u_outFIFO/FIFO_reg[27][3]  ( .D(n994), .E(\u_outFIFO/n455 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[27][3] ) );
  DFE1 \u_outFIFO/FIFO_reg[28][0]  ( .D(n995), .E(\u_outFIFO/n456 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[28][0] ) );
  DFE1 \u_outFIFO/FIFO_reg[28][1]  ( .D(n995), .E(\u_outFIFO/n457 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[28][1] ) );
  DFE1 \u_outFIFO/FIFO_reg[28][2]  ( .D(n995), .E(\u_outFIFO/n458 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[28][2] ) );
  DFE1 \u_outFIFO/FIFO_reg[28][3]  ( .D(n995), .E(\u_outFIFO/n459 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[28][3] ) );
  DFE1 \u_outFIFO/FIFO_reg[29][0]  ( .D(n995), .E(\u_outFIFO/n460 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[29][0] ) );
  DFE1 \u_outFIFO/FIFO_reg[29][1]  ( .D(n995), .E(\u_outFIFO/n461 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[29][1] ) );
  DFE1 \u_outFIFO/FIFO_reg[29][2]  ( .D(n995), .E(\u_outFIFO/n462 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[29][2] ) );
  DFE1 \u_outFIFO/FIFO_reg[29][3]  ( .D(n995), .E(\u_outFIFO/n463 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[29][3] ) );
  DFE1 \u_outFIFO/FIFO_reg[31][0]  ( .D(n996), .E(\u_outFIFO/n468 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[31][0] ) );
  DFE1 \u_outFIFO/FIFO_reg[31][1]  ( .D(n996), .E(\u_outFIFO/n470 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[31][1] ) );
  DFE1 \u_outFIFO/FIFO_reg[31][2]  ( .D(n996), .E(\u_outFIFO/n471 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[31][2] ) );
  DFE1 \u_outFIFO/FIFO_reg[31][3]  ( .D(n996), .E(\u_outFIFO/n472 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[31][3] ) );
  DFE1 \u_outFIFO/FIFO_reg[32][0]  ( .D(n997), .E(\u_outFIFO/n473 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[32][0] ) );
  DFE1 \u_outFIFO/FIFO_reg[32][1]  ( .D(n997), .E(\u_outFIFO/n475 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[32][1] ) );
  DFE1 \u_outFIFO/FIFO_reg[32][2]  ( .D(n997), .E(\u_outFIFO/n477 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[32][2] ) );
  DFE1 \u_outFIFO/FIFO_reg[32][3]  ( .D(n997), .E(\u_outFIFO/n479 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[32][3] ) );
  DFE1 \u_outFIFO/FIFO_reg[33][0]  ( .D(n997), .E(\u_outFIFO/n481 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[33][0] ) );
  DFE1 \u_outFIFO/FIFO_reg[33][1]  ( .D(n997), .E(\u_outFIFO/n482 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[33][1] ) );
  DFE1 \u_outFIFO/FIFO_reg[33][2]  ( .D(n997), .E(\u_outFIFO/n483 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[33][2] ) );
  DFE1 \u_outFIFO/FIFO_reg[33][3]  ( .D(n997), .E(\u_outFIFO/n484 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[33][3] ) );
  DFE1 \u_outFIFO/FIFO_reg[35][0]  ( .D(n998), .E(\u_outFIFO/n489 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[35][0] ) );
  DFE1 \u_outFIFO/FIFO_reg[35][1]  ( .D(n998), .E(\u_outFIFO/n490 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[35][1] ) );
  DFE1 \u_outFIFO/FIFO_reg[35][2]  ( .D(n998), .E(\u_outFIFO/n491 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[35][2] ) );
  DFE1 \u_outFIFO/FIFO_reg[35][3]  ( .D(n998), .E(\u_outFIFO/n492 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[35][3] ) );
  DFE1 \u_outFIFO/FIFO_reg[36][0]  ( .D(n999), .E(\u_outFIFO/n493 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[36][0] ) );
  DFE1 \u_outFIFO/FIFO_reg[36][1]  ( .D(n999), .E(\u_outFIFO/n494 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[36][1] ) );
  DFE1 \u_outFIFO/FIFO_reg[36][2]  ( .D(n999), .E(\u_outFIFO/n495 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[36][2] ) );
  DFE1 \u_outFIFO/FIFO_reg[36][3]  ( .D(n999), .E(\u_outFIFO/n496 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[36][3] ) );
  DFE1 \u_outFIFO/FIFO_reg[37][0]  ( .D(n999), .E(\u_outFIFO/n497 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[37][0] ) );
  DFE1 \u_outFIFO/FIFO_reg[37][1]  ( .D(n999), .E(\u_outFIFO/n498 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[37][1] ) );
  DFE1 \u_outFIFO/FIFO_reg[37][2]  ( .D(n999), .E(\u_outFIFO/n499 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[37][2] ) );
  DFE1 \u_outFIFO/FIFO_reg[37][3]  ( .D(n999), .E(\u_outFIFO/n500 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[37][3] ) );
  DFE1 \u_outFIFO/FIFO_reg[39][0]  ( .D(n1000), .E(\u_outFIFO/n505 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[39][0] ) );
  DFE1 \u_outFIFO/FIFO_reg[39][1]  ( .D(n1000), .E(\u_outFIFO/n506 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[39][1] ) );
  DFE1 \u_outFIFO/FIFO_reg[39][2]  ( .D(n1000), .E(\u_outFIFO/n507 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[39][2] ) );
  DFE1 \u_outFIFO/FIFO_reg[39][3]  ( .D(n1000), .E(\u_outFIFO/n508 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[39][3] ) );
  DFE1 \u_outFIFO/FIFO_reg[40][0]  ( .D(n1001), .E(\u_outFIFO/n509 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[40][0] ) );
  DFE1 \u_outFIFO/FIFO_reg[40][1]  ( .D(n1001), .E(\u_outFIFO/n510 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[40][1] ) );
  DFE1 \u_outFIFO/FIFO_reg[40][2]  ( .D(n1001), .E(\u_outFIFO/n511 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[40][2] ) );
  DFE1 \u_outFIFO/FIFO_reg[40][3]  ( .D(n1001), .E(\u_outFIFO/n512 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[40][3] ) );
  DFE1 \u_outFIFO/FIFO_reg[41][0]  ( .D(n1001), .E(\u_outFIFO/n513 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[41][0] ) );
  DFE1 \u_outFIFO/FIFO_reg[41][1]  ( .D(n1001), .E(\u_outFIFO/n514 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[41][1] ) );
  DFE1 \u_outFIFO/FIFO_reg[41][2]  ( .D(n1001), .E(\u_outFIFO/n515 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[41][2] ) );
  DFE1 \u_outFIFO/FIFO_reg[41][3]  ( .D(n1001), .E(\u_outFIFO/n516 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[41][3] ) );
  DFE1 \u_outFIFO/FIFO_reg[43][0]  ( .D(n1002), .E(\u_outFIFO/n521 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[43][0] ) );
  DFE1 \u_outFIFO/FIFO_reg[43][1]  ( .D(n1002), .E(\u_outFIFO/n522 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[43][1] ) );
  DFE1 \u_outFIFO/FIFO_reg[43][2]  ( .D(n1002), .E(\u_outFIFO/n523 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[43][2] ) );
  DFE1 \u_outFIFO/FIFO_reg[43][3]  ( .D(n1002), .E(\u_outFIFO/n524 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[43][3] ) );
  DFE1 \u_outFIFO/FIFO_reg[44][0]  ( .D(n1003), .E(\u_outFIFO/n525 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[44][0] ) );
  DFE1 \u_outFIFO/FIFO_reg[44][1]  ( .D(n1003), .E(\u_outFIFO/n526 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[44][1] ) );
  DFE1 \u_outFIFO/FIFO_reg[44][2]  ( .D(n1003), .E(\u_outFIFO/n527 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[44][2] ) );
  DFE1 \u_outFIFO/FIFO_reg[44][3]  ( .D(n1003), .E(\u_outFIFO/n528 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[44][3] ) );
  DFE1 \u_outFIFO/FIFO_reg[45][0]  ( .D(n1003), .E(\u_outFIFO/n529 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[45][0] ) );
  DFE1 \u_outFIFO/FIFO_reg[45][1]  ( .D(n1003), .E(\u_outFIFO/n530 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[45][1] ) );
  DFE1 \u_outFIFO/FIFO_reg[45][2]  ( .D(n1003), .E(\u_outFIFO/n531 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[45][2] ) );
  DFE1 \u_outFIFO/FIFO_reg[45][3]  ( .D(n1003), .E(\u_outFIFO/n532 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[45][3] ) );
  DFE1 \u_outFIFO/FIFO_reg[47][0]  ( .D(n1004), .E(\u_outFIFO/n537 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[47][0] ) );
  DFE1 \u_outFIFO/FIFO_reg[47][1]  ( .D(n1004), .E(\u_outFIFO/n539 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[47][1] ) );
  DFE1 \u_outFIFO/FIFO_reg[47][2]  ( .D(n1004), .E(\u_outFIFO/n540 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[47][2] ) );
  DFE1 \u_outFIFO/FIFO_reg[47][3]  ( .D(n1004), .E(\u_outFIFO/n541 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[47][3] ) );
  DFE1 \u_outFIFO/FIFO_reg[48][0]  ( .D(n1005), .E(\u_outFIFO/n542 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[48][0] ) );
  DFE1 \u_outFIFO/FIFO_reg[48][1]  ( .D(n1005), .E(\u_outFIFO/n544 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[48][1] ) );
  DFE1 \u_outFIFO/FIFO_reg[48][2]  ( .D(n1005), .E(\u_outFIFO/n546 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[48][2] ) );
  DFE1 \u_outFIFO/FIFO_reg[48][3]  ( .D(n1005), .E(\u_outFIFO/n548 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[48][3] ) );
  DFE1 \u_outFIFO/FIFO_reg[49][0]  ( .D(n1005), .E(\u_outFIFO/n550 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[49][0] ) );
  DFE1 \u_outFIFO/FIFO_reg[49][1]  ( .D(n1005), .E(\u_outFIFO/n551 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[49][1] ) );
  DFE1 \u_outFIFO/FIFO_reg[49][2]  ( .D(n1005), .E(\u_outFIFO/n552 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[49][2] ) );
  DFE1 \u_outFIFO/FIFO_reg[49][3]  ( .D(n1005), .E(\u_outFIFO/n553 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[49][3] ) );
  DFE1 \u_outFIFO/FIFO_reg[51][0]  ( .D(n1006), .E(\u_outFIFO/n558 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[51][0] ) );
  DFE1 \u_outFIFO/FIFO_reg[51][1]  ( .D(n1006), .E(\u_outFIFO/n559 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[51][1] ) );
  DFE1 \u_outFIFO/FIFO_reg[51][2]  ( .D(n1006), .E(\u_outFIFO/n560 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[51][2] ) );
  DFE1 \u_outFIFO/FIFO_reg[51][3]  ( .D(n1006), .E(\u_outFIFO/n561 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[51][3] ) );
  DFE1 \u_outFIFO/FIFO_reg[52][0]  ( .D(n1007), .E(\u_outFIFO/n562 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[52][0] ) );
  DFE1 \u_outFIFO/FIFO_reg[52][1]  ( .D(n1007), .E(\u_outFIFO/n563 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[52][1] ) );
  DFE1 \u_outFIFO/FIFO_reg[52][2]  ( .D(n1007), .E(\u_outFIFO/n564 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[52][2] ) );
  DFE1 \u_outFIFO/FIFO_reg[52][3]  ( .D(n1007), .E(\u_outFIFO/n565 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[52][3] ) );
  DFE1 \u_outFIFO/FIFO_reg[53][0]  ( .D(n1007), .E(\u_outFIFO/n566 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[53][0] ) );
  DFE1 \u_outFIFO/FIFO_reg[53][1]  ( .D(n1007), .E(\u_outFIFO/n567 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[53][1] ) );
  DFE1 \u_outFIFO/FIFO_reg[53][2]  ( .D(n1007), .E(\u_outFIFO/n568 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[53][2] ) );
  DFE1 \u_outFIFO/FIFO_reg[53][3]  ( .D(n1007), .E(\u_outFIFO/n569 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[53][3] ) );
  DFE1 \u_outFIFO/FIFO_reg[55][0]  ( .D(n1008), .E(\u_outFIFO/n574 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[55][0] ) );
  DFE1 \u_outFIFO/FIFO_reg[55][1]  ( .D(n1008), .E(\u_outFIFO/n575 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[55][1] ) );
  DFE1 \u_outFIFO/FIFO_reg[55][2]  ( .D(n1008), .E(\u_outFIFO/n576 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[55][2] ) );
  DFE1 \u_outFIFO/FIFO_reg[55][3]  ( .D(n1008), .E(\u_outFIFO/n577 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[55][3] ) );
  DFE1 \u_outFIFO/FIFO_reg[56][0]  ( .D(n1009), .E(\u_outFIFO/n578 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[56][0] ) );
  DFE1 \u_outFIFO/FIFO_reg[56][1]  ( .D(n1009), .E(\u_outFIFO/n579 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[56][1] ) );
  DFE1 \u_outFIFO/FIFO_reg[56][2]  ( .D(n1009), .E(\u_outFIFO/n580 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[56][2] ) );
  DFE1 \u_outFIFO/FIFO_reg[56][3]  ( .D(n1009), .E(\u_outFIFO/n581 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[56][3] ) );
  DFE1 \u_outFIFO/FIFO_reg[57][0]  ( .D(n1009), .E(\u_outFIFO/n582 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[57][0] ) );
  DFE1 \u_outFIFO/FIFO_reg[57][1]  ( .D(n1009), .E(\u_outFIFO/n583 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[57][1] ) );
  DFE1 \u_outFIFO/FIFO_reg[57][2]  ( .D(n1009), .E(\u_outFIFO/n584 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[57][2] ) );
  DFE1 \u_outFIFO/FIFO_reg[57][3]  ( .D(n1009), .E(\u_outFIFO/n585 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[57][3] ) );
  DFE1 \u_outFIFO/FIFO_reg[59][0]  ( .D(n1010), .E(\u_outFIFO/n590 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[59][0] ) );
  DFE1 \u_outFIFO/FIFO_reg[59][1]  ( .D(n1010), .E(\u_outFIFO/n591 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[59][1] ) );
  DFE1 \u_outFIFO/FIFO_reg[59][2]  ( .D(n1010), .E(\u_outFIFO/n592 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[59][2] ) );
  DFE1 \u_outFIFO/FIFO_reg[59][3]  ( .D(n1010), .E(\u_outFIFO/n593 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[59][3] ) );
  DFE1 \u_outFIFO/FIFO_reg[60][0]  ( .D(n1011), .E(\u_outFIFO/n594 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[60][0] ) );
  DFE1 \u_outFIFO/FIFO_reg[60][1]  ( .D(n1011), .E(\u_outFIFO/n595 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[60][1] ) );
  DFE1 \u_outFIFO/FIFO_reg[60][2]  ( .D(n1011), .E(\u_outFIFO/n596 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[60][2] ) );
  DFE1 \u_outFIFO/FIFO_reg[60][3]  ( .D(n1011), .E(\u_outFIFO/n597 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[60][3] ) );
  DFE1 \u_outFIFO/FIFO_reg[61][0]  ( .D(n1011), .E(\u_outFIFO/n598 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[61][0] ) );
  DFE1 \u_outFIFO/FIFO_reg[61][1]  ( .D(n1011), .E(\u_outFIFO/n599 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[61][1] ) );
  DFE1 \u_outFIFO/FIFO_reg[61][2]  ( .D(n1011), .E(\u_outFIFO/n600 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[61][2] ) );
  DFE1 \u_outFIFO/FIFO_reg[61][3]  ( .D(n1011), .E(\u_outFIFO/n601 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[61][3] ) );
  DFE1 \u_outFIFO/FIFO_reg[63][0]  ( .D(n1012), .E(\u_outFIFO/n606 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[63][0] ) );
  DFE1 \u_outFIFO/FIFO_reg[63][1]  ( .D(n1012), .E(\u_outFIFO/n608 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[63][1] ) );
  DFE1 \u_outFIFO/FIFO_reg[63][2]  ( .D(n1012), .E(\u_outFIFO/n609 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[63][2] ) );
  DFE1 \u_outFIFO/FIFO_reg[63][3]  ( .D(n1012), .E(\u_outFIFO/n610 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[63][3] ) );
  DFE1 \u_outFIFO/FIFO_reg[64][0]  ( .D(n1013), .E(\u_outFIFO/n611 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[64][0] ) );
  DFE1 \u_outFIFO/FIFO_reg[64][1]  ( .D(n1013), .E(\u_outFIFO/n613 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[64][1] ) );
  DFE1 \u_outFIFO/FIFO_reg[64][2]  ( .D(n1013), .E(\u_outFIFO/n615 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[64][2] ) );
  DFE1 \u_outFIFO/FIFO_reg[64][3]  ( .D(n1013), .E(\u_outFIFO/n617 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[64][3] ) );
  DFE1 \u_outFIFO/FIFO_reg[65][0]  ( .D(n1013), .E(\u_outFIFO/n619 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[65][0] ) );
  DFE1 \u_outFIFO/FIFO_reg[65][1]  ( .D(n1013), .E(\u_outFIFO/n620 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[65][1] ) );
  DFE1 \u_outFIFO/FIFO_reg[65][2]  ( .D(n1013), .E(\u_outFIFO/n621 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[65][2] ) );
  DFE1 \u_outFIFO/FIFO_reg[65][3]  ( .D(n1013), .E(\u_outFIFO/n622 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[65][3] ) );
  DFE1 \u_outFIFO/FIFO_reg[67][0]  ( .D(n1014), .E(\u_outFIFO/n627 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[67][0] ) );
  DFE1 \u_outFIFO/FIFO_reg[67][1]  ( .D(n1014), .E(\u_outFIFO/n628 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[67][1] ) );
  DFE1 \u_outFIFO/FIFO_reg[67][2]  ( .D(n1014), .E(\u_outFIFO/n629 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[67][2] ) );
  DFE1 \u_outFIFO/FIFO_reg[67][3]  ( .D(n1014), .E(\u_outFIFO/n630 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[67][3] ) );
  DFE1 \u_outFIFO/FIFO_reg[68][0]  ( .D(n1015), .E(\u_outFIFO/n631 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[68][0] ) );
  DFE1 \u_outFIFO/FIFO_reg[68][1]  ( .D(n1015), .E(\u_outFIFO/n632 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[68][1] ) );
  DFE1 \u_outFIFO/FIFO_reg[68][2]  ( .D(n1015), .E(\u_outFIFO/n633 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[68][2] ) );
  DFE1 \u_outFIFO/FIFO_reg[68][3]  ( .D(n1015), .E(\u_outFIFO/n634 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[68][3] ) );
  DFE1 \u_outFIFO/FIFO_reg[69][0]  ( .D(n1015), .E(\u_outFIFO/n635 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[69][0] ) );
  DFE1 \u_outFIFO/FIFO_reg[69][1]  ( .D(n1015), .E(\u_outFIFO/n636 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[69][1] ) );
  DFE1 \u_outFIFO/FIFO_reg[69][2]  ( .D(n1015), .E(\u_outFIFO/n637 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[69][2] ) );
  DFE1 \u_outFIFO/FIFO_reg[69][3]  ( .D(n1015), .E(\u_outFIFO/n638 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[69][3] ) );
  DFE1 \u_outFIFO/FIFO_reg[71][0]  ( .D(n1016), .E(\u_outFIFO/n643 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[71][0] ) );
  DFE1 \u_outFIFO/FIFO_reg[71][1]  ( .D(n1016), .E(\u_outFIFO/n644 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[71][1] ) );
  DFE1 \u_outFIFO/FIFO_reg[71][2]  ( .D(n1016), .E(\u_outFIFO/n645 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[71][2] ) );
  DFE1 \u_outFIFO/FIFO_reg[71][3]  ( .D(n1016), .E(\u_outFIFO/n646 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[71][3] ) );
  DFE1 \u_outFIFO/FIFO_reg[72][0]  ( .D(n1017), .E(\u_outFIFO/n647 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[72][0] ) );
  DFE1 \u_outFIFO/FIFO_reg[72][1]  ( .D(n1017), .E(\u_outFIFO/n648 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[72][1] ) );
  DFE1 \u_outFIFO/FIFO_reg[72][2]  ( .D(n1017), .E(\u_outFIFO/n649 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[72][2] ) );
  DFE1 \u_outFIFO/FIFO_reg[72][3]  ( .D(n1017), .E(\u_outFIFO/n650 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[72][3] ) );
  DFE1 \u_outFIFO/FIFO_reg[73][0]  ( .D(n1017), .E(\u_outFIFO/n651 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[73][0] ) );
  DFE1 \u_outFIFO/FIFO_reg[73][1]  ( .D(n1017), .E(\u_outFIFO/n652 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[73][1] ) );
  DFE1 \u_outFIFO/FIFO_reg[73][2]  ( .D(n1017), .E(\u_outFIFO/n653 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[73][2] ) );
  DFE1 \u_outFIFO/FIFO_reg[73][3]  ( .D(n1017), .E(\u_outFIFO/n654 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[73][3] ) );
  DFE1 \u_outFIFO/FIFO_reg[75][0]  ( .D(n1018), .E(\u_outFIFO/n662 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[75][0] ) );
  DFE1 \u_outFIFO/FIFO_reg[75][1]  ( .D(n1018), .E(\u_outFIFO/n663 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[75][1] ) );
  DFE1 \u_outFIFO/FIFO_reg[75][2]  ( .D(n1018), .E(\u_outFIFO/n665 ), .C(
        inClock), .Q(\u_outFIFO/FIFO[75][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[2][0]  ( .D(n1019), .E(n2091), .C(inClock), .Q(
        \u_inFIFO/FIFO[2][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[2][1]  ( .D(n1035), .E(n2091), .C(inClock), .Q(
        \u_inFIFO/FIFO[2][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[2][2]  ( .D(n1051), .E(n2091), .C(inClock), .Q(
        \u_inFIFO/FIFO[2][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[2][3]  ( .D(n1067), .E(n2091), .C(inClock), .Q(
        \u_inFIFO/FIFO[2][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[6][0]  ( .D(n1019), .E(n2087), .C(inClock), .Q(
        \u_inFIFO/FIFO[6][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[6][1]  ( .D(n1035), .E(n2087), .C(inClock), .Q(
        \u_inFIFO/FIFO[6][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[6][2]  ( .D(n1051), .E(n2087), .C(inClock), .Q(
        \u_inFIFO/FIFO[6][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[6][3]  ( .D(n1067), .E(n2087), .C(inClock), .Q(
        \u_inFIFO/FIFO[6][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[10][0]  ( .D(n1020), .E(n2083), .C(inClock), .Q(
        \u_inFIFO/FIFO[10][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[10][1]  ( .D(n1036), .E(n2083), .C(inClock), .Q(
        \u_inFIFO/FIFO[10][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[10][2]  ( .D(n1052), .E(n2083), .C(inClock), .Q(
        \u_inFIFO/FIFO[10][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[10][3]  ( .D(n1068), .E(n2083), .C(inClock), .Q(
        \u_inFIFO/FIFO[10][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[14][0]  ( .D(n1020), .E(n2079), .C(inClock), .Q(
        \u_inFIFO/FIFO[14][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[14][1]  ( .D(n1036), .E(n2079), .C(inClock), .Q(
        \u_inFIFO/FIFO[14][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[14][2]  ( .D(n1052), .E(n2079), .C(inClock), .Q(
        \u_inFIFO/FIFO[14][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[14][3]  ( .D(n1068), .E(n2079), .C(inClock), .Q(
        \u_inFIFO/FIFO[14][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[18][0]  ( .D(n1021), .E(n2075), .C(inClock), .Q(
        \u_inFIFO/FIFO[18][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[18][1]  ( .D(n1037), .E(n2075), .C(inClock), .Q(
        \u_inFIFO/FIFO[18][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[18][2]  ( .D(n1053), .E(n2075), .C(inClock), .Q(
        \u_inFIFO/FIFO[18][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[18][3]  ( .D(n1069), .E(n2075), .C(inClock), .Q(
        \u_inFIFO/FIFO[18][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[22][0]  ( .D(n1021), .E(n2071), .C(inClock), .Q(
        \u_inFIFO/FIFO[22][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[22][1]  ( .D(n1037), .E(n2071), .C(inClock), .Q(
        \u_inFIFO/FIFO[22][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[22][2]  ( .D(n1053), .E(n2071), .C(inClock), .Q(
        \u_inFIFO/FIFO[22][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[22][3]  ( .D(n1069), .E(n2071), .C(inClock), .Q(
        \u_inFIFO/FIFO[22][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[26][0]  ( .D(n1022), .E(n2067), .C(inClock), .Q(
        \u_inFIFO/FIFO[26][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[26][1]  ( .D(n1038), .E(n2067), .C(inClock), .Q(
        \u_inFIFO/FIFO[26][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[26][2]  ( .D(n1054), .E(n2067), .C(inClock), .Q(
        \u_inFIFO/FIFO[26][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[26][3]  ( .D(n1070), .E(n2067), .C(inClock), .Q(
        \u_inFIFO/FIFO[26][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[30][0]  ( .D(n1022), .E(n2063), .C(inClock), .Q(
        \u_inFIFO/FIFO[30][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[30][1]  ( .D(n1038), .E(n2063), .C(inClock), .Q(
        \u_inFIFO/FIFO[30][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[30][2]  ( .D(n1054), .E(n2063), .C(inClock), .Q(
        \u_inFIFO/FIFO[30][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[30][3]  ( .D(n1070), .E(n2063), .C(inClock), .Q(
        \u_inFIFO/FIFO[30][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[34][0]  ( .D(n1023), .E(n2059), .C(inClock), .Q(
        \u_inFIFO/FIFO[34][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[34][1]  ( .D(n1039), .E(n2059), .C(inClock), .Q(
        \u_inFIFO/FIFO[34][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[34][2]  ( .D(n1055), .E(n2059), .C(inClock), .Q(
        \u_inFIFO/FIFO[34][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[34][3]  ( .D(n1071), .E(n2059), .C(inClock), .Q(
        \u_inFIFO/FIFO[34][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[38][0]  ( .D(n1023), .E(n2055), .C(inClock), .Q(
        \u_inFIFO/FIFO[38][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[38][1]  ( .D(n1039), .E(n2055), .C(inClock), .Q(
        \u_inFIFO/FIFO[38][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[38][2]  ( .D(n1055), .E(n2055), .C(inClock), .Q(
        \u_inFIFO/FIFO[38][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[38][3]  ( .D(n1071), .E(n2055), .C(inClock), .Q(
        \u_inFIFO/FIFO[38][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[42][0]  ( .D(n1024), .E(n2051), .C(inClock), .Q(
        \u_inFIFO/FIFO[42][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[42][1]  ( .D(n1040), .E(n2051), .C(inClock), .Q(
        \u_inFIFO/FIFO[42][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[42][2]  ( .D(n1056), .E(n2051), .C(inClock), .Q(
        \u_inFIFO/FIFO[42][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[42][3]  ( .D(n1072), .E(n2051), .C(inClock), .Q(
        \u_inFIFO/FIFO[42][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[46][0]  ( .D(n1024), .E(n2047), .C(inClock), .Q(
        \u_inFIFO/FIFO[46][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[46][1]  ( .D(n1040), .E(n2047), .C(inClock), .Q(
        \u_inFIFO/FIFO[46][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[46][2]  ( .D(n1056), .E(n2047), .C(inClock), .Q(
        \u_inFIFO/FIFO[46][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[46][3]  ( .D(n1072), .E(n2047), .C(inClock), .Q(
        \u_inFIFO/FIFO[46][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[50][0]  ( .D(n1025), .E(n2043), .C(inClock), .Q(
        \u_inFIFO/FIFO[50][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[50][1]  ( .D(n1041), .E(n2043), .C(inClock), .Q(
        \u_inFIFO/FIFO[50][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[50][2]  ( .D(n1057), .E(n2043), .C(inClock), .Q(
        \u_inFIFO/FIFO[50][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[50][3]  ( .D(n1073), .E(n2043), .C(inClock), .Q(
        \u_inFIFO/FIFO[50][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[54][0]  ( .D(n1025), .E(n2039), .C(inClock), .Q(
        \u_inFIFO/FIFO[54][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[54][1]  ( .D(n1041), .E(n2039), .C(inClock), .Q(
        \u_inFIFO/FIFO[54][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[54][2]  ( .D(n1057), .E(n2039), .C(inClock), .Q(
        \u_inFIFO/FIFO[54][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[54][3]  ( .D(n1073), .E(n2039), .C(inClock), .Q(
        \u_inFIFO/FIFO[54][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[58][0]  ( .D(n1026), .E(n2035), .C(inClock), .Q(
        \u_inFIFO/FIFO[58][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[58][1]  ( .D(n1042), .E(n2035), .C(inClock), .Q(
        \u_inFIFO/FIFO[58][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[58][2]  ( .D(n1058), .E(n2035), .C(inClock), .Q(
        \u_inFIFO/FIFO[58][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[58][3]  ( .D(n1074), .E(n2035), .C(inClock), .Q(
        \u_inFIFO/FIFO[58][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[62][0]  ( .D(n1026), .E(n2031), .C(inClock), .Q(
        \u_inFIFO/FIFO[62][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[62][1]  ( .D(n1042), .E(n2031), .C(inClock), .Q(
        \u_inFIFO/FIFO[62][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[62][2]  ( .D(n1058), .E(n2031), .C(inClock), .Q(
        \u_inFIFO/FIFO[62][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[62][3]  ( .D(n1074), .E(n2031), .C(inClock), .Q(
        \u_inFIFO/FIFO[62][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[66][0]  ( .D(n1027), .E(n2027), .C(inClock), .Q(
        \u_inFIFO/FIFO[66][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[66][1]  ( .D(n1043), .E(n2027), .C(inClock), .Q(
        \u_inFIFO/FIFO[66][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[66][2]  ( .D(n1059), .E(n2027), .C(inClock), .Q(
        \u_inFIFO/FIFO[66][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[66][3]  ( .D(n1075), .E(n2027), .C(inClock), .Q(
        \u_inFIFO/FIFO[66][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[70][0]  ( .D(n1027), .E(n2023), .C(inClock), .Q(
        \u_inFIFO/FIFO[70][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[70][1]  ( .D(n1043), .E(n2023), .C(inClock), .Q(
        \u_inFIFO/FIFO[70][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[70][2]  ( .D(n1059), .E(n2023), .C(inClock), .Q(
        \u_inFIFO/FIFO[70][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[70][3]  ( .D(n1075), .E(n2023), .C(inClock), .Q(
        \u_inFIFO/FIFO[70][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[74][0]  ( .D(n1028), .E(n2019), .C(inClock), .Q(
        \u_inFIFO/FIFO[74][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[74][1]  ( .D(n1044), .E(n2019), .C(inClock), .Q(
        \u_inFIFO/FIFO[74][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[74][2]  ( .D(n1060), .E(n2019), .C(inClock), .Q(
        \u_inFIFO/FIFO[74][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[74][3]  ( .D(n1076), .E(n2019), .C(inClock), .Q(
        \u_inFIFO/FIFO[74][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[78][0]  ( .D(n1028), .E(n2015), .C(inClock), .Q(
        \u_inFIFO/FIFO[78][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[78][1]  ( .D(n1044), .E(n2015), .C(inClock), .Q(
        \u_inFIFO/FIFO[78][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[78][2]  ( .D(n1060), .E(n2015), .C(inClock), .Q(
        \u_inFIFO/FIFO[78][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[78][3]  ( .D(n1076), .E(n2015), .C(inClock), .Q(
        \u_inFIFO/FIFO[78][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[82][0]  ( .D(n1029), .E(n2011), .C(inClock), .Q(
        \u_inFIFO/FIFO[82][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[82][1]  ( .D(n1045), .E(n2011), .C(inClock), .Q(
        \u_inFIFO/FIFO[82][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[82][2]  ( .D(n1061), .E(n2011), .C(inClock), .Q(
        \u_inFIFO/FIFO[82][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[82][3]  ( .D(n1077), .E(n2011), .C(inClock), .Q(
        \u_inFIFO/FIFO[82][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[86][0]  ( .D(n1029), .E(n2007), .C(inClock), .Q(
        \u_inFIFO/FIFO[86][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[86][1]  ( .D(n1045), .E(n2007), .C(inClock), .Q(
        \u_inFIFO/FIFO[86][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[86][2]  ( .D(n1061), .E(n2007), .C(inClock), .Q(
        \u_inFIFO/FIFO[86][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[86][3]  ( .D(n1077), .E(n2007), .C(inClock), .Q(
        \u_inFIFO/FIFO[86][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[90][0]  ( .D(n1030), .E(n2003), .C(inClock), .Q(
        \u_inFIFO/FIFO[90][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[90][1]  ( .D(n1046), .E(n2003), .C(inClock), .Q(
        \u_inFIFO/FIFO[90][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[90][2]  ( .D(n1062), .E(n2003), .C(inClock), .Q(
        \u_inFIFO/FIFO[90][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[90][3]  ( .D(n1078), .E(n2003), .C(inClock), .Q(
        \u_inFIFO/FIFO[90][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[94][0]  ( .D(n1030), .E(n1999), .C(inClock), .Q(
        \u_inFIFO/FIFO[94][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[94][1]  ( .D(n1046), .E(n1999), .C(inClock), .Q(
        \u_inFIFO/FIFO[94][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[94][2]  ( .D(n1062), .E(n1999), .C(inClock), .Q(
        \u_inFIFO/FIFO[94][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[94][3]  ( .D(n1078), .E(n1999), .C(inClock), .Q(
        \u_inFIFO/FIFO[94][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[98][0]  ( .D(n1031), .E(n1995), .C(inClock), .Q(
        \u_inFIFO/FIFO[98][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[98][1]  ( .D(n1047), .E(n1995), .C(inClock), .Q(
        \u_inFIFO/FIFO[98][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[98][2]  ( .D(n1063), .E(n1995), .C(inClock), .Q(
        \u_inFIFO/FIFO[98][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[98][3]  ( .D(n1079), .E(n1995), .C(inClock), .Q(
        \u_inFIFO/FIFO[98][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[102][0]  ( .D(n1031), .E(n1991), .C(inClock), .Q(
        \u_inFIFO/FIFO[102][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[102][1]  ( .D(n1047), .E(n1991), .C(inClock), .Q(
        \u_inFIFO/FIFO[102][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[102][2]  ( .D(n1063), .E(n1991), .C(inClock), .Q(
        \u_inFIFO/FIFO[102][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[102][3]  ( .D(n1079), .E(n1991), .C(inClock), .Q(
        \u_inFIFO/FIFO[102][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[106][0]  ( .D(n1032), .E(n1987), .C(inClock), .Q(
        \u_inFIFO/FIFO[106][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[106][1]  ( .D(n1048), .E(n1987), .C(inClock), .Q(
        \u_inFIFO/FIFO[106][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[106][2]  ( .D(n1064), .E(n1987), .C(inClock), .Q(
        \u_inFIFO/FIFO[106][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[106][3]  ( .D(n1080), .E(n1987), .C(inClock), .Q(
        \u_inFIFO/FIFO[106][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[110][0]  ( .D(n1032), .E(n1983), .C(inClock), .Q(
        \u_inFIFO/FIFO[110][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[110][1]  ( .D(n1048), .E(n1983), .C(inClock), .Q(
        \u_inFIFO/FIFO[110][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[110][2]  ( .D(n1064), .E(n1983), .C(inClock), .Q(
        \u_inFIFO/FIFO[110][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[110][3]  ( .D(n1080), .E(n1983), .C(inClock), .Q(
        \u_inFIFO/FIFO[110][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[114][0]  ( .D(n1033), .E(n1979), .C(inClock), .Q(
        \u_inFIFO/FIFO[114][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[114][1]  ( .D(n1049), .E(n1979), .C(inClock), .Q(
        \u_inFIFO/FIFO[114][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[114][2]  ( .D(n1065), .E(n1979), .C(inClock), .Q(
        \u_inFIFO/FIFO[114][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[114][3]  ( .D(n1081), .E(n1979), .C(inClock), .Q(
        \u_inFIFO/FIFO[114][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[118][0]  ( .D(n1033), .E(n1975), .C(inClock), .Q(
        \u_inFIFO/FIFO[118][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[118][1]  ( .D(n1049), .E(n1975), .C(inClock), .Q(
        \u_inFIFO/FIFO[118][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[118][2]  ( .D(n1065), .E(n1975), .C(inClock), .Q(
        \u_inFIFO/FIFO[118][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[118][3]  ( .D(n1081), .E(n1975), .C(inClock), .Q(
        \u_inFIFO/FIFO[118][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[122][0]  ( .D(n1034), .E(n1971), .C(inClock), .Q(
        \u_inFIFO/FIFO[122][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[122][1]  ( .D(n1050), .E(n1971), .C(inClock), .Q(
        \u_inFIFO/FIFO[122][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[122][2]  ( .D(n1066), .E(n1971), .C(inClock), .Q(
        \u_inFIFO/FIFO[122][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[122][3]  ( .D(n1082), .E(n1971), .C(inClock), .Q(
        \u_inFIFO/FIFO[122][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[126][0]  ( .D(n1034), .E(n1967), .C(inClock), .Q(
        \u_inFIFO/FIFO[126][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[126][1]  ( .D(n1050), .E(n1967), .C(inClock), .Q(
        \u_inFIFO/FIFO[126][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[126][2]  ( .D(n1066), .E(n1967), .C(inClock), .Q(
        \u_inFIFO/FIFO[126][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[126][3]  ( .D(n1082), .E(n1967), .C(inClock), .Q(
        \u_inFIFO/FIFO[126][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[0][0]  ( .D(n1019), .E(n2093), .C(inClock), .Q(
        \u_inFIFO/FIFO[0][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[0][1]  ( .D(n1035), .E(n2093), .C(inClock), .Q(
        \u_inFIFO/FIFO[0][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[0][2]  ( .D(n1051), .E(n2093), .C(inClock), .Q(
        \u_inFIFO/FIFO[0][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[0][3]  ( .D(n1067), .E(n2093), .C(inClock), .Q(
        \u_inFIFO/FIFO[0][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[1][0]  ( .D(n1019), .E(n2092), .C(inClock), .Q(
        \u_inFIFO/FIFO[1][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[1][1]  ( .D(n1035), .E(n2092), .C(inClock), .Q(
        \u_inFIFO/FIFO[1][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[1][2]  ( .D(n1051), .E(n2092), .C(inClock), .Q(
        \u_inFIFO/FIFO[1][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[1][3]  ( .D(n1067), .E(n2092), .C(inClock), .Q(
        \u_inFIFO/FIFO[1][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[3][0]  ( .D(n1019), .E(n2090), .C(inClock), .Q(
        \u_inFIFO/FIFO[3][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[3][1]  ( .D(n1035), .E(n2090), .C(inClock), .Q(
        \u_inFIFO/FIFO[3][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[3][2]  ( .D(n1051), .E(n2090), .C(inClock), .Q(
        \u_inFIFO/FIFO[3][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[3][3]  ( .D(n1067), .E(n2090), .C(inClock), .Q(
        \u_inFIFO/FIFO[3][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[4][0]  ( .D(n1019), .E(n2089), .C(inClock), .Q(
        \u_inFIFO/FIFO[4][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[4][1]  ( .D(n1035), .E(n2089), .C(inClock), .Q(
        \u_inFIFO/FIFO[4][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[4][2]  ( .D(n1051), .E(n2089), .C(inClock), .Q(
        \u_inFIFO/FIFO[4][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[4][3]  ( .D(n1067), .E(n2089), .C(inClock), .Q(
        \u_inFIFO/FIFO[4][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[5][0]  ( .D(n1019), .E(n2088), .C(inClock), .Q(
        \u_inFIFO/FIFO[5][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[5][1]  ( .D(n1035), .E(n2088), .C(inClock), .Q(
        \u_inFIFO/FIFO[5][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[5][2]  ( .D(n1051), .E(n2088), .C(inClock), .Q(
        \u_inFIFO/FIFO[5][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[5][3]  ( .D(n1067), .E(n2088), .C(inClock), .Q(
        \u_inFIFO/FIFO[5][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[7][0]  ( .D(n1019), .E(n2086), .C(inClock), .Q(
        \u_inFIFO/FIFO[7][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[7][1]  ( .D(n1035), .E(n2086), .C(inClock), .Q(
        \u_inFIFO/FIFO[7][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[7][2]  ( .D(n1051), .E(n2086), .C(inClock), .Q(
        \u_inFIFO/FIFO[7][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[7][3]  ( .D(n1067), .E(n2086), .C(inClock), .Q(
        \u_inFIFO/FIFO[7][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[8][0]  ( .D(n1020), .E(n2085), .C(inClock), .Q(
        \u_inFIFO/FIFO[8][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[8][1]  ( .D(n1036), .E(n2085), .C(inClock), .Q(
        \u_inFIFO/FIFO[8][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[8][2]  ( .D(n1052), .E(n2085), .C(inClock), .Q(
        \u_inFIFO/FIFO[8][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[8][3]  ( .D(n1068), .E(n2085), .C(inClock), .Q(
        \u_inFIFO/FIFO[8][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[9][0]  ( .D(n1020), .E(n2084), .C(inClock), .Q(
        \u_inFIFO/FIFO[9][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[9][1]  ( .D(n1036), .E(n2084), .C(inClock), .Q(
        \u_inFIFO/FIFO[9][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[9][2]  ( .D(n1052), .E(n2084), .C(inClock), .Q(
        \u_inFIFO/FIFO[9][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[9][3]  ( .D(n1068), .E(n2084), .C(inClock), .Q(
        \u_inFIFO/FIFO[9][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[11][0]  ( .D(n1020), .E(n2082), .C(inClock), .Q(
        \u_inFIFO/FIFO[11][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[11][1]  ( .D(n1036), .E(n2082), .C(inClock), .Q(
        \u_inFIFO/FIFO[11][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[11][2]  ( .D(n1052), .E(n2082), .C(inClock), .Q(
        \u_inFIFO/FIFO[11][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[11][3]  ( .D(n1068), .E(n2082), .C(inClock), .Q(
        \u_inFIFO/FIFO[11][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[12][0]  ( .D(n1020), .E(n2081), .C(inClock), .Q(
        \u_inFIFO/FIFO[12][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[12][1]  ( .D(n1036), .E(n2081), .C(inClock), .Q(
        \u_inFIFO/FIFO[12][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[12][2]  ( .D(n1052), .E(n2081), .C(inClock), .Q(
        \u_inFIFO/FIFO[12][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[12][3]  ( .D(n1068), .E(n2081), .C(inClock), .Q(
        \u_inFIFO/FIFO[12][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[13][0]  ( .D(n1020), .E(n2080), .C(inClock), .Q(
        \u_inFIFO/FIFO[13][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[13][1]  ( .D(n1036), .E(n2080), .C(inClock), .Q(
        \u_inFIFO/FIFO[13][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[13][2]  ( .D(n1052), .E(n2080), .C(inClock), .Q(
        \u_inFIFO/FIFO[13][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[13][3]  ( .D(n1068), .E(n2080), .C(inClock), .Q(
        \u_inFIFO/FIFO[13][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[15][0]  ( .D(n1020), .E(n2078), .C(inClock), .Q(
        \u_inFIFO/FIFO[15][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[15][1]  ( .D(n1036), .E(n2078), .C(inClock), .Q(
        \u_inFIFO/FIFO[15][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[15][2]  ( .D(n1052), .E(n2078), .C(inClock), .Q(
        \u_inFIFO/FIFO[15][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[15][3]  ( .D(n1068), .E(n2078), .C(inClock), .Q(
        \u_inFIFO/FIFO[15][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[16][0]  ( .D(n1021), .E(n2077), .C(inClock), .Q(
        \u_inFIFO/FIFO[16][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[16][1]  ( .D(n1037), .E(n2077), .C(inClock), .Q(
        \u_inFIFO/FIFO[16][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[16][2]  ( .D(n1053), .E(n2077), .C(inClock), .Q(
        \u_inFIFO/FIFO[16][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[16][3]  ( .D(n1069), .E(n2077), .C(inClock), .Q(
        \u_inFIFO/FIFO[16][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[17][0]  ( .D(n1021), .E(n2076), .C(inClock), .Q(
        \u_inFIFO/FIFO[17][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[17][1]  ( .D(n1037), .E(n2076), .C(inClock), .Q(
        \u_inFIFO/FIFO[17][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[17][2]  ( .D(n1053), .E(n2076), .C(inClock), .Q(
        \u_inFIFO/FIFO[17][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[17][3]  ( .D(n1069), .E(n2076), .C(inClock), .Q(
        \u_inFIFO/FIFO[17][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[19][0]  ( .D(n1021), .E(n2074), .C(inClock), .Q(
        \u_inFIFO/FIFO[19][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[19][1]  ( .D(n1037), .E(n2074), .C(inClock), .Q(
        \u_inFIFO/FIFO[19][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[19][2]  ( .D(n1053), .E(n2074), .C(inClock), .Q(
        \u_inFIFO/FIFO[19][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[19][3]  ( .D(n1069), .E(n2074), .C(inClock), .Q(
        \u_inFIFO/FIFO[19][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[20][0]  ( .D(n1021), .E(n2073), .C(inClock), .Q(
        \u_inFIFO/FIFO[20][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[20][1]  ( .D(n1037), .E(n2073), .C(inClock), .Q(
        \u_inFIFO/FIFO[20][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[20][2]  ( .D(n1053), .E(n2073), .C(inClock), .Q(
        \u_inFIFO/FIFO[20][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[20][3]  ( .D(n1069), .E(n2073), .C(inClock), .Q(
        \u_inFIFO/FIFO[20][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[21][0]  ( .D(n1021), .E(n2072), .C(inClock), .Q(
        \u_inFIFO/FIFO[21][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[21][1]  ( .D(n1037), .E(n2072), .C(inClock), .Q(
        \u_inFIFO/FIFO[21][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[21][2]  ( .D(n1053), .E(n2072), .C(inClock), .Q(
        \u_inFIFO/FIFO[21][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[21][3]  ( .D(n1069), .E(n2072), .C(inClock), .Q(
        \u_inFIFO/FIFO[21][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[23][0]  ( .D(n1021), .E(n2070), .C(inClock), .Q(
        \u_inFIFO/FIFO[23][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[23][1]  ( .D(n1037), .E(n2070), .C(inClock), .Q(
        \u_inFIFO/FIFO[23][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[23][2]  ( .D(n1053), .E(n2070), .C(inClock), .Q(
        \u_inFIFO/FIFO[23][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[23][3]  ( .D(n1069), .E(n2070), .C(inClock), .Q(
        \u_inFIFO/FIFO[23][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[24][0]  ( .D(n1022), .E(n2069), .C(inClock), .Q(
        \u_inFIFO/FIFO[24][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[24][1]  ( .D(n1038), .E(n2069), .C(inClock), .Q(
        \u_inFIFO/FIFO[24][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[24][2]  ( .D(n1054), .E(n2069), .C(inClock), .Q(
        \u_inFIFO/FIFO[24][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[24][3]  ( .D(n1070), .E(n2069), .C(inClock), .Q(
        \u_inFIFO/FIFO[24][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[25][0]  ( .D(n1022), .E(n2068), .C(inClock), .Q(
        \u_inFIFO/FIFO[25][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[25][1]  ( .D(n1038), .E(n2068), .C(inClock), .Q(
        \u_inFIFO/FIFO[25][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[25][2]  ( .D(n1054), .E(n2068), .C(inClock), .Q(
        \u_inFIFO/FIFO[25][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[25][3]  ( .D(n1070), .E(n2068), .C(inClock), .Q(
        \u_inFIFO/FIFO[25][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[27][0]  ( .D(n1022), .E(n2066), .C(inClock), .Q(
        \u_inFIFO/FIFO[27][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[27][1]  ( .D(n1038), .E(n2066), .C(inClock), .Q(
        \u_inFIFO/FIFO[27][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[27][2]  ( .D(n1054), .E(n2066), .C(inClock), .Q(
        \u_inFIFO/FIFO[27][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[27][3]  ( .D(n1070), .E(n2066), .C(inClock), .Q(
        \u_inFIFO/FIFO[27][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[28][0]  ( .D(n1022), .E(n2065), .C(inClock), .Q(
        \u_inFIFO/FIFO[28][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[28][1]  ( .D(n1038), .E(n2065), .C(inClock), .Q(
        \u_inFIFO/FIFO[28][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[28][2]  ( .D(n1054), .E(n2065), .C(inClock), .Q(
        \u_inFIFO/FIFO[28][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[28][3]  ( .D(n1070), .E(n2065), .C(inClock), .Q(
        \u_inFIFO/FIFO[28][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[29][0]  ( .D(n1022), .E(n2064), .C(inClock), .Q(
        \u_inFIFO/FIFO[29][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[29][1]  ( .D(n1038), .E(n2064), .C(inClock), .Q(
        \u_inFIFO/FIFO[29][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[29][2]  ( .D(n1054), .E(n2064), .C(inClock), .Q(
        \u_inFIFO/FIFO[29][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[29][3]  ( .D(n1070), .E(n2064), .C(inClock), .Q(
        \u_inFIFO/FIFO[29][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[31][0]  ( .D(n1022), .E(n2062), .C(inClock), .Q(
        \u_inFIFO/FIFO[31][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[31][1]  ( .D(n1038), .E(n2062), .C(inClock), .Q(
        \u_inFIFO/FIFO[31][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[31][2]  ( .D(n1054), .E(n2062), .C(inClock), .Q(
        \u_inFIFO/FIFO[31][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[31][3]  ( .D(n1070), .E(n2062), .C(inClock), .Q(
        \u_inFIFO/FIFO[31][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[32][0]  ( .D(n1023), .E(n2061), .C(inClock), .Q(
        \u_inFIFO/FIFO[32][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[32][1]  ( .D(n1039), .E(n2061), .C(inClock), .Q(
        \u_inFIFO/FIFO[32][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[32][2]  ( .D(n1055), .E(n2061), .C(inClock), .Q(
        \u_inFIFO/FIFO[32][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[32][3]  ( .D(n1071), .E(n2061), .C(inClock), .Q(
        \u_inFIFO/FIFO[32][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[33][0]  ( .D(n1023), .E(n2060), .C(inClock), .Q(
        \u_inFIFO/FIFO[33][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[33][1]  ( .D(n1039), .E(n2060), .C(inClock), .Q(
        \u_inFIFO/FIFO[33][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[33][2]  ( .D(n1055), .E(n2060), .C(inClock), .Q(
        \u_inFIFO/FIFO[33][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[33][3]  ( .D(n1071), .E(n2060), .C(inClock), .Q(
        \u_inFIFO/FIFO[33][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[35][0]  ( .D(n1023), .E(n2058), .C(inClock), .Q(
        \u_inFIFO/FIFO[35][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[35][1]  ( .D(n1039), .E(n2058), .C(inClock), .Q(
        \u_inFIFO/FIFO[35][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[35][2]  ( .D(n1055), .E(n2058), .C(inClock), .Q(
        \u_inFIFO/FIFO[35][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[35][3]  ( .D(n1071), .E(n2058), .C(inClock), .Q(
        \u_inFIFO/FIFO[35][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[36][0]  ( .D(n1023), .E(n2057), .C(inClock), .Q(
        \u_inFIFO/FIFO[36][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[36][1]  ( .D(n1039), .E(n2057), .C(inClock), .Q(
        \u_inFIFO/FIFO[36][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[36][2]  ( .D(n1055), .E(n2057), .C(inClock), .Q(
        \u_inFIFO/FIFO[36][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[36][3]  ( .D(n1071), .E(n2057), .C(inClock), .Q(
        \u_inFIFO/FIFO[36][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[37][0]  ( .D(n1023), .E(n2056), .C(inClock), .Q(
        \u_inFIFO/FIFO[37][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[37][1]  ( .D(n1039), .E(n2056), .C(inClock), .Q(
        \u_inFIFO/FIFO[37][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[37][2]  ( .D(n1055), .E(n2056), .C(inClock), .Q(
        \u_inFIFO/FIFO[37][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[37][3]  ( .D(n1071), .E(n2056), .C(inClock), .Q(
        \u_inFIFO/FIFO[37][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[39][0]  ( .D(n1023), .E(n2054), .C(inClock), .Q(
        \u_inFIFO/FIFO[39][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[39][1]  ( .D(n1039), .E(n2054), .C(inClock), .Q(
        \u_inFIFO/FIFO[39][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[39][2]  ( .D(n1055), .E(n2054), .C(inClock), .Q(
        \u_inFIFO/FIFO[39][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[39][3]  ( .D(n1071), .E(n2054), .C(inClock), .Q(
        \u_inFIFO/FIFO[39][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[40][0]  ( .D(n1024), .E(n2053), .C(inClock), .Q(
        \u_inFIFO/FIFO[40][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[40][1]  ( .D(n1040), .E(n2053), .C(inClock), .Q(
        \u_inFIFO/FIFO[40][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[40][2]  ( .D(n1056), .E(n2053), .C(inClock), .Q(
        \u_inFIFO/FIFO[40][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[40][3]  ( .D(n1072), .E(n2053), .C(inClock), .Q(
        \u_inFIFO/FIFO[40][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[41][0]  ( .D(n1024), .E(n2052), .C(inClock), .Q(
        \u_inFIFO/FIFO[41][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[41][1]  ( .D(n1040), .E(n2052), .C(inClock), .Q(
        \u_inFIFO/FIFO[41][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[41][2]  ( .D(n1056), .E(n2052), .C(inClock), .Q(
        \u_inFIFO/FIFO[41][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[41][3]  ( .D(n1072), .E(n2052), .C(inClock), .Q(
        \u_inFIFO/FIFO[41][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[43][0]  ( .D(n1024), .E(n2050), .C(inClock), .Q(
        \u_inFIFO/FIFO[43][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[43][1]  ( .D(n1040), .E(n2050), .C(inClock), .Q(
        \u_inFIFO/FIFO[43][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[43][2]  ( .D(n1056), .E(n2050), .C(inClock), .Q(
        \u_inFIFO/FIFO[43][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[43][3]  ( .D(n1072), .E(n2050), .C(inClock), .Q(
        \u_inFIFO/FIFO[43][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[44][0]  ( .D(n1024), .E(n2049), .C(inClock), .Q(
        \u_inFIFO/FIFO[44][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[44][1]  ( .D(n1040), .E(n2049), .C(inClock), .Q(
        \u_inFIFO/FIFO[44][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[44][2]  ( .D(n1056), .E(n2049), .C(inClock), .Q(
        \u_inFIFO/FIFO[44][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[44][3]  ( .D(n1072), .E(n2049), .C(inClock), .Q(
        \u_inFIFO/FIFO[44][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[45][0]  ( .D(n1024), .E(n2048), .C(inClock), .Q(
        \u_inFIFO/FIFO[45][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[45][1]  ( .D(n1040), .E(n2048), .C(inClock), .Q(
        \u_inFIFO/FIFO[45][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[45][2]  ( .D(n1056), .E(n2048), .C(inClock), .Q(
        \u_inFIFO/FIFO[45][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[45][3]  ( .D(n1072), .E(n2048), .C(inClock), .Q(
        \u_inFIFO/FIFO[45][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[47][0]  ( .D(n1024), .E(n2046), .C(inClock), .Q(
        \u_inFIFO/FIFO[47][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[47][1]  ( .D(n1040), .E(n2046), .C(inClock), .Q(
        \u_inFIFO/FIFO[47][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[47][2]  ( .D(n1056), .E(n2046), .C(inClock), .Q(
        \u_inFIFO/FIFO[47][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[47][3]  ( .D(n1072), .E(n2046), .C(inClock), .Q(
        \u_inFIFO/FIFO[47][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[48][0]  ( .D(n1025), .E(n2045), .C(inClock), .Q(
        \u_inFIFO/FIFO[48][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[48][1]  ( .D(n1041), .E(n2045), .C(inClock), .Q(
        \u_inFIFO/FIFO[48][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[48][2]  ( .D(n1057), .E(n2045), .C(inClock), .Q(
        \u_inFIFO/FIFO[48][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[48][3]  ( .D(n1073), .E(n2045), .C(inClock), .Q(
        \u_inFIFO/FIFO[48][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[49][0]  ( .D(n1025), .E(n2044), .C(inClock), .Q(
        \u_inFIFO/FIFO[49][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[49][1]  ( .D(n1041), .E(n2044), .C(inClock), .Q(
        \u_inFIFO/FIFO[49][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[49][2]  ( .D(n1057), .E(n2044), .C(inClock), .Q(
        \u_inFIFO/FIFO[49][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[49][3]  ( .D(n1073), .E(n2044), .C(inClock), .Q(
        \u_inFIFO/FIFO[49][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[51][0]  ( .D(n1025), .E(n2042), .C(inClock), .Q(
        \u_inFIFO/FIFO[51][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[51][1]  ( .D(n1041), .E(n2042), .C(inClock), .Q(
        \u_inFIFO/FIFO[51][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[51][2]  ( .D(n1057), .E(n2042), .C(inClock), .Q(
        \u_inFIFO/FIFO[51][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[51][3]  ( .D(n1073), .E(n2042), .C(inClock), .Q(
        \u_inFIFO/FIFO[51][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[52][0]  ( .D(n1025), .E(n2041), .C(inClock), .Q(
        \u_inFIFO/FIFO[52][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[52][1]  ( .D(n1041), .E(n2041), .C(inClock), .Q(
        \u_inFIFO/FIFO[52][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[52][2]  ( .D(n1057), .E(n2041), .C(inClock), .Q(
        \u_inFIFO/FIFO[52][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[52][3]  ( .D(n1073), .E(n2041), .C(inClock), .Q(
        \u_inFIFO/FIFO[52][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[53][0]  ( .D(n1025), .E(n2040), .C(inClock), .Q(
        \u_inFIFO/FIFO[53][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[53][1]  ( .D(n1041), .E(n2040), .C(inClock), .Q(
        \u_inFIFO/FIFO[53][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[53][2]  ( .D(n1057), .E(n2040), .C(inClock), .Q(
        \u_inFIFO/FIFO[53][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[53][3]  ( .D(n1073), .E(n2040), .C(inClock), .Q(
        \u_inFIFO/FIFO[53][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[55][0]  ( .D(n1025), .E(n2038), .C(inClock), .Q(
        \u_inFIFO/FIFO[55][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[55][1]  ( .D(n1041), .E(n2038), .C(inClock), .Q(
        \u_inFIFO/FIFO[55][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[55][2]  ( .D(n1057), .E(n2038), .C(inClock), .Q(
        \u_inFIFO/FIFO[55][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[55][3]  ( .D(n1073), .E(n2038), .C(inClock), .Q(
        \u_inFIFO/FIFO[55][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[56][0]  ( .D(n1026), .E(n2037), .C(inClock), .Q(
        \u_inFIFO/FIFO[56][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[56][1]  ( .D(n1042), .E(n2037), .C(inClock), .Q(
        \u_inFIFO/FIFO[56][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[56][2]  ( .D(n1058), .E(n2037), .C(inClock), .Q(
        \u_inFIFO/FIFO[56][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[56][3]  ( .D(n1074), .E(n2037), .C(inClock), .Q(
        \u_inFIFO/FIFO[56][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[57][0]  ( .D(n1026), .E(n2036), .C(inClock), .Q(
        \u_inFIFO/FIFO[57][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[57][1]  ( .D(n1042), .E(n2036), .C(inClock), .Q(
        \u_inFIFO/FIFO[57][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[57][2]  ( .D(n1058), .E(n2036), .C(inClock), .Q(
        \u_inFIFO/FIFO[57][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[57][3]  ( .D(n1074), .E(n2036), .C(inClock), .Q(
        \u_inFIFO/FIFO[57][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[59][0]  ( .D(n1026), .E(n2034), .C(inClock), .Q(
        \u_inFIFO/FIFO[59][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[59][1]  ( .D(n1042), .E(n2034), .C(inClock), .Q(
        \u_inFIFO/FIFO[59][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[59][2]  ( .D(n1058), .E(n2034), .C(inClock), .Q(
        \u_inFIFO/FIFO[59][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[59][3]  ( .D(n1074), .E(n2034), .C(inClock), .Q(
        \u_inFIFO/FIFO[59][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[60][0]  ( .D(n1026), .E(n2033), .C(inClock), .Q(
        \u_inFIFO/FIFO[60][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[60][1]  ( .D(n1042), .E(n2033), .C(inClock), .Q(
        \u_inFIFO/FIFO[60][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[60][2]  ( .D(n1058), .E(n2033), .C(inClock), .Q(
        \u_inFIFO/FIFO[60][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[60][3]  ( .D(n1074), .E(n2033), .C(inClock), .Q(
        \u_inFIFO/FIFO[60][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[61][0]  ( .D(n1026), .E(n2032), .C(inClock), .Q(
        \u_inFIFO/FIFO[61][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[61][1]  ( .D(n1042), .E(n2032), .C(inClock), .Q(
        \u_inFIFO/FIFO[61][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[61][2]  ( .D(n1058), .E(n2032), .C(inClock), .Q(
        \u_inFIFO/FIFO[61][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[61][3]  ( .D(n1074), .E(n2032), .C(inClock), .Q(
        \u_inFIFO/FIFO[61][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[63][0]  ( .D(n1026), .E(n2030), .C(inClock), .Q(
        \u_inFIFO/FIFO[63][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[63][1]  ( .D(n1042), .E(n2030), .C(inClock), .Q(
        \u_inFIFO/FIFO[63][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[63][2]  ( .D(n1058), .E(n2030), .C(inClock), .Q(
        \u_inFIFO/FIFO[63][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[63][3]  ( .D(n1074), .E(n2030), .C(inClock), .Q(
        \u_inFIFO/FIFO[63][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[64][0]  ( .D(n1027), .E(n2029), .C(inClock), .Q(
        \u_inFIFO/FIFO[64][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[64][1]  ( .D(n1043), .E(n2029), .C(inClock), .Q(
        \u_inFIFO/FIFO[64][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[64][2]  ( .D(n1059), .E(n2029), .C(inClock), .Q(
        \u_inFIFO/FIFO[64][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[64][3]  ( .D(n1075), .E(n2029), .C(inClock), .Q(
        \u_inFIFO/FIFO[64][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[65][0]  ( .D(n1027), .E(n2028), .C(inClock), .Q(
        \u_inFIFO/FIFO[65][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[65][1]  ( .D(n1043), .E(n2028), .C(inClock), .Q(
        \u_inFIFO/FIFO[65][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[65][2]  ( .D(n1059), .E(n2028), .C(inClock), .Q(
        \u_inFIFO/FIFO[65][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[65][3]  ( .D(n1075), .E(n2028), .C(inClock), .Q(
        \u_inFIFO/FIFO[65][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[67][0]  ( .D(n1027), .E(n2026), .C(inClock), .Q(
        \u_inFIFO/FIFO[67][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[67][1]  ( .D(n1043), .E(n2026), .C(inClock), .Q(
        \u_inFIFO/FIFO[67][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[67][2]  ( .D(n1059), .E(n2026), .C(inClock), .Q(
        \u_inFIFO/FIFO[67][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[67][3]  ( .D(n1075), .E(n2026), .C(inClock), .Q(
        \u_inFIFO/FIFO[67][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[68][0]  ( .D(n1027), .E(n2025), .C(inClock), .Q(
        \u_inFIFO/FIFO[68][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[68][1]  ( .D(n1043), .E(n2025), .C(inClock), .Q(
        \u_inFIFO/FIFO[68][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[68][2]  ( .D(n1059), .E(n2025), .C(inClock), .Q(
        \u_inFIFO/FIFO[68][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[68][3]  ( .D(n1075), .E(n2025), .C(inClock), .Q(
        \u_inFIFO/FIFO[68][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[69][0]  ( .D(n1027), .E(n2024), .C(inClock), .Q(
        \u_inFIFO/FIFO[69][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[69][1]  ( .D(n1043), .E(n2024), .C(inClock), .Q(
        \u_inFIFO/FIFO[69][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[69][2]  ( .D(n1059), .E(n2024), .C(inClock), .Q(
        \u_inFIFO/FIFO[69][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[69][3]  ( .D(n1075), .E(n2024), .C(inClock), .Q(
        \u_inFIFO/FIFO[69][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[71][0]  ( .D(n1027), .E(n2022), .C(inClock), .Q(
        \u_inFIFO/FIFO[71][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[71][1]  ( .D(n1043), .E(n2022), .C(inClock), .Q(
        \u_inFIFO/FIFO[71][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[71][2]  ( .D(n1059), .E(n2022), .C(inClock), .Q(
        \u_inFIFO/FIFO[71][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[71][3]  ( .D(n1075), .E(n2022), .C(inClock), .Q(
        \u_inFIFO/FIFO[71][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[72][0]  ( .D(n1028), .E(n2021), .C(inClock), .Q(
        \u_inFIFO/FIFO[72][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[72][1]  ( .D(n1044), .E(n2021), .C(inClock), .Q(
        \u_inFIFO/FIFO[72][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[72][2]  ( .D(n1060), .E(n2021), .C(inClock), .Q(
        \u_inFIFO/FIFO[72][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[72][3]  ( .D(n1076), .E(n2021), .C(inClock), .Q(
        \u_inFIFO/FIFO[72][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[73][0]  ( .D(n1028), .E(n2020), .C(inClock), .Q(
        \u_inFIFO/FIFO[73][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[73][1]  ( .D(n1044), .E(n2020), .C(inClock), .Q(
        \u_inFIFO/FIFO[73][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[73][2]  ( .D(n1060), .E(n2020), .C(inClock), .Q(
        \u_inFIFO/FIFO[73][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[73][3]  ( .D(n1076), .E(n2020), .C(inClock), .Q(
        \u_inFIFO/FIFO[73][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[75][0]  ( .D(n1028), .E(n2018), .C(inClock), .Q(
        \u_inFIFO/FIFO[75][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[75][1]  ( .D(n1044), .E(n2018), .C(inClock), .Q(
        \u_inFIFO/FIFO[75][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[75][2]  ( .D(n1060), .E(n2018), .C(inClock), .Q(
        \u_inFIFO/FIFO[75][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[75][3]  ( .D(n1076), .E(n2018), .C(inClock), .Q(
        \u_inFIFO/FIFO[75][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[76][0]  ( .D(n1028), .E(n2017), .C(inClock), .Q(
        \u_inFIFO/FIFO[76][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[76][1]  ( .D(n1044), .E(n2017), .C(inClock), .Q(
        \u_inFIFO/FIFO[76][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[76][2]  ( .D(n1060), .E(n2017), .C(inClock), .Q(
        \u_inFIFO/FIFO[76][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[76][3]  ( .D(n1076), .E(n2017), .C(inClock), .Q(
        \u_inFIFO/FIFO[76][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[77][0]  ( .D(n1028), .E(n2016), .C(inClock), .Q(
        \u_inFIFO/FIFO[77][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[77][1]  ( .D(n1044), .E(n2016), .C(inClock), .Q(
        \u_inFIFO/FIFO[77][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[77][2]  ( .D(n1060), .E(n2016), .C(inClock), .Q(
        \u_inFIFO/FIFO[77][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[77][3]  ( .D(n1076), .E(n2016), .C(inClock), .Q(
        \u_inFIFO/FIFO[77][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[79][0]  ( .D(n1028), .E(n2014), .C(inClock), .Q(
        \u_inFIFO/FIFO[79][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[79][1]  ( .D(n1044), .E(n2014), .C(inClock), .Q(
        \u_inFIFO/FIFO[79][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[79][2]  ( .D(n1060), .E(n2014), .C(inClock), .Q(
        \u_inFIFO/FIFO[79][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[79][3]  ( .D(n1076), .E(n2014), .C(inClock), .Q(
        \u_inFIFO/FIFO[79][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[80][0]  ( .D(n1029), .E(n2013), .C(inClock), .Q(
        \u_inFIFO/FIFO[80][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[80][1]  ( .D(n1045), .E(n2013), .C(inClock), .Q(
        \u_inFIFO/FIFO[80][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[80][2]  ( .D(n1061), .E(n2013), .C(inClock), .Q(
        \u_inFIFO/FIFO[80][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[80][3]  ( .D(n1077), .E(n2013), .C(inClock), .Q(
        \u_inFIFO/FIFO[80][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[81][0]  ( .D(n1029), .E(n2012), .C(inClock), .Q(
        \u_inFIFO/FIFO[81][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[81][1]  ( .D(n1045), .E(n2012), .C(inClock), .Q(
        \u_inFIFO/FIFO[81][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[81][2]  ( .D(n1061), .E(n2012), .C(inClock), .Q(
        \u_inFIFO/FIFO[81][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[81][3]  ( .D(n1077), .E(n2012), .C(inClock), .Q(
        \u_inFIFO/FIFO[81][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[83][0]  ( .D(n1029), .E(n2010), .C(inClock), .Q(
        \u_inFIFO/FIFO[83][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[83][1]  ( .D(n1045), .E(n2010), .C(inClock), .Q(
        \u_inFIFO/FIFO[83][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[83][2]  ( .D(n1061), .E(n2010), .C(inClock), .Q(
        \u_inFIFO/FIFO[83][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[83][3]  ( .D(n1077), .E(n2010), .C(inClock), .Q(
        \u_inFIFO/FIFO[83][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[84][0]  ( .D(n1029), .E(n2009), .C(inClock), .Q(
        \u_inFIFO/FIFO[84][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[84][1]  ( .D(n1045), .E(n2009), .C(inClock), .Q(
        \u_inFIFO/FIFO[84][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[84][2]  ( .D(n1061), .E(n2009), .C(inClock), .Q(
        \u_inFIFO/FIFO[84][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[84][3]  ( .D(n1077), .E(n2009), .C(inClock), .Q(
        \u_inFIFO/FIFO[84][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[85][0]  ( .D(n1029), .E(n2008), .C(inClock), .Q(
        \u_inFIFO/FIFO[85][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[85][1]  ( .D(n1045), .E(n2008), .C(inClock), .Q(
        \u_inFIFO/FIFO[85][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[85][2]  ( .D(n1061), .E(n2008), .C(inClock), .Q(
        \u_inFIFO/FIFO[85][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[85][3]  ( .D(n1077), .E(n2008), .C(inClock), .Q(
        \u_inFIFO/FIFO[85][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[87][0]  ( .D(n1029), .E(n2006), .C(inClock), .Q(
        \u_inFIFO/FIFO[87][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[87][1]  ( .D(n1045), .E(n2006), .C(inClock), .Q(
        \u_inFIFO/FIFO[87][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[87][2]  ( .D(n1061), .E(n2006), .C(inClock), .Q(
        \u_inFIFO/FIFO[87][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[87][3]  ( .D(n1077), .E(n2006), .C(inClock), .Q(
        \u_inFIFO/FIFO[87][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[88][0]  ( .D(n1030), .E(n2005), .C(inClock), .Q(
        \u_inFIFO/FIFO[88][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[88][1]  ( .D(n1046), .E(n2005), .C(inClock), .Q(
        \u_inFIFO/FIFO[88][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[88][2]  ( .D(n1062), .E(n2005), .C(inClock), .Q(
        \u_inFIFO/FIFO[88][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[88][3]  ( .D(n1078), .E(n2005), .C(inClock), .Q(
        \u_inFIFO/FIFO[88][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[89][0]  ( .D(n1030), .E(n2004), .C(inClock), .Q(
        \u_inFIFO/FIFO[89][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[89][1]  ( .D(n1046), .E(n2004), .C(inClock), .Q(
        \u_inFIFO/FIFO[89][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[89][2]  ( .D(n1062), .E(n2004), .C(inClock), .Q(
        \u_inFIFO/FIFO[89][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[89][3]  ( .D(n1078), .E(n2004), .C(inClock), .Q(
        \u_inFIFO/FIFO[89][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[91][0]  ( .D(n1030), .E(n2002), .C(inClock), .Q(
        \u_inFIFO/FIFO[91][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[91][1]  ( .D(n1046), .E(n2002), .C(inClock), .Q(
        \u_inFIFO/FIFO[91][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[91][2]  ( .D(n1062), .E(n2002), .C(inClock), .Q(
        \u_inFIFO/FIFO[91][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[91][3]  ( .D(n1078), .E(n2002), .C(inClock), .Q(
        \u_inFIFO/FIFO[91][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[92][0]  ( .D(n1030), .E(n2001), .C(inClock), .Q(
        \u_inFIFO/FIFO[92][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[92][1]  ( .D(n1046), .E(n2001), .C(inClock), .Q(
        \u_inFIFO/FIFO[92][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[92][2]  ( .D(n1062), .E(n2001), .C(inClock), .Q(
        \u_inFIFO/FIFO[92][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[92][3]  ( .D(n1078), .E(n2001), .C(inClock), .Q(
        \u_inFIFO/FIFO[92][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[93][0]  ( .D(n1030), .E(n2000), .C(inClock), .Q(
        \u_inFIFO/FIFO[93][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[93][1]  ( .D(n1046), .E(n2000), .C(inClock), .Q(
        \u_inFIFO/FIFO[93][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[93][2]  ( .D(n1062), .E(n2000), .C(inClock), .Q(
        \u_inFIFO/FIFO[93][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[93][3]  ( .D(n1078), .E(n2000), .C(inClock), .Q(
        \u_inFIFO/FIFO[93][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[95][0]  ( .D(n1030), .E(n1998), .C(inClock), .Q(
        \u_inFIFO/FIFO[95][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[95][1]  ( .D(n1046), .E(n1998), .C(inClock), .Q(
        \u_inFIFO/FIFO[95][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[95][2]  ( .D(n1062), .E(n1998), .C(inClock), .Q(
        \u_inFIFO/FIFO[95][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[95][3]  ( .D(n1078), .E(n1998), .C(inClock), .Q(
        \u_inFIFO/FIFO[95][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[96][0]  ( .D(n1031), .E(n1997), .C(inClock), .Q(
        \u_inFIFO/FIFO[96][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[96][1]  ( .D(n1047), .E(n1997), .C(inClock), .Q(
        \u_inFIFO/FIFO[96][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[96][2]  ( .D(n1063), .E(n1997), .C(inClock), .Q(
        \u_inFIFO/FIFO[96][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[96][3]  ( .D(n1079), .E(n1997), .C(inClock), .Q(
        \u_inFIFO/FIFO[96][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[97][0]  ( .D(n1031), .E(n1996), .C(inClock), .Q(
        \u_inFIFO/FIFO[97][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[97][1]  ( .D(n1047), .E(n1996), .C(inClock), .Q(
        \u_inFIFO/FIFO[97][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[97][2]  ( .D(n1063), .E(n1996), .C(inClock), .Q(
        \u_inFIFO/FIFO[97][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[97][3]  ( .D(n1079), .E(n1996), .C(inClock), .Q(
        \u_inFIFO/FIFO[97][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[99][0]  ( .D(n1031), .E(n1994), .C(inClock), .Q(
        \u_inFIFO/FIFO[99][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[99][1]  ( .D(n1047), .E(n1994), .C(inClock), .Q(
        \u_inFIFO/FIFO[99][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[99][2]  ( .D(n1063), .E(n1994), .C(inClock), .Q(
        \u_inFIFO/FIFO[99][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[99][3]  ( .D(n1079), .E(n1994), .C(inClock), .Q(
        \u_inFIFO/FIFO[99][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[100][0]  ( .D(n1031), .E(n1993), .C(inClock), .Q(
        \u_inFIFO/FIFO[100][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[100][1]  ( .D(n1047), .E(n1993), .C(inClock), .Q(
        \u_inFIFO/FIFO[100][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[100][2]  ( .D(n1063), .E(n1993), .C(inClock), .Q(
        \u_inFIFO/FIFO[100][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[100][3]  ( .D(n1079), .E(n1993), .C(inClock), .Q(
        \u_inFIFO/FIFO[100][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[101][0]  ( .D(n1031), .E(n1992), .C(inClock), .Q(
        \u_inFIFO/FIFO[101][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[101][1]  ( .D(n1047), .E(n1992), .C(inClock), .Q(
        \u_inFIFO/FIFO[101][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[101][2]  ( .D(n1063), .E(n1992), .C(inClock), .Q(
        \u_inFIFO/FIFO[101][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[101][3]  ( .D(n1079), .E(n1992), .C(inClock), .Q(
        \u_inFIFO/FIFO[101][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[103][0]  ( .D(n1031), .E(n1990), .C(inClock), .Q(
        \u_inFIFO/FIFO[103][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[103][1]  ( .D(n1047), .E(n1990), .C(inClock), .Q(
        \u_inFIFO/FIFO[103][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[103][2]  ( .D(n1063), .E(n1990), .C(inClock), .Q(
        \u_inFIFO/FIFO[103][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[103][3]  ( .D(n1079), .E(n1990), .C(inClock), .Q(
        \u_inFIFO/FIFO[103][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[104][0]  ( .D(n1032), .E(n1989), .C(inClock), .Q(
        \u_inFIFO/FIFO[104][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[104][1]  ( .D(n1048), .E(n1989), .C(inClock), .Q(
        \u_inFIFO/FIFO[104][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[104][2]  ( .D(n1064), .E(n1989), .C(inClock), .Q(
        \u_inFIFO/FIFO[104][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[104][3]  ( .D(n1080), .E(n1989), .C(inClock), .Q(
        \u_inFIFO/FIFO[104][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[105][0]  ( .D(n1032), .E(n1988), .C(inClock), .Q(
        \u_inFIFO/FIFO[105][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[105][1]  ( .D(n1048), .E(n1988), .C(inClock), .Q(
        \u_inFIFO/FIFO[105][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[105][2]  ( .D(n1064), .E(n1988), .C(inClock), .Q(
        \u_inFIFO/FIFO[105][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[105][3]  ( .D(n1080), .E(n1988), .C(inClock), .Q(
        \u_inFIFO/FIFO[105][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[107][0]  ( .D(n1032), .E(n1986), .C(inClock), .Q(
        \u_inFIFO/FIFO[107][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[107][1]  ( .D(n1048), .E(n1986), .C(inClock), .Q(
        \u_inFIFO/FIFO[107][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[107][2]  ( .D(n1064), .E(n1986), .C(inClock), .Q(
        \u_inFIFO/FIFO[107][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[107][3]  ( .D(n1080), .E(n1986), .C(inClock), .Q(
        \u_inFIFO/FIFO[107][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[108][0]  ( .D(n1032), .E(n1985), .C(inClock), .Q(
        \u_inFIFO/FIFO[108][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[108][1]  ( .D(n1048), .E(n1985), .C(inClock), .Q(
        \u_inFIFO/FIFO[108][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[108][2]  ( .D(n1064), .E(n1985), .C(inClock), .Q(
        \u_inFIFO/FIFO[108][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[108][3]  ( .D(n1080), .E(n1985), .C(inClock), .Q(
        \u_inFIFO/FIFO[108][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[109][0]  ( .D(n1032), .E(n1984), .C(inClock), .Q(
        \u_inFIFO/FIFO[109][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[109][1]  ( .D(n1048), .E(n1984), .C(inClock), .Q(
        \u_inFIFO/FIFO[109][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[109][2]  ( .D(n1064), .E(n1984), .C(inClock), .Q(
        \u_inFIFO/FIFO[109][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[109][3]  ( .D(n1080), .E(n1984), .C(inClock), .Q(
        \u_inFIFO/FIFO[109][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[111][0]  ( .D(n1032), .E(n1982), .C(inClock), .Q(
        \u_inFIFO/FIFO[111][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[111][1]  ( .D(n1048), .E(n1982), .C(inClock), .Q(
        \u_inFIFO/FIFO[111][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[111][2]  ( .D(n1064), .E(n1982), .C(inClock), .Q(
        \u_inFIFO/FIFO[111][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[111][3]  ( .D(n1080), .E(n1982), .C(inClock), .Q(
        \u_inFIFO/FIFO[111][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[112][0]  ( .D(n1033), .E(n1981), .C(inClock), .Q(
        \u_inFIFO/FIFO[112][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[112][1]  ( .D(n1049), .E(n1981), .C(inClock), .Q(
        \u_inFIFO/FIFO[112][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[112][2]  ( .D(n1065), .E(n1981), .C(inClock), .Q(
        \u_inFIFO/FIFO[112][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[112][3]  ( .D(n1081), .E(n1981), .C(inClock), .Q(
        \u_inFIFO/FIFO[112][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[113][0]  ( .D(n1033), .E(n1980), .C(inClock), .Q(
        \u_inFIFO/FIFO[113][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[113][1]  ( .D(n1049), .E(n1980), .C(inClock), .Q(
        \u_inFIFO/FIFO[113][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[113][2]  ( .D(n1065), .E(n1980), .C(inClock), .Q(
        \u_inFIFO/FIFO[113][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[113][3]  ( .D(n1081), .E(n1980), .C(inClock), .Q(
        \u_inFIFO/FIFO[113][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[115][0]  ( .D(n1033), .E(n1978), .C(inClock), .Q(
        \u_inFIFO/FIFO[115][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[115][1]  ( .D(n1049), .E(n1978), .C(inClock), .Q(
        \u_inFIFO/FIFO[115][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[115][2]  ( .D(n1065), .E(n1978), .C(inClock), .Q(
        \u_inFIFO/FIFO[115][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[115][3]  ( .D(n1081), .E(n1978), .C(inClock), .Q(
        \u_inFIFO/FIFO[115][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[116][0]  ( .D(n1033), .E(n1977), .C(inClock), .Q(
        \u_inFIFO/FIFO[116][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[116][1]  ( .D(n1049), .E(n1977), .C(inClock), .Q(
        \u_inFIFO/FIFO[116][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[116][2]  ( .D(n1065), .E(n1977), .C(inClock), .Q(
        \u_inFIFO/FIFO[116][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[116][3]  ( .D(n1081), .E(n1977), .C(inClock), .Q(
        \u_inFIFO/FIFO[116][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[117][0]  ( .D(n1033), .E(n1976), .C(inClock), .Q(
        \u_inFIFO/FIFO[117][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[117][1]  ( .D(n1049), .E(n1976), .C(inClock), .Q(
        \u_inFIFO/FIFO[117][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[117][2]  ( .D(n1065), .E(n1976), .C(inClock), .Q(
        \u_inFIFO/FIFO[117][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[117][3]  ( .D(n1081), .E(n1976), .C(inClock), .Q(
        \u_inFIFO/FIFO[117][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[119][0]  ( .D(n1033), .E(n1974), .C(inClock), .Q(
        \u_inFIFO/FIFO[119][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[119][1]  ( .D(n1049), .E(n1974), .C(inClock), .Q(
        \u_inFIFO/FIFO[119][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[119][2]  ( .D(n1065), .E(n1974), .C(inClock), .Q(
        \u_inFIFO/FIFO[119][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[119][3]  ( .D(n1081), .E(n1974), .C(inClock), .Q(
        \u_inFIFO/FIFO[119][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[120][0]  ( .D(n1034), .E(n1973), .C(inClock), .Q(
        \u_inFIFO/FIFO[120][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[120][1]  ( .D(n1050), .E(n1973), .C(inClock), .Q(
        \u_inFIFO/FIFO[120][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[120][2]  ( .D(n1066), .E(n1973), .C(inClock), .Q(
        \u_inFIFO/FIFO[120][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[120][3]  ( .D(n1082), .E(n1973), .C(inClock), .Q(
        \u_inFIFO/FIFO[120][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[121][0]  ( .D(n1034), .E(n1972), .C(inClock), .Q(
        \u_inFIFO/FIFO[121][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[121][1]  ( .D(n1050), .E(n1972), .C(inClock), .Q(
        \u_inFIFO/FIFO[121][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[121][2]  ( .D(n1066), .E(n1972), .C(inClock), .Q(
        \u_inFIFO/FIFO[121][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[121][3]  ( .D(n1082), .E(n1972), .C(inClock), .Q(
        \u_inFIFO/FIFO[121][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[123][0]  ( .D(n1034), .E(n1970), .C(inClock), .Q(
        \u_inFIFO/FIFO[123][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[123][1]  ( .D(n1050), .E(n1970), .C(inClock), .Q(
        \u_inFIFO/FIFO[123][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[123][2]  ( .D(n1066), .E(n1970), .C(inClock), .Q(
        \u_inFIFO/FIFO[123][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[123][3]  ( .D(n1082), .E(n1970), .C(inClock), .Q(
        \u_inFIFO/FIFO[123][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[124][0]  ( .D(n1034), .E(n1969), .C(inClock), .Q(
        \u_inFIFO/FIFO[124][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[124][1]  ( .D(n1050), .E(n1969), .C(inClock), .Q(
        \u_inFIFO/FIFO[124][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[124][2]  ( .D(n1066), .E(n1969), .C(inClock), .Q(
        \u_inFIFO/FIFO[124][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[124][3]  ( .D(n1082), .E(n1969), .C(inClock), .Q(
        \u_inFIFO/FIFO[124][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[125][0]  ( .D(n1034), .E(n1968), .C(inClock), .Q(
        \u_inFIFO/FIFO[125][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[125][1]  ( .D(n1050), .E(n1968), .C(inClock), .Q(
        \u_inFIFO/FIFO[125][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[125][2]  ( .D(n1066), .E(n1968), .C(inClock), .Q(
        \u_inFIFO/FIFO[125][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[125][3]  ( .D(n1082), .E(n1968), .C(inClock), .Q(
        \u_inFIFO/FIFO[125][3] ) );
  DFE1 \u_inFIFO/FIFO_reg[127][0]  ( .D(n1034), .E(n1966), .C(inClock), .Q(
        \u_inFIFO/FIFO[127][0] ) );
  DFE1 \u_inFIFO/FIFO_reg[127][1]  ( .D(n1050), .E(n1966), .C(inClock), .Q(
        \u_inFIFO/FIFO[127][1] ) );
  DFE1 \u_inFIFO/FIFO_reg[127][2]  ( .D(n1066), .E(n1966), .C(inClock), .Q(
        \u_inFIFO/FIFO[127][2] ) );
  DFE1 \u_inFIFO/FIFO_reg[127][3]  ( .D(n1082), .E(n1966), .C(inClock), .Q(
        \u_inFIFO/FIFO[127][3] ) );
  DFE1 \u_coder/my_clk_10M_reg  ( .D(\u_coder/clk_10M ), .E(n1231), .C(inClock), .Q(\u_coder/my_clk_10M ), .QN(\u_coder/n88 ) );
  DFE1 \u_cordic/my_rotation/present_angle_reg[1][13]  ( .D(
        \u_cordic/my_rotation/present_angle[0][13] ), .E(n1231), .C(inClock), 
        .QN(n172) );
  DFE1 \u_cordic/my_rotation/present_angle_reg[1][14]  ( .D(
        \u_cordic/my_rotation/present_angle[0][14] ), .E(n1231), .C(inClock), 
        .QN(n171) );
  DFE1 \u_cordic/my_rotation/present_angle_reg[1][15]  ( .D(
        \u_cordic/my_rotation/present_angle[0][15] ), .E(n1231), .C(inClock), 
        .QN(n193) );
  DFE1 \u_cordic/my_rotation/present_angle_reg[1][11]  ( .D(
        \u_cordic/my_rotation/present_angle[0][11] ), .E(n1231), .C(inClock), 
        .QN(n134) );
  DFE1 \u_cordic/my_rotation/present_angle_reg[1][12]  ( .D(
        \u_cordic/my_rotation/present_angle[0][12] ), .E(n1231), .C(inClock), 
        .QN(n133) );
  DFE1 \u_cordic/my_rotation/present_angle_reg[1][8]  ( .D(
        \u_cordic/my_rotation/present_angle[0][8] ), .E(n1231), .C(inClock), 
        .QN(n87) );
  DFE1 \u_cordic/my_rotation/present_angle_reg[1][9]  ( .D(
        \u_cordic/my_rotation/present_angle[0][9] ), .E(n1231), .C(inClock), 
        .QN(n86) );
  DFE1 \u_cordic/my_rotation/present_angle_reg[1][10]  ( .D(
        \u_cordic/my_rotation/present_angle[0][10] ), .E(n1231), .C(inClock), 
        .QN(n85) );
  DFE1 \u_cordic/my_rotation/present_angle_reg[1][6]  ( .D(
        \u_cordic/my_rotation/present_angle[0][6] ), .E(n1231), .C(inClock), 
        .QN(n72) );
  DFE1 \u_cordic/my_rotation/present_angle_reg[1][7]  ( .D(
        \u_cordic/my_rotation/present_angle[0][7] ), .E(n1231), .C(inClock), 
        .QN(n71) );
  DFE1 \u_cordic/my_rotation/present_angle_reg[1][3]  ( .D(
        \u_cordic/my_rotation/present_angle[0][3] ), .E(n1231), .C(inClock), 
        .QN(n21) );
  DFE1 \u_cordic/my_rotation/present_angle_reg[1][4]  ( .D(
        \u_cordic/my_rotation/present_angle[0][4] ), .E(n1231), .C(inClock), 
        .QN(n66) );
  DFE1 \u_cordic/my_rotation/present_angle_reg[1][5]  ( .D(
        \u_cordic/my_rotation/present_angle[0][5] ), .E(n1231), .C(inClock), 
        .QN(n73) );
  DFE1 \u_cordic/my_rotation/present_angle_reg[1][0]  ( .D(
        \u_cordic/my_rotation/present_angle[0][0] ), .E(n1231), .C(inClock), 
        .QN(n65) );
  DFE1 \u_cordic/my_rotation/present_angle_reg[1][1]  ( .D(
        \u_cordic/my_rotation/present_angle[0][1] ), .E(n1231), .C(inClock), 
        .QN(n64) );
  DFE1 \u_cordic/my_rotation/present_angle_reg[1][2]  ( .D(
        \u_cordic/my_rotation/present_angle[0][2] ), .E(n1231), .C(inClock), 
        .QN(n63) );
  NOR21 \u_decoder/iq_demod/cossin_dig/U51  ( .A(
        \u_decoder/iq_demod/cossin_dig/N55 ), .B(
        \u_decoder/iq_demod/cossin_dig/n54 ), .Q(
        \u_decoder/iq_demod/cossin_dig/N60 ) );
  NOR21 \u_decoder/iq_demod/cossin_dig/U49  ( .A(
        \u_decoder/iq_demod/cossin_dig/n21 ), .B(
        \u_decoder/iq_demod/cossin_dig/n19 ), .Q(
        \u_decoder/iq_demod/cossin_dig/N52 ) );
  NAND22 \u_cordic/mycordic/U561  ( .A(\u_cordic/mycordic/N619 ), .B(n758), 
        .Q(\u_cordic/mycordic/n564 ) );
  NAND22 \u_cordic/mycordic/U559  ( .A(
        \u_cordic/mycordic/present_ANGLE_table[6][2] ), .B(n758), .Q(
        \u_cordic/mycordic/n560 ) );
  NAND22 \u_cordic/mycordic/U557  ( .A(\u_cordic/mycordic/N615 ), .B(n758), 
        .Q(\u_cordic/mycordic/n556 ) );
  NAND22 \u_cordic/mycordic/U560  ( .A(n305), .B(n757), .Q(
        \u_cordic/mycordic/n562 ) );
  NAND22 \u_cordic/mycordic/U558  ( .A(
        \u_cordic/mycordic/present_ANGLE_table[6][1] ), .B(n757), .Q(
        \u_cordic/mycordic/n558 ) );
  NAND22 \u_decoder/iq_demod/cossin_dig/U50  ( .A(
        \u_decoder/iq_demod/cossin_dig/N55 ), .B(
        \u_decoder/iq_demod/cossin_dig/n19 ), .Q(
        \u_decoder/iq_demod/cossin_dig/n55 ) );
  IMUX21 \u_cordic/mycordic/U535  ( .A(\u_cordic/mycordic/n568 ), .B(n392), 
        .S(n766), .Q(\u_cordic/mycordic/n567 ) );
  MUX22 \u_cordic/mycordic/U536  ( .A(
        \u_cordic/mycordic/present_ANGLE_table[6][6] ), .B(
        \u_cordic/mycordic/n567 ), .S(n384), .Q(
        \u_cordic/mycordic/next_ANGLE_table[6][6] ) );
  IMUX21 \u_cordic/mycordic/U533  ( .A(\u_cordic/mycordic/n566 ), .B(n390), 
        .S(n766), .Q(\u_cordic/mycordic/n565 ) );
  MUX22 \u_cordic/mycordic/U534  ( .A(
        \u_cordic/mycordic/present_ANGLE_table[6][5] ), .B(
        \u_cordic/mycordic/n565 ), .S(n384), .Q(
        \u_cordic/mycordic/next_ANGLE_table[6][5] ) );
  IMUX21 \u_cordic/mycordic/U531  ( .A(\u_cordic/mycordic/n564 ), .B(n386), 
        .S(n766), .Q(\u_cordic/mycordic/n563 ) );
  MUX22 \u_cordic/mycordic/U532  ( .A(
        \u_cordic/mycordic/present_ANGLE_table[6][4] ), .B(
        \u_cordic/mycordic/n563 ), .S(n384), .Q(
        \u_cordic/mycordic/next_ANGLE_table[6][4] ) );
  IMUX21 \u_cordic/mycordic/U529  ( .A(\u_cordic/mycordic/n562 ), .B(n393), 
        .S(n766), .Q(\u_cordic/mycordic/n561 ) );
  MUX22 \u_cordic/mycordic/U530  ( .A(
        \u_cordic/mycordic/present_ANGLE_table[6][3] ), .B(
        \u_cordic/mycordic/n561 ), .S(n384), .Q(
        \u_cordic/mycordic/next_ANGLE_table[6][3] ) );
  IMUX40 \u_outFIFO/U1411  ( .A(\u_outFIFO/n1409 ), .B(\u_outFIFO/n1399 ), .C(
        \u_outFIFO/n1404 ), .D(\u_outFIFO/n1394 ), .S0(n761), .S1(
        \u_outFIFO/N43 ), .Q(\u_outFIFO/n1435 ) );
  IMUX21 \u_outFIFO/U1367  ( .A(\u_outFIFO/n1434 ), .B(\u_outFIFO/n1435 ), .S(
        \u_outFIFO/N45 ), .Q(\u_outFIFO/N205 ) );
  IMUX40 \u_outFIFO/U1445  ( .A(\u_outFIFO/n1451 ), .B(\u_outFIFO/n1441 ), .C(
        \u_outFIFO/n1446 ), .D(\u_outFIFO/n1436 ), .S0(n761), .S1(
        \u_outFIFO/N43 ), .Q(\u_outFIFO/n1477 ) );
  IMUX21 \u_outFIFO/U1376  ( .A(\u_outFIFO/n1476 ), .B(\u_outFIFO/n1477 ), .S(
        \u_outFIFO/N45 ), .Q(\u_outFIFO/N204 ) );
  IMUX40 \u_outFIFO/U1479  ( .A(\u_outFIFO/n1493 ), .B(\u_outFIFO/n1483 ), .C(
        \u_outFIFO/n1488 ), .D(\u_outFIFO/n1478 ), .S0(n761), .S1(
        \u_outFIFO/N43 ), .Q(\u_outFIFO/n1519 ) );
  IMUX21 \u_outFIFO/U1385  ( .A(\u_outFIFO/n1518 ), .B(\u_outFIFO/n1519 ), .S(
        \u_outFIFO/N45 ), .Q(\u_outFIFO/N203 ) );
  IMUX40 \u_outFIFO/U1513  ( .A(\u_outFIFO/n1535 ), .B(\u_outFIFO/n1525 ), .C(
        \u_outFIFO/n1530 ), .D(\u_outFIFO/n1520 ), .S0(n761), .S1(
        \u_outFIFO/N43 ), .Q(\u_outFIFO/n1561 ) );
  IMUX21 \u_outFIFO/U1394  ( .A(\u_outFIFO/n1560 ), .B(\u_outFIFO/n1561 ), .S(
        \u_outFIFO/N45 ), .Q(\u_outFIFO/N202 ) );
  IMUX21 \u_cordic/mycordic/U527  ( .A(\u_cordic/mycordic/n560 ), .B(
        \u_cordic/mycordic/present_ANGLE_table[6][2] ), .S(n766), .Q(
        \u_cordic/mycordic/n559 ) );
  MUX22 \u_cordic/mycordic/U528  ( .A(
        \u_cordic/mycordic/present_ANGLE_table[6][2] ), .B(
        \u_cordic/mycordic/n559 ), .S(n384), .Q(
        \u_cordic/mycordic/next_ANGLE_table[6][2] ) );
  IMUX21 \u_cordic/mycordic/U537  ( .A(\u_cordic/mycordic/n570 ), .B(n388), 
        .S(n766), .Q(\u_cordic/mycordic/n569 ) );
  MUX22 \u_cordic/mycordic/U538  ( .A(
        \u_cordic/mycordic/present_ANGLE_table[6][7] ), .B(
        \u_cordic/mycordic/n569 ), .S(n384), .Q(
        \u_cordic/mycordic/next_ANGLE_table[6][7] ) );
  IMUX21 \u_cordic/mycordic/U525  ( .A(\u_cordic/mycordic/n558 ), .B(n314), 
        .S(n766), .Q(\u_cordic/mycordic/n557 ) );
  MUX22 \u_cordic/mycordic/U526  ( .A(
        \u_cordic/mycordic/present_ANGLE_table[6][1] ), .B(
        \u_cordic/mycordic/n557 ), .S(n384), .Q(
        \u_cordic/mycordic/next_ANGLE_table[6][1] ) );
  IMUX21 \u_cordic/mycordic/U523  ( .A(\u_cordic/mycordic/n556 ), .B(n313), 
        .S(n766), .Q(\u_cordic/mycordic/n555 ) );
  MUX22 \u_cordic/mycordic/U524  ( .A(\u_cordic/mycordic/N615 ), .B(
        \u_cordic/mycordic/n555 ), .S(n384), .Q(
        \u_cordic/mycordic/next_ANGLE_table[6][0] ) );
  NAND22 \u_cordic/mycordic/U565  ( .A(\u_cordic/mycordic/N623 ), .B(n758), 
        .Q(\u_cordic/mycordic/n572 ) );
  NAND22 \u_cordic/mycordic/U563  ( .A(\u_cordic/mycordic/N621 ), .B(n758), 
        .Q(\u_cordic/mycordic/n568 ) );
  NAND22 \u_cordic/mycordic/U564  ( .A(\u_cordic/mycordic/N622 ), .B(n757), 
        .Q(\u_cordic/mycordic/n570 ) );
  NAND22 \u_cordic/mycordic/U562  ( .A(\u_cordic/mycordic/N620 ), .B(n757), 
        .Q(\u_cordic/mycordic/n566 ) );
  XOR21 \u_cordic/mycordic/U555  ( .A(\u_cordic/mycordic/n110 ), .B(
        \u_cordic/mycordic/present_C_table[7][0] ), .Q(
        \u_cordic/mycordic/n587 ) );
  NAND22 \u_decoder/iq_demod/cossin_dig/U52  ( .A(
        \u_decoder/iq_demod/cossin_dig/n21 ), .B(
        \u_decoder/iq_demod/cossin_dig/n54 ), .Q(
        \u_decoder/iq_demod/cossin_dig/n56 ) );
  IMUX40 \u_outFIFO/U1422  ( .A(\u_outFIFO/FIFO[20][0] ), .B(
        \u_outFIFO/FIFO[21][0] ), .C(\u_outFIFO/FIFO[22][0] ), .D(
        \u_outFIFO/FIFO[23][0] ), .S0(n1179), .S1(n760), .Q(\u_outFIFO/n1427 )
         );
  IMUX40 \u_outFIFO/U1414  ( .A(\u_outFIFO/FIFO[52][0] ), .B(
        \u_outFIFO/FIFO[53][0] ), .C(\u_outFIFO/FIFO[54][0] ), .D(
        \u_outFIFO/FIFO[55][0] ), .S0(n759), .S1(n760), .Q(\u_outFIFO/n1417 )
         );
  IMUX40 \u_outFIFO/U1418  ( .A(\u_outFIFO/FIFO[36][0] ), .B(
        \u_outFIFO/FIFO[37][0] ), .C(\u_outFIFO/FIFO[38][0] ), .D(
        \u_outFIFO/FIFO[39][0] ), .S0(n1179), .S1(\u_outFIFO/N40 ), .Q(
        \u_outFIFO/n1422 ) );
  IMUX40 \u_outFIFO/U1456  ( .A(\u_outFIFO/FIFO[20][1] ), .B(
        \u_outFIFO/FIFO[21][1] ), .C(\u_outFIFO/FIFO[22][1] ), .D(
        \u_outFIFO/FIFO[23][1] ), .S0(n1177), .S1(\u_outFIFO/N40 ), .Q(
        \u_outFIFO/n1469 ) );
  IMUX40 \u_outFIFO/U1448  ( .A(\u_outFIFO/FIFO[52][1] ), .B(
        \u_outFIFO/FIFO[53][1] ), .C(\u_outFIFO/FIFO[54][1] ), .D(
        \u_outFIFO/FIFO[55][1] ), .S0(\u_outFIFO/N39 ), .S1(\u_outFIFO/N40 ), 
        .Q(\u_outFIFO/n1459 ) );
  IMUX40 \u_outFIFO/U1452  ( .A(\u_outFIFO/FIFO[36][1] ), .B(
        \u_outFIFO/FIFO[37][1] ), .C(\u_outFIFO/FIFO[38][1] ), .D(
        \u_outFIFO/FIFO[39][1] ), .S0(n1180), .S1(n1182), .Q(\u_outFIFO/n1464 ) );
  IMUX40 \u_outFIFO/U1490  ( .A(\u_outFIFO/FIFO[20][2] ), .B(
        \u_outFIFO/FIFO[21][2] ), .C(\u_outFIFO/FIFO[22][2] ), .D(
        \u_outFIFO/FIFO[23][2] ), .S0(n1180), .S1(n760), .Q(\u_outFIFO/n1511 )
         );
  IMUX40 \u_outFIFO/U1482  ( .A(\u_outFIFO/FIFO[52][2] ), .B(
        \u_outFIFO/FIFO[53][2] ), .C(\u_outFIFO/FIFO[54][2] ), .D(
        \u_outFIFO/FIFO[55][2] ), .S0(n1179), .S1(n760), .Q(\u_outFIFO/n1501 )
         );
  IMUX40 \u_outFIFO/U1486  ( .A(\u_outFIFO/FIFO[36][2] ), .B(
        \u_outFIFO/FIFO[37][2] ), .C(\u_outFIFO/FIFO[38][2] ), .D(
        \u_outFIFO/FIFO[39][2] ), .S0(n1180), .S1(n760), .Q(\u_outFIFO/n1506 )
         );
  IMUX40 \u_outFIFO/U1524  ( .A(\u_outFIFO/FIFO[20][3] ), .B(
        \u_outFIFO/FIFO[21][3] ), .C(\u_outFIFO/FIFO[22][3] ), .D(
        \u_outFIFO/FIFO[23][3] ), .S0(n1176), .S1(\u_outFIFO/N40 ), .Q(
        \u_outFIFO/n1553 ) );
  IMUX40 \u_outFIFO/U1516  ( .A(\u_outFIFO/FIFO[52][3] ), .B(
        \u_outFIFO/FIFO[53][3] ), .C(\u_outFIFO/FIFO[54][3] ), .D(
        \u_outFIFO/FIFO[55][3] ), .S0(n759), .S1(\u_outFIFO/N40 ), .Q(
        \u_outFIFO/n1543 ) );
  IMUX40 \u_outFIFO/U1520  ( .A(\u_outFIFO/FIFO[36][3] ), .B(
        \u_outFIFO/FIFO[37][3] ), .C(\u_outFIFO/FIFO[38][3] ), .D(
        \u_outFIFO/FIFO[39][3] ), .S0(n1176), .S1(n1181), .Q(\u_outFIFO/n1548 ) );
  IMUX40 \u_outFIFO/U1406  ( .A(\u_outFIFO/FIFO[80][0] ), .B(
        \u_outFIFO/FIFO[81][0] ), .C(\u_outFIFO/FIFO[82][0] ), .D(
        \u_outFIFO/FIFO[83][0] ), .S0(n1179), .S1(\u_outFIFO/N40 ), .Q(
        \u_outFIFO/n1405 ) );
  IMUX40 \u_outFIFO/U1404  ( .A(\u_outFIFO/FIFO[88][0] ), .B(
        \u_outFIFO/FIFO[89][0] ), .C(\u_outFIFO/FIFO[90][0] ), .D(
        \u_outFIFO/FIFO[91][0] ), .S0(\u_outFIFO/N39 ), .S1(\u_outFIFO/N40 ), 
        .Q(\u_outFIFO/n1406 ) );
  IMUX40 \u_outFIFO/U1405  ( .A(\u_outFIFO/FIFO[84][0] ), .B(
        \u_outFIFO/FIFO[85][0] ), .C(\u_outFIFO/FIFO[86][0] ), .D(
        \u_outFIFO/FIFO[87][0] ), .S0(n1177), .S1(n1182), .Q(\u_outFIFO/n1407 ) );
  IMUX40 \u_outFIFO/U1361  ( .A(\u_outFIFO/n1405 ), .B(\u_outFIFO/n1406 ), .C(
        \u_outFIFO/n1407 ), .D(\u_outFIFO/n1408 ), .S0(n1183), .S1(n14), .Q(
        \u_outFIFO/n1404 ) );
  IMUX40 \u_outFIFO/U1440  ( .A(\u_outFIFO/FIFO[80][1] ), .B(
        \u_outFIFO/FIFO[81][1] ), .C(\u_outFIFO/FIFO[82][1] ), .D(
        \u_outFIFO/FIFO[83][1] ), .S0(n1178), .S1(\u_outFIFO/N40 ), .Q(
        \u_outFIFO/n1447 ) );
  IMUX40 \u_outFIFO/U1438  ( .A(\u_outFIFO/FIFO[88][1] ), .B(
        \u_outFIFO/FIFO[89][1] ), .C(\u_outFIFO/FIFO[90][1] ), .D(
        \u_outFIFO/FIFO[91][1] ), .S0(n1178), .S1(\u_outFIFO/N40 ), .Q(
        \u_outFIFO/n1448 ) );
  IMUX40 \u_outFIFO/U1439  ( .A(\u_outFIFO/FIFO[84][1] ), .B(
        \u_outFIFO/FIFO[85][1] ), .C(\u_outFIFO/FIFO[86][1] ), .D(
        \u_outFIFO/FIFO[87][1] ), .S0(n1178), .S1(\u_outFIFO/N40 ), .Q(
        \u_outFIFO/n1449 ) );
  IMUX40 \u_outFIFO/U1370  ( .A(\u_outFIFO/n1447 ), .B(\u_outFIFO/n1448 ), .C(
        \u_outFIFO/n1449 ), .D(\u_outFIFO/n1450 ), .S0(\u_outFIFO/N42 ), .S1(
        n14), .Q(\u_outFIFO/n1446 ) );
  IMUX40 \u_outFIFO/U1474  ( .A(\u_outFIFO/FIFO[80][2] ), .B(
        \u_outFIFO/FIFO[81][2] ), .C(\u_outFIFO/FIFO[82][2] ), .D(
        \u_outFIFO/FIFO[83][2] ), .S0(n759), .S1(n1181), .Q(\u_outFIFO/n1489 )
         );
  IMUX40 \u_outFIFO/U1472  ( .A(\u_outFIFO/FIFO[88][2] ), .B(
        \u_outFIFO/FIFO[89][2] ), .C(\u_outFIFO/FIFO[90][2] ), .D(
        \u_outFIFO/FIFO[91][2] ), .S0(n759), .S1(n1181), .Q(\u_outFIFO/n1490 )
         );
  IMUX40 \u_outFIFO/U1473  ( .A(\u_outFIFO/FIFO[84][2] ), .B(
        \u_outFIFO/FIFO[85][2] ), .C(\u_outFIFO/FIFO[86][2] ), .D(
        \u_outFIFO/FIFO[87][2] ), .S0(n759), .S1(n1181), .Q(\u_outFIFO/n1491 )
         );
  IMUX40 \u_outFIFO/U1379  ( .A(\u_outFIFO/n1489 ), .B(\u_outFIFO/n1490 ), .C(
        \u_outFIFO/n1491 ), .D(\u_outFIFO/n1492 ), .S0(\u_outFIFO/N42 ), .S1(
        n14), .Q(\u_outFIFO/n1488 ) );
  IMUX40 \u_outFIFO/U1508  ( .A(\u_outFIFO/FIFO[80][3] ), .B(
        \u_outFIFO/FIFO[81][3] ), .C(\u_outFIFO/FIFO[82][3] ), .D(
        \u_outFIFO/FIFO[83][3] ), .S0(n1179), .S1(\u_outFIFO/N40 ), .Q(
        \u_outFIFO/n1531 ) );
  IMUX40 \u_outFIFO/U1506  ( .A(\u_outFIFO/FIFO[88][3] ), .B(
        \u_outFIFO/FIFO[89][3] ), .C(\u_outFIFO/FIFO[90][3] ), .D(
        \u_outFIFO/FIFO[91][3] ), .S0(\u_outFIFO/N39 ), .S1(\u_outFIFO/N40 ), 
        .Q(\u_outFIFO/n1532 ) );
  IMUX40 \u_outFIFO/U1507  ( .A(\u_outFIFO/FIFO[84][3] ), .B(
        \u_outFIFO/FIFO[85][3] ), .C(\u_outFIFO/FIFO[86][3] ), .D(
        \u_outFIFO/FIFO[87][3] ), .S0(n1177), .S1(\u_outFIFO/N40 ), .Q(
        \u_outFIFO/n1533 ) );
  IMUX40 \u_outFIFO/U1388  ( .A(\u_outFIFO/n1531 ), .B(\u_outFIFO/n1532 ), .C(
        \u_outFIFO/n1533 ), .D(\u_outFIFO/n1534 ), .S0(\u_outFIFO/N42 ), .S1(
        n14), .Q(\u_outFIFO/n1530 ) );
  IMUX40 \u_outFIFO/U1421  ( .A(\u_outFIFO/FIFO[24][0] ), .B(
        \u_outFIFO/FIFO[25][0] ), .C(\u_outFIFO/FIFO[26][0] ), .D(
        \u_outFIFO/FIFO[27][0] ), .S0(n1179), .S1(n1181), .Q(\u_outFIFO/n1426 ) );
  IMUX40 \u_outFIFO/U1423  ( .A(\u_outFIFO/FIFO[16][0] ), .B(
        \u_outFIFO/FIFO[17][0] ), .C(\u_outFIFO/FIFO[18][0] ), .D(
        \u_outFIFO/FIFO[19][0] ), .S0(n1179), .S1(n760), .Q(\u_outFIFO/n1425 )
         );
  IMUX40 \u_outFIFO/U1420  ( .A(\u_outFIFO/FIFO[28][0] ), .B(
        \u_outFIFO/FIFO[29][0] ), .C(\u_outFIFO/FIFO[30][0] ), .D(
        \u_outFIFO/FIFO[31][0] ), .S0(n1179), .S1(n1181), .Q(\u_outFIFO/n1428 ) );
  IMUX40 \u_outFIFO/U1413  ( .A(\u_outFIFO/FIFO[56][0] ), .B(
        \u_outFIFO/FIFO[57][0] ), .C(\u_outFIFO/FIFO[58][0] ), .D(
        \u_outFIFO/FIFO[59][0] ), .S0(n1178), .S1(\u_outFIFO/N40 ), .Q(
        \u_outFIFO/n1416 ) );
  IMUX40 \u_outFIFO/U1415  ( .A(\u_outFIFO/FIFO[48][0] ), .B(
        \u_outFIFO/FIFO[49][0] ), .C(\u_outFIFO/FIFO[50][0] ), .D(
        \u_outFIFO/FIFO[51][0] ), .S0(n1176), .S1(n760), .Q(\u_outFIFO/n1415 )
         );
  IMUX40 \u_outFIFO/U1412  ( .A(\u_outFIFO/FIFO[60][0] ), .B(
        \u_outFIFO/FIFO[61][0] ), .C(\u_outFIFO/FIFO[62][0] ), .D(
        \u_outFIFO/FIFO[63][0] ), .S0(n1179), .S1(n760), .Q(\u_outFIFO/n1418 )
         );
  IMUX40 \u_outFIFO/U1417  ( .A(\u_outFIFO/FIFO[40][0] ), .B(
        \u_outFIFO/FIFO[41][0] ), .C(\u_outFIFO/FIFO[42][0] ), .D(
        \u_outFIFO/FIFO[43][0] ), .S0(n1179), .S1(n1182), .Q(\u_outFIFO/n1421 ) );
  IMUX40 \u_outFIFO/U1419  ( .A(\u_outFIFO/FIFO[32][0] ), .B(
        \u_outFIFO/FIFO[33][0] ), .C(\u_outFIFO/FIFO[34][0] ), .D(
        \u_outFIFO/FIFO[35][0] ), .S0(n1179), .S1(n1182), .Q(\u_outFIFO/n1420 ) );
  IMUX40 \u_outFIFO/U1416  ( .A(\u_outFIFO/FIFO[44][0] ), .B(
        \u_outFIFO/FIFO[45][0] ), .C(\u_outFIFO/FIFO[46][0] ), .D(
        \u_outFIFO/FIFO[47][0] ), .S0(n1179), .S1(n760), .Q(\u_outFIFO/n1423 )
         );
  IMUX40 \u_outFIFO/U1424  ( .A(\u_outFIFO/FIFO[12][0] ), .B(
        \u_outFIFO/FIFO[13][0] ), .C(\u_outFIFO/FIFO[14][0] ), .D(
        \u_outFIFO/FIFO[15][0] ), .S0(n1179), .S1(n1182), .Q(\u_outFIFO/n1433 ) );
  IMUX40 \u_outFIFO/U1455  ( .A(\u_outFIFO/FIFO[24][1] ), .B(
        \u_outFIFO/FIFO[25][1] ), .C(\u_outFIFO/FIFO[26][1] ), .D(
        \u_outFIFO/FIFO[27][1] ), .S0(n1177), .S1(\u_outFIFO/N40 ), .Q(
        \u_outFIFO/n1468 ) );
  IMUX40 \u_outFIFO/U1457  ( .A(\u_outFIFO/FIFO[16][1] ), .B(
        \u_outFIFO/FIFO[17][1] ), .C(\u_outFIFO/FIFO[18][1] ), .D(
        \u_outFIFO/FIFO[19][1] ), .S0(n1177), .S1(n760), .Q(\u_outFIFO/n1467 )
         );
  IMUX40 \u_outFIFO/U1454  ( .A(\u_outFIFO/FIFO[28][1] ), .B(
        \u_outFIFO/FIFO[29][1] ), .C(\u_outFIFO/FIFO[30][1] ), .D(
        \u_outFIFO/FIFO[31][1] ), .S0(n1177), .S1(n1182), .Q(\u_outFIFO/n1470 ) );
  IMUX40 \u_outFIFO/U1447  ( .A(\u_outFIFO/FIFO[56][1] ), .B(
        \u_outFIFO/FIFO[57][1] ), .C(\u_outFIFO/FIFO[58][1] ), .D(
        \u_outFIFO/FIFO[59][1] ), .S0(\u_outFIFO/N39 ), .S1(\u_outFIFO/N40 ), 
        .Q(\u_outFIFO/n1458 ) );
  IMUX40 \u_outFIFO/U1449  ( .A(\u_outFIFO/FIFO[48][1] ), .B(
        \u_outFIFO/FIFO[49][1] ), .C(\u_outFIFO/FIFO[50][1] ), .D(
        \u_outFIFO/FIFO[51][1] ), .S0(\u_outFIFO/N39 ), .S1(n1181), .Q(
        \u_outFIFO/n1457 ) );
  IMUX40 \u_outFIFO/U1446  ( .A(\u_outFIFO/FIFO[60][1] ), .B(
        \u_outFIFO/FIFO[61][1] ), .C(\u_outFIFO/FIFO[62][1] ), .D(
        \u_outFIFO/FIFO[63][1] ), .S0(\u_outFIFO/N39 ), .S1(\u_outFIFO/N40 ), 
        .Q(\u_outFIFO/n1460 ) );
  IMUX40 \u_outFIFO/U1451  ( .A(\u_outFIFO/FIFO[40][1] ), .B(
        \u_outFIFO/FIFO[41][1] ), .C(\u_outFIFO/FIFO[42][1] ), .D(
        \u_outFIFO/FIFO[43][1] ), .S0(\u_outFIFO/N39 ), .S1(\u_outFIFO/N40 ), 
        .Q(\u_outFIFO/n1463 ) );
  IMUX40 \u_outFIFO/U1453  ( .A(\u_outFIFO/FIFO[32][1] ), .B(
        \u_outFIFO/FIFO[33][1] ), .C(\u_outFIFO/FIFO[34][1] ), .D(
        \u_outFIFO/FIFO[35][1] ), .S0(\u_outFIFO/N39 ), .S1(n1181), .Q(
        \u_outFIFO/n1462 ) );
  IMUX40 \u_outFIFO/U1450  ( .A(\u_outFIFO/FIFO[44][1] ), .B(
        \u_outFIFO/FIFO[45][1] ), .C(\u_outFIFO/FIFO[46][1] ), .D(
        \u_outFIFO/FIFO[47][1] ), .S0(\u_outFIFO/N39 ), .S1(\u_outFIFO/N40 ), 
        .Q(\u_outFIFO/n1465 ) );
  IMUX40 \u_outFIFO/U1458  ( .A(\u_outFIFO/FIFO[12][1] ), .B(
        \u_outFIFO/FIFO[13][1] ), .C(\u_outFIFO/FIFO[14][1] ), .D(
        \u_outFIFO/FIFO[15][1] ), .S0(n1177), .S1(\u_outFIFO/N40 ), .Q(
        \u_outFIFO/n1475 ) );
  IMUX40 \u_outFIFO/U1489  ( .A(\u_outFIFO/FIFO[24][2] ), .B(
        \u_outFIFO/FIFO[25][2] ), .C(\u_outFIFO/FIFO[26][2] ), .D(
        \u_outFIFO/FIFO[27][2] ), .S0(n759), .S1(n760), .Q(\u_outFIFO/n1510 )
         );
  IMUX40 \u_outFIFO/U1491  ( .A(\u_outFIFO/FIFO[16][2] ), .B(
        \u_outFIFO/FIFO[17][2] ), .C(\u_outFIFO/FIFO[18][2] ), .D(
        \u_outFIFO/FIFO[19][2] ), .S0(n759), .S1(n760), .Q(\u_outFIFO/n1509 )
         );
  IMUX40 \u_outFIFO/U1488  ( .A(\u_outFIFO/FIFO[28][2] ), .B(
        \u_outFIFO/FIFO[29][2] ), .C(\u_outFIFO/FIFO[30][2] ), .D(
        \u_outFIFO/FIFO[31][2] ), .S0(n1177), .S1(n760), .Q(\u_outFIFO/n1512 )
         );
  IMUX40 \u_outFIFO/U1481  ( .A(\u_outFIFO/FIFO[56][2] ), .B(
        \u_outFIFO/FIFO[57][2] ), .C(\u_outFIFO/FIFO[58][2] ), .D(
        \u_outFIFO/FIFO[59][2] ), .S0(n759), .S1(n1181), .Q(\u_outFIFO/n1500 )
         );
  IMUX40 \u_outFIFO/U1483  ( .A(\u_outFIFO/FIFO[48][2] ), .B(
        \u_outFIFO/FIFO[49][2] ), .C(\u_outFIFO/FIFO[50][2] ), .D(
        \u_outFIFO/FIFO[51][2] ), .S0(n759), .S1(n760), .Q(\u_outFIFO/n1499 )
         );
  IMUX40 \u_outFIFO/U1480  ( .A(\u_outFIFO/FIFO[60][2] ), .B(
        \u_outFIFO/FIFO[61][2] ), .C(\u_outFIFO/FIFO[62][2] ), .D(
        \u_outFIFO/FIFO[63][2] ), .S0(\u_outFIFO/N39 ), .S1(n1181), .Q(
        \u_outFIFO/n1502 ) );
  IMUX40 \u_outFIFO/U1485  ( .A(\u_outFIFO/FIFO[40][2] ), .B(
        \u_outFIFO/FIFO[41][2] ), .C(\u_outFIFO/FIFO[42][2] ), .D(
        \u_outFIFO/FIFO[43][2] ), .S0(n1176), .S1(n760), .Q(\u_outFIFO/n1505 )
         );
  IMUX40 \u_outFIFO/U1487  ( .A(\u_outFIFO/FIFO[32][2] ), .B(
        \u_outFIFO/FIFO[33][2] ), .C(\u_outFIFO/FIFO[34][2] ), .D(
        \u_outFIFO/FIFO[35][2] ), .S0(n759), .S1(n760), .Q(\u_outFIFO/n1504 )
         );
  IMUX40 \u_outFIFO/U1484  ( .A(\u_outFIFO/FIFO[44][2] ), .B(
        \u_outFIFO/FIFO[45][2] ), .C(\u_outFIFO/FIFO[46][2] ), .D(
        \u_outFIFO/FIFO[47][2] ), .S0(\u_outFIFO/N39 ), .S1(n760), .Q(
        \u_outFIFO/n1507 ) );
  IMUX40 \u_outFIFO/U1492  ( .A(\u_outFIFO/FIFO[12][2] ), .B(
        \u_outFIFO/FIFO[13][2] ), .C(\u_outFIFO/FIFO[14][2] ), .D(
        \u_outFIFO/FIFO[15][2] ), .S0(\u_outFIFO/N39 ), .S1(n760), .Q(
        \u_outFIFO/n1517 ) );
  IMUX40 \u_outFIFO/U1523  ( .A(\u_outFIFO/FIFO[24][3] ), .B(
        \u_outFIFO/FIFO[25][3] ), .C(\u_outFIFO/FIFO[26][3] ), .D(
        \u_outFIFO/FIFO[27][3] ), .S0(n1176), .S1(n1181), .Q(\u_outFIFO/n1552 ) );
  IMUX40 \u_outFIFO/U1525  ( .A(\u_outFIFO/FIFO[16][3] ), .B(
        \u_outFIFO/FIFO[17][3] ), .C(\u_outFIFO/FIFO[18][3] ), .D(
        \u_outFIFO/FIFO[19][3] ), .S0(n1176), .S1(\u_outFIFO/N40 ), .Q(
        \u_outFIFO/n1551 ) );
  IMUX40 \u_outFIFO/U1522  ( .A(\u_outFIFO/FIFO[28][3] ), .B(
        \u_outFIFO/FIFO[29][3] ), .C(\u_outFIFO/FIFO[30][3] ), .D(
        \u_outFIFO/FIFO[31][3] ), .S0(n1176), .S1(n760), .Q(\u_outFIFO/n1554 )
         );
  IMUX40 \u_outFIFO/U1515  ( .A(\u_outFIFO/FIFO[56][3] ), .B(
        \u_outFIFO/FIFO[57][3] ), .C(\u_outFIFO/FIFO[58][3] ), .D(
        \u_outFIFO/FIFO[59][3] ), .S0(n1178), .S1(n1181), .Q(\u_outFIFO/n1542 ) );
  IMUX40 \u_outFIFO/U1517  ( .A(\u_outFIFO/FIFO[48][3] ), .B(
        \u_outFIFO/FIFO[49][3] ), .C(\u_outFIFO/FIFO[50][3] ), .D(
        \u_outFIFO/FIFO[51][3] ), .S0(n1176), .S1(n760), .Q(\u_outFIFO/n1541 )
         );
  IMUX40 \u_outFIFO/U1514  ( .A(\u_outFIFO/FIFO[60][3] ), .B(
        \u_outFIFO/FIFO[61][3] ), .C(\u_outFIFO/FIFO[62][3] ), .D(
        \u_outFIFO/FIFO[63][3] ), .S0(n1178), .S1(n1181), .Q(\u_outFIFO/n1544 ) );
  IMUX40 \u_outFIFO/U1519  ( .A(\u_outFIFO/FIFO[40][3] ), .B(
        \u_outFIFO/FIFO[41][3] ), .C(\u_outFIFO/FIFO[42][3] ), .D(
        \u_outFIFO/FIFO[43][3] ), .S0(n1176), .S1(\u_outFIFO/N40 ), .Q(
        \u_outFIFO/n1547 ) );
  IMUX40 \u_outFIFO/U1521  ( .A(\u_outFIFO/FIFO[32][3] ), .B(
        \u_outFIFO/FIFO[33][3] ), .C(\u_outFIFO/FIFO[34][3] ), .D(
        \u_outFIFO/FIFO[35][3] ), .S0(n1176), .S1(n1182), .Q(\u_outFIFO/n1546 ) );
  IMUX40 \u_outFIFO/U1518  ( .A(\u_outFIFO/FIFO[44][3] ), .B(
        \u_outFIFO/FIFO[45][3] ), .C(\u_outFIFO/FIFO[46][3] ), .D(
        \u_outFIFO/FIFO[47][3] ), .S0(n1176), .S1(\u_outFIFO/N40 ), .Q(
        \u_outFIFO/n1549 ) );
  IMUX40 \u_outFIFO/U1526  ( .A(\u_outFIFO/FIFO[12][3] ), .B(
        \u_outFIFO/FIFO[13][3] ), .C(\u_outFIFO/FIFO[14][3] ), .D(
        \u_outFIFO/FIFO[15][3] ), .S0(n1176), .S1(n1182), .Q(\u_outFIFO/n1559 ) );
  IMUX40 \u_outFIFO/U1402  ( .A(\u_outFIFO/FIFO[96][0] ), .B(
        \u_outFIFO/FIFO[97][0] ), .C(\u_outFIFO/FIFO[98][0] ), .D(
        \u_outFIFO/FIFO[99][0] ), .S0(n1180), .S1(\u_outFIFO/N40 ), .Q(
        \u_outFIFO/n1400 ) );
  IMUX40 \u_outFIFO/U1398  ( .A(\u_outFIFO/FIFO[112][0] ), .B(
        \u_outFIFO/FIFO[113][0] ), .C(\u_outFIFO/FIFO[114][0] ), .D(
        \u_outFIFO/FIFO[115][0] ), .S0(n1180), .S1(\u_outFIFO/N40 ), .Q(
        \u_outFIFO/n1395 ) );
  IMUX40 \u_outFIFO/U1403  ( .A(\u_outFIFO/FIFO[92][0] ), .B(
        \u_outFIFO/FIFO[93][0] ), .C(\u_outFIFO/FIFO[94][0] ), .D(
        \u_outFIFO/FIFO[95][0] ), .S0(n1176), .S1(n1182), .Q(\u_outFIFO/n1408 ) );
  IMUX40 \u_outFIFO/U1407  ( .A(\u_outFIFO/FIFO[76][0] ), .B(
        \u_outFIFO/FIFO[77][0] ), .C(\u_outFIFO/FIFO[78][0] ), .D(
        \u_outFIFO/FIFO[79][0] ), .S0(\u_outFIFO/N39 ), .S1(\u_outFIFO/N40 ), 
        .Q(\u_outFIFO/n1413 ) );
  IMUX40 \u_outFIFO/U1437  ( .A(\u_outFIFO/FIFO[92][1] ), .B(
        \u_outFIFO/FIFO[93][1] ), .C(\u_outFIFO/FIFO[94][1] ), .D(
        \u_outFIFO/FIFO[95][1] ), .S0(n1178), .S1(\u_outFIFO/N40 ), .Q(
        \u_outFIFO/n1450 ) );
  IMUX40 \u_outFIFO/U1433  ( .A(\u_outFIFO/FIFO[108][1] ), .B(
        \u_outFIFO/FIFO[109][1] ), .C(\u_outFIFO/FIFO[110][1] ), .D(
        \u_outFIFO/FIFO[111][1] ), .S0(n1178), .S1(n1182), .Q(
        \u_outFIFO/n1445 ) );
  IMUX40 \u_outFIFO/U1441  ( .A(\u_outFIFO/FIFO[76][1] ), .B(
        \u_outFIFO/FIFO[77][1] ), .C(\u_outFIFO/FIFO[78][1] ), .D(
        \u_outFIFO/FIFO[79][1] ), .S0(n1180), .S1(\u_outFIFO/N40 ), .Q(
        \u_outFIFO/n1455 ) );
  IMUX40 \u_outFIFO/U1432  ( .A(\u_outFIFO/FIFO[112][1] ), .B(
        \u_outFIFO/FIFO[113][1] ), .C(\u_outFIFO/FIFO[114][1] ), .D(
        \u_outFIFO/FIFO[115][1] ), .S0(n1178), .S1(n1182), .Q(
        \u_outFIFO/n1437 ) );
  IMUX40 \u_outFIFO/U1471  ( .A(\u_outFIFO/FIFO[92][2] ), .B(
        \u_outFIFO/FIFO[93][2] ), .C(\u_outFIFO/FIFO[94][2] ), .D(
        \u_outFIFO/FIFO[95][2] ), .S0(n1178), .S1(n1181), .Q(\u_outFIFO/n1492 ) );
  IMUX40 \u_outFIFO/U1467  ( .A(\u_outFIFO/FIFO[108][2] ), .B(
        \u_outFIFO/FIFO[109][2] ), .C(\u_outFIFO/FIFO[110][2] ), .D(
        \u_outFIFO/FIFO[111][2] ), .S0(n1180), .S1(n1181), .Q(
        \u_outFIFO/n1487 ) );
  IMUX40 \u_outFIFO/U1475  ( .A(\u_outFIFO/FIFO[76][2] ), .B(
        \u_outFIFO/FIFO[77][2] ), .C(\u_outFIFO/FIFO[78][2] ), .D(
        \u_outFIFO/FIFO[79][2] ), .S0(n1176), .S1(n1181), .Q(\u_outFIFO/n1497 ) );
  IMUX40 \u_outFIFO/U1466  ( .A(\u_outFIFO/FIFO[112][2] ), .B(
        \u_outFIFO/FIFO[113][2] ), .C(\u_outFIFO/FIFO[114][2] ), .D(
        \u_outFIFO/FIFO[115][2] ), .S0(n1177), .S1(n1181), .Q(
        \u_outFIFO/n1479 ) );
  IMUX40 \u_outFIFO/U1505  ( .A(\u_outFIFO/FIFO[92][3] ), .B(
        \u_outFIFO/FIFO[93][3] ), .C(\u_outFIFO/FIFO[94][3] ), .D(
        \u_outFIFO/FIFO[95][3] ), .S0(\u_outFIFO/N39 ), .S1(\u_outFIFO/N40 ), 
        .Q(\u_outFIFO/n1534 ) );
  IMUX40 \u_outFIFO/U1501  ( .A(\u_outFIFO/FIFO[108][3] ), .B(
        \u_outFIFO/FIFO[109][3] ), .C(\u_outFIFO/FIFO[110][3] ), .D(
        \u_outFIFO/FIFO[111][3] ), .S0(n1180), .S1(\u_outFIFO/N40 ), .Q(
        \u_outFIFO/n1529 ) );
  IMUX40 \u_outFIFO/U1509  ( .A(\u_outFIFO/FIFO[76][3] ), .B(
        \u_outFIFO/FIFO[77][3] ), .C(\u_outFIFO/FIFO[78][3] ), .D(
        \u_outFIFO/FIFO[79][3] ), .S0(n1177), .S1(\u_outFIFO/N40 ), .Q(
        \u_outFIFO/n1539 ) );
  IMUX40 \u_outFIFO/U1500  ( .A(\u_outFIFO/FIFO[112][3] ), .B(
        \u_outFIFO/FIFO[113][3] ), .C(\u_outFIFO/FIFO[114][3] ), .D(
        \u_outFIFO/FIFO[115][3] ), .S0(n1180), .S1(\u_outFIFO/N40 ), .Q(
        \u_outFIFO/n1521 ) );
  IMUX40 \u_outFIFO/U1529  ( .A(\u_outFIFO/FIFO[0][3] ), .B(
        \u_outFIFO/FIFO[1][3] ), .C(\u_outFIFO/FIFO[2][3] ), .D(
        \u_outFIFO/FIFO[3][3] ), .S0(n1176), .S1(n1182), .Q(\u_outFIFO/n1556 )
         );
  IMUX40 \u_outFIFO/U1527  ( .A(\u_outFIFO/FIFO[8][3] ), .B(
        \u_outFIFO/FIFO[9][3] ), .C(\u_outFIFO/FIFO[10][3] ), .D(
        \u_outFIFO/FIFO[11][3] ), .S0(n1176), .S1(n1182), .Q(\u_outFIFO/n1557 ) );
  IMUX40 \u_outFIFO/U1528  ( .A(\u_outFIFO/FIFO[4][3] ), .B(
        \u_outFIFO/FIFO[5][3] ), .C(\u_outFIFO/FIFO[6][3] ), .D(
        \u_outFIFO/FIFO[7][3] ), .S0(n1176), .S1(n1182), .Q(\u_outFIFO/n1558 )
         );
  IMUX40 \u_outFIFO/U1393  ( .A(\u_outFIFO/n1556 ), .B(\u_outFIFO/n1557 ), .C(
        \u_outFIFO/n1558 ), .D(\u_outFIFO/n1559 ), .S0(\u_outFIFO/N42 ), .S1(
        n14), .Q(\u_outFIFO/n1555 ) );
  IMUX40 \u_outFIFO/U1400  ( .A(\u_outFIFO/FIFO[104][0] ), .B(
        \u_outFIFO/FIFO[105][0] ), .C(\u_outFIFO/FIFO[106][0] ), .D(
        \u_outFIFO/FIFO[107][0] ), .S0(n1180), .S1(n1182), .Q(
        \u_outFIFO/n1401 ) );
  IMUX40 \u_outFIFO/U1399  ( .A(\u_outFIFO/FIFO[108][0] ), .B(
        \u_outFIFO/FIFO[109][0] ), .C(\u_outFIFO/FIFO[110][0] ), .D(
        \u_outFIFO/FIFO[111][0] ), .S0(n1180), .S1(n1181), .Q(
        \u_outFIFO/n1403 ) );
  IMUX40 \u_outFIFO/U1401  ( .A(\u_outFIFO/FIFO[100][0] ), .B(
        \u_outFIFO/FIFO[101][0] ), .C(\u_outFIFO/FIFO[102][0] ), .D(
        \u_outFIFO/FIFO[103][0] ), .S0(n1180), .S1(n1181), .Q(
        \u_outFIFO/n1402 ) );
  IMUX40 \u_outFIFO/U1360  ( .A(\u_outFIFO/n1400 ), .B(\u_outFIFO/n1401 ), .C(
        \u_outFIFO/n1402 ), .D(\u_outFIFO/n1403 ), .S0(n1183), .S1(n14), .Q(
        \u_outFIFO/n1399 ) );
  IMUX40 \u_outFIFO/U1396  ( .A(\u_outFIFO/FIFO[120][0] ), .B(
        \u_outFIFO/FIFO[121][0] ), .C(\u_outFIFO/FIFO[122][0] ), .D(
        \u_outFIFO/FIFO[123][0] ), .S0(n1180), .S1(n1181), .Q(
        \u_outFIFO/n1396 ) );
  IMUX40 \u_outFIFO/U1395  ( .A(\u_outFIFO/FIFO[124][0] ), .B(
        \u_outFIFO/FIFO[125][0] ), .C(\u_outFIFO/FIFO[126][0] ), .D(
        \u_outFIFO/FIFO[127][0] ), .S0(n1180), .S1(\u_outFIFO/N40 ), .Q(
        \u_outFIFO/n1398 ) );
  IMUX40 \u_outFIFO/U1397  ( .A(\u_outFIFO/FIFO[116][0] ), .B(
        \u_outFIFO/FIFO[117][0] ), .C(\u_outFIFO/FIFO[118][0] ), .D(
        \u_outFIFO/FIFO[119][0] ), .S0(n1180), .S1(\u_outFIFO/N40 ), .Q(
        \u_outFIFO/n1397 ) );
  IMUX40 \u_outFIFO/U1359  ( .A(\u_outFIFO/n1395 ), .B(\u_outFIFO/n1396 ), .C(
        \u_outFIFO/n1397 ), .D(\u_outFIFO/n1398 ), .S0(n1183), .S1(n14), .Q(
        \u_outFIFO/n1394 ) );
  IMUX40 \u_outFIFO/U1410  ( .A(\u_outFIFO/FIFO[64][0] ), .B(
        \u_outFIFO/FIFO[65][0] ), .C(\u_outFIFO/FIFO[66][0] ), .D(
        \u_outFIFO/FIFO[67][0] ), .S0(n759), .S1(n1182), .Q(\u_outFIFO/n1410 )
         );
  IMUX40 \u_outFIFO/U1408  ( .A(\u_outFIFO/FIFO[72][0] ), .B(
        \u_outFIFO/FIFO[73][0] ), .C(\u_outFIFO/FIFO[74][0] ), .D(
        \u_outFIFO/FIFO[75][0] ), .S0(\u_outFIFO/N39 ), .S1(\u_outFIFO/N40 ), 
        .Q(\u_outFIFO/n1411 ) );
  IMUX40 \u_outFIFO/U1409  ( .A(\u_outFIFO/FIFO[68][0] ), .B(
        \u_outFIFO/FIFO[69][0] ), .C(\u_outFIFO/FIFO[70][0] ), .D(
        \u_outFIFO/FIFO[71][0] ), .S0(\u_outFIFO/N39 ), .S1(\u_outFIFO/N40 ), 
        .Q(\u_outFIFO/n1412 ) );
  IMUX40 \u_outFIFO/U1362  ( .A(\u_outFIFO/n1410 ), .B(\u_outFIFO/n1411 ), .C(
        \u_outFIFO/n1412 ), .D(\u_outFIFO/n1413 ), .S0(n1183), .S1(n14), .Q(
        \u_outFIFO/n1409 ) );
  IMUX40 \u_outFIFO/U1427  ( .A(\u_outFIFO/FIFO[0][0] ), .B(
        \u_outFIFO/FIFO[1][0] ), .C(\u_outFIFO/FIFO[2][0] ), .D(
        \u_outFIFO/FIFO[3][0] ), .S0(n1179), .S1(n1182), .Q(\u_outFIFO/n1430 )
         );
  IMUX40 \u_outFIFO/U1425  ( .A(\u_outFIFO/FIFO[8][0] ), .B(
        \u_outFIFO/FIFO[9][0] ), .C(\u_outFIFO/FIFO[10][0] ), .D(
        \u_outFIFO/FIFO[11][0] ), .S0(n1179), .S1(\u_outFIFO/N40 ), .Q(
        \u_outFIFO/n1431 ) );
  IMUX40 \u_outFIFO/U1426  ( .A(\u_outFIFO/FIFO[4][0] ), .B(
        \u_outFIFO/FIFO[5][0] ), .C(\u_outFIFO/FIFO[6][0] ), .D(
        \u_outFIFO/FIFO[7][0] ), .S0(n1179), .S1(n1182), .Q(\u_outFIFO/n1432 )
         );
  IMUX40 \u_outFIFO/U1366  ( .A(\u_outFIFO/n1430 ), .B(\u_outFIFO/n1431 ), .C(
        \u_outFIFO/n1432 ), .D(\u_outFIFO/n1433 ), .S0(n1183), .S1(n14), .Q(
        \u_outFIFO/n1429 ) );
  IMUX40 \u_outFIFO/U1436  ( .A(\u_outFIFO/FIFO[96][1] ), .B(
        \u_outFIFO/FIFO[97][1] ), .C(\u_outFIFO/FIFO[98][1] ), .D(
        \u_outFIFO/FIFO[99][1] ), .S0(n1178), .S1(n1182), .Q(\u_outFIFO/n1442 ) );
  IMUX40 \u_outFIFO/U1434  ( .A(\u_outFIFO/FIFO[104][1] ), .B(
        \u_outFIFO/FIFO[105][1] ), .C(\u_outFIFO/FIFO[106][1] ), .D(
        \u_outFIFO/FIFO[107][1] ), .S0(n1178), .S1(n1182), .Q(
        \u_outFIFO/n1443 ) );
  IMUX40 \u_outFIFO/U1435  ( .A(\u_outFIFO/FIFO[100][1] ), .B(
        \u_outFIFO/FIFO[101][1] ), .C(\u_outFIFO/FIFO[102][1] ), .D(
        \u_outFIFO/FIFO[103][1] ), .S0(n1178), .S1(n1182), .Q(
        \u_outFIFO/n1444 ) );
  IMUX40 \u_outFIFO/U1369  ( .A(\u_outFIFO/n1442 ), .B(\u_outFIFO/n1443 ), .C(
        \u_outFIFO/n1444 ), .D(\u_outFIFO/n1445 ), .S0(\u_outFIFO/N42 ), .S1(
        n14), .Q(\u_outFIFO/n1441 ) );
  IMUX40 \u_outFIFO/U1444  ( .A(\u_outFIFO/FIFO[64][1] ), .B(
        \u_outFIFO/FIFO[65][1] ), .C(\u_outFIFO/FIFO[66][1] ), .D(
        \u_outFIFO/FIFO[67][1] ), .S0(\u_outFIFO/N39 ), .S1(\u_outFIFO/N40 ), 
        .Q(\u_outFIFO/n1452 ) );
  IMUX40 \u_outFIFO/U1442  ( .A(\u_outFIFO/FIFO[72][1] ), .B(
        \u_outFIFO/FIFO[73][1] ), .C(\u_outFIFO/FIFO[74][1] ), .D(
        \u_outFIFO/FIFO[75][1] ), .S0(\u_outFIFO/N39 ), .S1(\u_outFIFO/N40 ), 
        .Q(\u_outFIFO/n1453 ) );
  IMUX40 \u_outFIFO/U1443  ( .A(\u_outFIFO/FIFO[68][1] ), .B(
        \u_outFIFO/FIFO[69][1] ), .C(\u_outFIFO/FIFO[70][1] ), .D(
        \u_outFIFO/FIFO[71][1] ), .S0(\u_outFIFO/N39 ), .S1(\u_outFIFO/N40 ), 
        .Q(\u_outFIFO/n1454 ) );
  IMUX40 \u_outFIFO/U1371  ( .A(\u_outFIFO/n1452 ), .B(\u_outFIFO/n1453 ), .C(
        \u_outFIFO/n1454 ), .D(\u_outFIFO/n1455 ), .S0(\u_outFIFO/N42 ), .S1(
        n14), .Q(\u_outFIFO/n1451 ) );
  IMUX40 \u_outFIFO/U1430  ( .A(\u_outFIFO/FIFO[120][1] ), .B(
        \u_outFIFO/FIFO[121][1] ), .C(\u_outFIFO/FIFO[122][1] ), .D(
        \u_outFIFO/FIFO[123][1] ), .S0(n1178), .S1(n1182), .Q(
        \u_outFIFO/n1438 ) );
  IMUX40 \u_outFIFO/U1429  ( .A(\u_outFIFO/FIFO[124][1] ), .B(
        \u_outFIFO/FIFO[125][1] ), .C(\u_outFIFO/FIFO[126][1] ), .D(
        \u_outFIFO/FIFO[127][1] ), .S0(n1178), .S1(n1182), .Q(
        \u_outFIFO/n1440 ) );
  IMUX40 \u_outFIFO/U1431  ( .A(\u_outFIFO/FIFO[116][1] ), .B(
        \u_outFIFO/FIFO[117][1] ), .C(\u_outFIFO/FIFO[118][1] ), .D(
        \u_outFIFO/FIFO[119][1] ), .S0(n1178), .S1(n1182), .Q(
        \u_outFIFO/n1439 ) );
  IMUX40 \u_outFIFO/U1368  ( .A(\u_outFIFO/n1437 ), .B(\u_outFIFO/n1438 ), .C(
        \u_outFIFO/n1439 ), .D(\u_outFIFO/n1440 ), .S0(n1183), .S1(n14), .Q(
        \u_outFIFO/n1436 ) );
  IMUX40 \u_outFIFO/U1461  ( .A(\u_outFIFO/FIFO[0][1] ), .B(
        \u_outFIFO/FIFO[1][1] ), .C(\u_outFIFO/FIFO[2][1] ), .D(
        \u_outFIFO/FIFO[3][1] ), .S0(n1177), .S1(n1182), .Q(\u_outFIFO/n1472 )
         );
  IMUX40 \u_outFIFO/U1459  ( .A(\u_outFIFO/FIFO[8][1] ), .B(
        \u_outFIFO/FIFO[9][1] ), .C(\u_outFIFO/FIFO[10][1] ), .D(
        \u_outFIFO/FIFO[11][1] ), .S0(n1177), .S1(\u_outFIFO/N40 ), .Q(
        \u_outFIFO/n1473 ) );
  IMUX40 \u_outFIFO/U1460  ( .A(\u_outFIFO/FIFO[4][1] ), .B(
        \u_outFIFO/FIFO[5][1] ), .C(\u_outFIFO/FIFO[6][1] ), .D(
        \u_outFIFO/FIFO[7][1] ), .S0(n1177), .S1(n760), .Q(\u_outFIFO/n1474 )
         );
  IMUX40 \u_outFIFO/U1375  ( .A(\u_outFIFO/n1472 ), .B(\u_outFIFO/n1473 ), .C(
        \u_outFIFO/n1474 ), .D(\u_outFIFO/n1475 ), .S0(\u_outFIFO/N42 ), .S1(
        n14), .Q(\u_outFIFO/n1471 ) );
  IMUX40 \u_outFIFO/U1470  ( .A(\u_outFIFO/FIFO[96][2] ), .B(
        \u_outFIFO/FIFO[97][2] ), .C(\u_outFIFO/FIFO[98][2] ), .D(
        \u_outFIFO/FIFO[99][2] ), .S0(n759), .S1(n1181), .Q(\u_outFIFO/n1484 )
         );
  IMUX40 \u_outFIFO/U1468  ( .A(\u_outFIFO/FIFO[104][2] ), .B(
        \u_outFIFO/FIFO[105][2] ), .C(\u_outFIFO/FIFO[106][2] ), .D(
        \u_outFIFO/FIFO[107][2] ), .S0(n1177), .S1(n1181), .Q(
        \u_outFIFO/n1485 ) );
  IMUX40 \u_outFIFO/U1469  ( .A(\u_outFIFO/FIFO[100][2] ), .B(
        \u_outFIFO/FIFO[101][2] ), .C(\u_outFIFO/FIFO[102][2] ), .D(
        \u_outFIFO/FIFO[103][2] ), .S0(n1179), .S1(n1181), .Q(
        \u_outFIFO/n1486 ) );
  IMUX40 \u_outFIFO/U1378  ( .A(\u_outFIFO/n1484 ), .B(\u_outFIFO/n1485 ), .C(
        \u_outFIFO/n1486 ), .D(\u_outFIFO/n1487 ), .S0(\u_outFIFO/N42 ), .S1(
        n14), .Q(\u_outFIFO/n1483 ) );
  IMUX40 \u_outFIFO/U1478  ( .A(\u_outFIFO/FIFO[64][2] ), .B(
        \u_outFIFO/FIFO[65][2] ), .C(\u_outFIFO/FIFO[66][2] ), .D(
        \u_outFIFO/FIFO[67][2] ), .S0(n759), .S1(n1181), .Q(\u_outFIFO/n1494 )
         );
  IMUX40 \u_outFIFO/U1476  ( .A(\u_outFIFO/FIFO[72][2] ), .B(
        \u_outFIFO/FIFO[73][2] ), .C(\u_outFIFO/FIFO[74][2] ), .D(
        \u_outFIFO/FIFO[75][2] ), .S0(n759), .S1(n1181), .Q(\u_outFIFO/n1495 )
         );
  IMUX40 \u_outFIFO/U1477  ( .A(\u_outFIFO/FIFO[68][2] ), .B(
        \u_outFIFO/FIFO[69][2] ), .C(\u_outFIFO/FIFO[70][2] ), .D(
        \u_outFIFO/FIFO[71][2] ), .S0(n759), .S1(n1181), .Q(\u_outFIFO/n1496 )
         );
  IMUX40 \u_outFIFO/U1380  ( .A(\u_outFIFO/n1494 ), .B(\u_outFIFO/n1495 ), .C(
        \u_outFIFO/n1496 ), .D(\u_outFIFO/n1497 ), .S0(\u_outFIFO/N42 ), .S1(
        n14), .Q(\u_outFIFO/n1493 ) );
  IMUX40 \u_outFIFO/U1464  ( .A(\u_outFIFO/FIFO[120][2] ), .B(
        \u_outFIFO/FIFO[121][2] ), .C(\u_outFIFO/FIFO[122][2] ), .D(
        \u_outFIFO/FIFO[123][2] ), .S0(n1177), .S1(n1182), .Q(
        \u_outFIFO/n1480 ) );
  IMUX40 \u_outFIFO/U1463  ( .A(\u_outFIFO/FIFO[124][2] ), .B(
        \u_outFIFO/FIFO[125][2] ), .C(\u_outFIFO/FIFO[126][2] ), .D(
        \u_outFIFO/FIFO[127][2] ), .S0(n1177), .S1(\u_outFIFO/N40 ), .Q(
        \u_outFIFO/n1482 ) );
  IMUX40 \u_outFIFO/U1465  ( .A(\u_outFIFO/FIFO[116][2] ), .B(
        \u_outFIFO/FIFO[117][2] ), .C(\u_outFIFO/FIFO[118][2] ), .D(
        \u_outFIFO/FIFO[119][2] ), .S0(n1177), .S1(n1181), .Q(
        \u_outFIFO/n1481 ) );
  IMUX40 \u_outFIFO/U1377  ( .A(\u_outFIFO/n1479 ), .B(\u_outFIFO/n1480 ), .C(
        \u_outFIFO/n1481 ), .D(\u_outFIFO/n1482 ), .S0(n1183), .S1(n14), .Q(
        \u_outFIFO/n1478 ) );
  IMUX40 \u_outFIFO/U1495  ( .A(\u_outFIFO/FIFO[0][2] ), .B(
        \u_outFIFO/FIFO[1][2] ), .C(\u_outFIFO/FIFO[2][2] ), .D(
        \u_outFIFO/FIFO[3][2] ), .S0(\u_outFIFO/N39 ), .S1(n760), .Q(
        \u_outFIFO/n1514 ) );
  IMUX40 \u_outFIFO/U1493  ( .A(\u_outFIFO/FIFO[8][2] ), .B(
        \u_outFIFO/FIFO[9][2] ), .C(\u_outFIFO/FIFO[10][2] ), .D(
        \u_outFIFO/FIFO[11][2] ), .S0(\u_outFIFO/N39 ), .S1(n760), .Q(
        \u_outFIFO/n1515 ) );
  IMUX40 \u_outFIFO/U1494  ( .A(\u_outFIFO/FIFO[4][2] ), .B(
        \u_outFIFO/FIFO[5][2] ), .C(\u_outFIFO/FIFO[6][2] ), .D(
        \u_outFIFO/FIFO[7][2] ), .S0(\u_outFIFO/N39 ), .S1(n760), .Q(
        \u_outFIFO/n1516 ) );
  IMUX40 \u_outFIFO/U1384  ( .A(\u_outFIFO/n1514 ), .B(\u_outFIFO/n1515 ), .C(
        \u_outFIFO/n1516 ), .D(\u_outFIFO/n1517 ), .S0(\u_outFIFO/N42 ), .S1(
        n14), .Q(\u_outFIFO/n1513 ) );
  IMUX40 \u_outFIFO/U1504  ( .A(\u_outFIFO/FIFO[96][3] ), .B(
        \u_outFIFO/FIFO[97][3] ), .C(\u_outFIFO/FIFO[98][3] ), .D(
        \u_outFIFO/FIFO[99][3] ), .S0(\u_outFIFO/N39 ), .S1(\u_outFIFO/N40 ), 
        .Q(\u_outFIFO/n1526 ) );
  IMUX40 \u_outFIFO/U1502  ( .A(\u_outFIFO/FIFO[104][3] ), .B(
        \u_outFIFO/FIFO[105][3] ), .C(\u_outFIFO/FIFO[106][3] ), .D(
        \u_outFIFO/FIFO[107][3] ), .S0(\u_outFIFO/N39 ), .S1(\u_outFIFO/N40 ), 
        .Q(\u_outFIFO/n1527 ) );
  IMUX40 \u_outFIFO/U1503  ( .A(\u_outFIFO/FIFO[100][3] ), .B(
        \u_outFIFO/FIFO[101][3] ), .C(\u_outFIFO/FIFO[102][3] ), .D(
        \u_outFIFO/FIFO[103][3] ), .S0(\u_outFIFO/N39 ), .S1(\u_outFIFO/N40 ), 
        .Q(\u_outFIFO/n1528 ) );
  IMUX40 \u_outFIFO/U1387  ( .A(\u_outFIFO/n1526 ), .B(\u_outFIFO/n1527 ), .C(
        \u_outFIFO/n1528 ), .D(\u_outFIFO/n1529 ), .S0(\u_outFIFO/N42 ), .S1(
        n14), .Q(\u_outFIFO/n1525 ) );
  IMUX40 \u_outFIFO/U1512  ( .A(\u_outFIFO/FIFO[64][3] ), .B(
        \u_outFIFO/FIFO[65][3] ), .C(\u_outFIFO/FIFO[66][3] ), .D(
        \u_outFIFO/FIFO[67][3] ), .S0(n1178), .S1(n760), .Q(\u_outFIFO/n1536 )
         );
  IMUX40 \u_outFIFO/U1510  ( .A(\u_outFIFO/FIFO[72][3] ), .B(
        \u_outFIFO/FIFO[73][3] ), .C(\u_outFIFO/FIFO[74][3] ), .D(
        \u_outFIFO/FIFO[75][3] ), .S0(\u_outFIFO/N39 ), .S1(\u_outFIFO/N40 ), 
        .Q(\u_outFIFO/n1537 ) );
  IMUX40 \u_outFIFO/U1511  ( .A(\u_outFIFO/FIFO[68][3] ), .B(
        \u_outFIFO/FIFO[69][3] ), .C(\u_outFIFO/FIFO[70][3] ), .D(
        \u_outFIFO/FIFO[71][3] ), .S0(n759), .S1(n1182), .Q(\u_outFIFO/n1538 )
         );
  IMUX40 \u_outFIFO/U1389  ( .A(\u_outFIFO/n1536 ), .B(\u_outFIFO/n1537 ), .C(
        \u_outFIFO/n1538 ), .D(\u_outFIFO/n1539 ), .S0(\u_outFIFO/N42 ), .S1(
        n14), .Q(\u_outFIFO/n1535 ) );
  IMUX40 \u_outFIFO/U1498  ( .A(\u_outFIFO/FIFO[120][3] ), .B(
        \u_outFIFO/FIFO[121][3] ), .C(\u_outFIFO/FIFO[122][3] ), .D(
        \u_outFIFO/FIFO[123][3] ), .S0(\u_outFIFO/N39 ), .S1(\u_outFIFO/N40 ), 
        .Q(\u_outFIFO/n1522 ) );
  IMUX40 \u_outFIFO/U1497  ( .A(\u_outFIFO/FIFO[124][3] ), .B(
        \u_outFIFO/FIFO[125][3] ), .C(\u_outFIFO/FIFO[126][3] ), .D(
        \u_outFIFO/FIFO[127][3] ), .S0(\u_outFIFO/N39 ), .S1(\u_outFIFO/N40 ), 
        .Q(\u_outFIFO/n1524 ) );
  IMUX40 \u_outFIFO/U1499  ( .A(\u_outFIFO/FIFO[116][3] ), .B(
        \u_outFIFO/FIFO[117][3] ), .C(\u_outFIFO/FIFO[118][3] ), .D(
        \u_outFIFO/FIFO[119][3] ), .S0(\u_outFIFO/N39 ), .S1(\u_outFIFO/N40 ), 
        .Q(\u_outFIFO/n1523 ) );
  IMUX40 \u_outFIFO/U1386  ( .A(\u_outFIFO/n1521 ), .B(\u_outFIFO/n1522 ), .C(
        \u_outFIFO/n1523 ), .D(\u_outFIFO/n1524 ), .S0(\u_outFIFO/N42 ), .S1(
        n14), .Q(\u_outFIFO/n1520 ) );
  IMUX40 \u_outFIFO/U1364  ( .A(\u_outFIFO/n1420 ), .B(\u_outFIFO/n1421 ), .C(
        \u_outFIFO/n1422 ), .D(\u_outFIFO/n1423 ), .S0(n1183), .S1(n14), .Q(
        \u_outFIFO/n1419 ) );
  IMUX40 \u_outFIFO/U1363  ( .A(\u_outFIFO/n1415 ), .B(\u_outFIFO/n1416 ), .C(
        \u_outFIFO/n1417 ), .D(\u_outFIFO/n1418 ), .S0(n1183), .S1(n14), .Q(
        \u_outFIFO/n1414 ) );
  IMUX40 \u_outFIFO/U1365  ( .A(\u_outFIFO/n1425 ), .B(\u_outFIFO/n1426 ), .C(
        \u_outFIFO/n1427 ), .D(\u_outFIFO/n1428 ), .S0(n1183), .S1(n14), .Q(
        \u_outFIFO/n1424 ) );
  IMUX40 \u_outFIFO/U1428  ( .A(\u_outFIFO/n1429 ), .B(\u_outFIFO/n1419 ), .C(
        \u_outFIFO/n1424 ), .D(\u_outFIFO/n1414 ), .S0(n761), .S1(
        \u_outFIFO/N43 ), .Q(\u_outFIFO/n1434 ) );
  IMUX40 \u_outFIFO/U1373  ( .A(\u_outFIFO/n1462 ), .B(\u_outFIFO/n1463 ), .C(
        \u_outFIFO/n1464 ), .D(\u_outFIFO/n1465 ), .S0(\u_outFIFO/N42 ), .S1(
        n14), .Q(\u_outFIFO/n1461 ) );
  IMUX40 \u_outFIFO/U1372  ( .A(\u_outFIFO/n1457 ), .B(\u_outFIFO/n1458 ), .C(
        \u_outFIFO/n1459 ), .D(\u_outFIFO/n1460 ), .S0(n1183), .S1(n14), .Q(
        \u_outFIFO/n1456 ) );
  IMUX40 \u_outFIFO/U1374  ( .A(\u_outFIFO/n1467 ), .B(\u_outFIFO/n1468 ), .C(
        \u_outFIFO/n1469 ), .D(\u_outFIFO/n1470 ), .S0(\u_outFIFO/N42 ), .S1(
        n14), .Q(\u_outFIFO/n1466 ) );
  IMUX40 \u_outFIFO/U1462  ( .A(\u_outFIFO/n1471 ), .B(\u_outFIFO/n1461 ), .C(
        \u_outFIFO/n1466 ), .D(\u_outFIFO/n1456 ), .S0(n761), .S1(
        \u_outFIFO/N43 ), .Q(\u_outFIFO/n1476 ) );
  IMUX40 \u_outFIFO/U1382  ( .A(\u_outFIFO/n1504 ), .B(\u_outFIFO/n1505 ), .C(
        \u_outFIFO/n1506 ), .D(\u_outFIFO/n1507 ), .S0(\u_outFIFO/N42 ), .S1(
        n14), .Q(\u_outFIFO/n1503 ) );
  IMUX40 \u_outFIFO/U1381  ( .A(\u_outFIFO/n1499 ), .B(\u_outFIFO/n1500 ), .C(
        \u_outFIFO/n1501 ), .D(\u_outFIFO/n1502 ), .S0(\u_outFIFO/N42 ), .S1(
        n14), .Q(\u_outFIFO/n1498 ) );
  IMUX40 \u_outFIFO/U1383  ( .A(\u_outFIFO/n1509 ), .B(\u_outFIFO/n1510 ), .C(
        \u_outFIFO/n1511 ), .D(\u_outFIFO/n1512 ), .S0(\u_outFIFO/N42 ), .S1(
        n14), .Q(\u_outFIFO/n1508 ) );
  IMUX40 \u_outFIFO/U1496  ( .A(\u_outFIFO/n1513 ), .B(\u_outFIFO/n1503 ), .C(
        \u_outFIFO/n1508 ), .D(\u_outFIFO/n1498 ), .S0(n761), .S1(
        \u_outFIFO/N43 ), .Q(\u_outFIFO/n1518 ) );
  IMUX40 \u_outFIFO/U1391  ( .A(\u_outFIFO/n1546 ), .B(\u_outFIFO/n1547 ), .C(
        \u_outFIFO/n1548 ), .D(\u_outFIFO/n1549 ), .S0(\u_outFIFO/N42 ), .S1(
        n14), .Q(\u_outFIFO/n1545 ) );
  IMUX40 \u_outFIFO/U1390  ( .A(\u_outFIFO/n1541 ), .B(\u_outFIFO/n1542 ), .C(
        \u_outFIFO/n1543 ), .D(\u_outFIFO/n1544 ), .S0(\u_outFIFO/N42 ), .S1(
        n14), .Q(\u_outFIFO/n1540 ) );
  IMUX40 \u_outFIFO/U1392  ( .A(\u_outFIFO/n1551 ), .B(\u_outFIFO/n1552 ), .C(
        \u_outFIFO/n1553 ), .D(\u_outFIFO/n1554 ), .S0(\u_outFIFO/N42 ), .S1(
        n14), .Q(\u_outFIFO/n1550 ) );
  IMUX40 \u_outFIFO/U1530  ( .A(\u_outFIFO/n1555 ), .B(\u_outFIFO/n1545 ), .C(
        \u_outFIFO/n1550 ), .D(\u_outFIFO/n1540 ), .S0(n761), .S1(
        \u_outFIFO/N43 ), .Q(\u_outFIFO/n1560 ) );
  XOR31 \u_cordic/mycordic/sub_182/U2_7  ( .A(
        \u_cordic/mycordic/present_I_table[1][7] ), .B(n304), .C(
        \u_cordic/mycordic/sub_182/carry [7]), .Q(\u_cordic/mycordic/N291 ) );
  IMUX21 \u_cordic/mycordic/U539  ( .A(\u_cordic/mycordic/n572 ), .B(n380), 
        .S(n766), .Q(\u_cordic/mycordic/n571 ) );
  MUX22 \u_cordic/mycordic/U540  ( .A(
        \u_cordic/mycordic/present_ANGLE_table[6][8] ), .B(
        \u_cordic/mycordic/n571 ), .S(n384), .Q(
        \u_cordic/mycordic/next_ANGLE_table[6][8] ) );
  IMUX21 \u_cordic/mycordic/U547  ( .A(\u_cordic/mycordic/n580 ), .B(n382), 
        .S(n766), .Q(\u_cordic/mycordic/n579 ) );
  MUX22 \u_cordic/mycordic/U548  ( .A(
        \u_cordic/mycordic/present_ANGLE_table[6][12] ), .B(
        \u_cordic/mycordic/n579 ), .S(n384), .Q(
        \u_cordic/mycordic/next_ANGLE_table[6][12] ) );
  IMUX21 \u_cordic/mycordic/U545  ( .A(\u_cordic/mycordic/n578 ), .B(n378), 
        .S(n766), .Q(\u_cordic/mycordic/n577 ) );
  MUX22 \u_cordic/mycordic/U546  ( .A(
        \u_cordic/mycordic/present_ANGLE_table[6][11] ), .B(
        \u_cordic/mycordic/n577 ), .S(n384), .Q(
        \u_cordic/mycordic/next_ANGLE_table[6][11] ) );
  IMUX21 \u_cordic/mycordic/U541  ( .A(\u_cordic/mycordic/n574 ), .B(n381), 
        .S(n766), .Q(\u_cordic/mycordic/n573 ) );
  MUX22 \u_cordic/mycordic/U542  ( .A(
        \u_cordic/mycordic/present_ANGLE_table[6][9] ), .B(
        \u_cordic/mycordic/n573 ), .S(n384), .Q(
        \u_cordic/mycordic/next_ANGLE_table[6][9] ) );
  NAND22 \u_cordic/mycordic/U569  ( .A(\u_cordic/mycordic/N627 ), .B(n758), 
        .Q(\u_cordic/mycordic/n580 ) );
  NAND22 \u_cordic/mycordic/U566  ( .A(\u_cordic/mycordic/N624 ), .B(n757), 
        .Q(\u_cordic/mycordic/n574 ) );
  IMUX40 \u_inFIFO/U568  ( .A(\u_inFIFO/n637 ), .B(\u_inFIFO/n638 ), .C(
        \u_inFIFO/n639 ), .D(\u_inFIFO/n640 ), .S0(\u_inFIFO/N40 ), .S1(n15), 
        .Q(\u_inFIFO/n636 ) );
  IMUX40 \u_inFIFO/U660  ( .A(\u_inFIFO/n661 ), .B(\u_inFIFO/n651 ), .C(
        \u_inFIFO/n656 ), .D(\u_inFIFO/n646 ), .S0(n49), .S1(n765), .Q(
        \u_inFIFO/n666 ) );
  IMUX40 \u_inFIFO/U643  ( .A(\u_inFIFO/n641 ), .B(\u_inFIFO/n631 ), .C(
        \u_inFIFO/n636 ), .D(\u_inFIFO/n626 ), .S0(n49), .S1(n765), .Q(
        \u_inFIFO/n667 ) );
  IMUX21 \u_inFIFO/U574  ( .A(\u_inFIFO/n666 ), .B(\u_inFIFO/n667 ), .S(
        \u_inFIFO/N43 ), .Q(\u_inFIFO/N202 ) );
  IMUX40 \u_inFIFO/U577  ( .A(\u_inFIFO/n679 ), .B(\u_inFIFO/n680 ), .C(
        \u_inFIFO/n681 ), .D(\u_inFIFO/n682 ), .S0(\u_inFIFO/N40 ), .S1(n15), 
        .Q(\u_inFIFO/n678 ) );
  IMUX40 \u_inFIFO/U694  ( .A(\u_inFIFO/n703 ), .B(\u_inFIFO/n693 ), .C(
        \u_inFIFO/n698 ), .D(\u_inFIFO/n688 ), .S0(n49), .S1(n765), .Q(
        \u_inFIFO/n708 ) );
  IMUX40 \u_inFIFO/U677  ( .A(\u_inFIFO/n683 ), .B(\u_inFIFO/n673 ), .C(
        \u_inFIFO/n678 ), .D(\u_inFIFO/n668 ), .S0(n49), .S1(n765), .Q(
        \u_inFIFO/n709 ) );
  IMUX21 \u_inFIFO/U583  ( .A(\u_inFIFO/n708 ), .B(\u_inFIFO/n709 ), .S(
        \u_inFIFO/N43 ), .Q(\u_inFIFO/N201 ) );
  IMUX40 \u_inFIFO/U558  ( .A(\u_inFIFO/n590 ), .B(\u_inFIFO/n591 ), .C(
        \u_inFIFO/n592 ), .D(\u_inFIFO/n593 ), .S0(n1202), .S1(n15), .Q(
        \u_inFIFO/n589 ) );
  IMUX40 \u_inFIFO/U626  ( .A(\u_inFIFO/n619 ), .B(\u_inFIFO/n609 ), .C(
        \u_inFIFO/n614 ), .D(\u_inFIFO/n604 ), .S0(n49), .S1(n765), .Q(
        \u_inFIFO/n624 ) );
  IMUX40 \u_inFIFO/U609  ( .A(\u_inFIFO/n599 ), .B(\u_inFIFO/n589 ), .C(
        \u_inFIFO/n594 ), .D(\u_inFIFO/n584 ), .S0(n49), .S1(n765), .Q(
        \u_inFIFO/n625 ) );
  IMUX21 \u_inFIFO/U565  ( .A(\u_inFIFO/n624 ), .B(\u_inFIFO/n625 ), .S(
        \u_inFIFO/N43 ), .Q(\u_inFIFO/N203 ) );
  IMUX21 \u_cordic/mycordic/U543  ( .A(\u_cordic/mycordic/n576 ), .B(n377), 
        .S(n766), .Q(\u_cordic/mycordic/n575 ) );
  MUX22 \u_cordic/mycordic/U544  ( .A(
        \u_cordic/mycordic/present_ANGLE_table[6][10] ), .B(
        \u_cordic/mycordic/n575 ), .S(n384), .Q(
        \u_cordic/mycordic/next_ANGLE_table[6][10] ) );
  NAND22 \u_cordic/mycordic/U570  ( .A(\u_cordic/mycordic/N628 ), .B(n757), 
        .Q(\u_cordic/mycordic/n582 ) );
  NAND22 \u_cordic/mycordic/U568  ( .A(\u_cordic/mycordic/N626 ), .B(n757), 
        .Q(\u_cordic/mycordic/n578 ) );
  NAND22 \u_cordic/mycordic/U567  ( .A(\u_cordic/mycordic/N625 ), .B(n758), 
        .Q(\u_cordic/mycordic/n576 ) );
  XOR31 \u_cordic/mycordic/sub_178/U2_7  ( .A(
        \u_cordic/mycordic/present_Q_table[1][7] ), .B(n307), .C(
        \u_cordic/mycordic/sub_178/carry [7]), .Q(\u_cordic/mycordic/N267 ) );
  IMUX40 \u_inFIFO/U599  ( .A(\u_inFIFO/FIFO[100][0] ), .B(
        \u_inFIFO/FIFO[101][0] ), .C(\u_inFIFO/FIFO[102][0] ), .D(
        \u_inFIFO/FIFO[103][0] ), .S0(n1196), .S1(n1201), .Q(\u_inFIFO/n592 )
         );
  IMUX40 \u_inFIFO/U722  ( .A(\u_inFIFO/FIFO[20][3] ), .B(
        \u_inFIFO/FIFO[21][3] ), .C(\u_inFIFO/FIFO[22][3] ), .D(
        \u_inFIFO/FIFO[23][3] ), .S0(n13), .S1(\u_inFIFO/N38 ), .Q(
        \u_inFIFO/n743 ) );
  IMUX40 \u_inFIFO/U714  ( .A(\u_inFIFO/FIFO[52][3] ), .B(
        \u_inFIFO/FIFO[53][3] ), .C(\u_inFIFO/FIFO[54][3] ), .D(
        \u_inFIFO/FIFO[55][3] ), .S0(n13), .S1(n764), .Q(\u_inFIFO/n733 ) );
  IMUX40 \u_inFIFO/U718  ( .A(\u_inFIFO/FIFO[36][3] ), .B(
        \u_inFIFO/FIFO[37][3] ), .C(\u_inFIFO/FIFO[38][3] ), .D(
        \u_inFIFO/FIFO[39][3] ), .S0(n13), .S1(\u_inFIFO/N38 ), .Q(
        \u_inFIFO/n738 ) );
  IMUX40 \u_inFIFO/U705  ( .A(\u_inFIFO/FIFO[84][3] ), .B(
        \u_inFIFO/FIFO[85][3] ), .C(\u_inFIFO/FIFO[86][3] ), .D(
        \u_inFIFO/FIFO[87][3] ), .S0(n13), .S1(\u_inFIFO/N38 ), .Q(
        \u_inFIFO/n723 ) );
  IMUX40 \u_inFIFO/U709  ( .A(\u_inFIFO/FIFO[68][3] ), .B(
        \u_inFIFO/FIFO[69][3] ), .C(\u_inFIFO/FIFO[70][3] ), .D(
        \u_inFIFO/FIFO[71][3] ), .S0(n13), .S1(\u_inFIFO/N38 ), .Q(
        \u_inFIFO/n728 ) );
  IMUX40 \u_inFIFO/U701  ( .A(\u_inFIFO/FIFO[100][3] ), .B(
        \u_inFIFO/FIFO[101][3] ), .C(\u_inFIFO/FIFO[102][3] ), .D(
        \u_inFIFO/FIFO[103][3] ), .S0(n1196), .S1(n1201), .Q(\u_inFIFO/n718 )
         );
  IMUX40 \u_inFIFO/U671  ( .A(\u_inFIFO/FIFO[84][2] ), .B(
        \u_inFIFO/FIFO[85][2] ), .C(\u_inFIFO/FIFO[86][2] ), .D(
        \u_inFIFO/FIFO[87][2] ), .S0(n1199), .S1(\u_inFIFO/N38 ), .Q(
        \u_inFIFO/n681 ) );
  IMUX40 \u_inFIFO/U637  ( .A(\u_inFIFO/FIFO[84][1] ), .B(
        \u_inFIFO/FIFO[85][1] ), .C(\u_inFIFO/FIFO[86][1] ), .D(
        \u_inFIFO/FIFO[87][1] ), .S0(n1197), .S1(\u_inFIFO/N38 ), .Q(
        \u_inFIFO/n639 ) );
  IMUX40 \u_inFIFO/U689  ( .A(\u_inFIFO/FIFO[16][2] ), .B(
        \u_inFIFO/FIFO[17][2] ), .C(\u_inFIFO/FIFO[18][2] ), .D(
        \u_inFIFO/FIFO[19][2] ), .S0(n1196), .S1(n764), .Q(\u_inFIFO/n699 ) );
  IMUX40 \u_inFIFO/U687  ( .A(\u_inFIFO/FIFO[24][2] ), .B(
        \u_inFIFO/FIFO[25][2] ), .C(\u_inFIFO/FIFO[26][2] ), .D(
        \u_inFIFO/FIFO[27][2] ), .S0(n1196), .S1(n764), .Q(\u_inFIFO/n700 ) );
  IMUX40 \u_inFIFO/U688  ( .A(\u_inFIFO/FIFO[20][2] ), .B(
        \u_inFIFO/FIFO[21][2] ), .C(\u_inFIFO/FIFO[22][2] ), .D(
        \u_inFIFO/FIFO[23][2] ), .S0(n1196), .S1(n764), .Q(\u_inFIFO/n701 ) );
  IMUX40 \u_inFIFO/U581  ( .A(\u_inFIFO/n699 ), .B(\u_inFIFO/n700 ), .C(
        \u_inFIFO/n701 ), .D(\u_inFIFO/n702 ), .S0(\u_inFIFO/N40 ), .S1(n15), 
        .Q(\u_inFIFO/n698 ) );
  IMUX40 \u_inFIFO/U655  ( .A(\u_inFIFO/FIFO[16][1] ), .B(
        \u_inFIFO/FIFO[17][1] ), .C(\u_inFIFO/FIFO[18][1] ), .D(
        \u_inFIFO/FIFO[19][1] ), .S0(n1199), .S1(n1200), .Q(\u_inFIFO/n657 )
         );
  IMUX40 \u_inFIFO/U653  ( .A(\u_inFIFO/FIFO[24][1] ), .B(
        \u_inFIFO/FIFO[25][1] ), .C(\u_inFIFO/FIFO[26][1] ), .D(
        \u_inFIFO/FIFO[27][1] ), .S0(n1198), .S1(n1200), .Q(\u_inFIFO/n658 )
         );
  IMUX40 \u_inFIFO/U654  ( .A(\u_inFIFO/FIFO[20][1] ), .B(
        \u_inFIFO/FIFO[21][1] ), .C(\u_inFIFO/FIFO[22][1] ), .D(
        \u_inFIFO/FIFO[23][1] ), .S0(n1197), .S1(n1200), .Q(\u_inFIFO/n659 )
         );
  IMUX40 \u_inFIFO/U572  ( .A(\u_inFIFO/n657 ), .B(\u_inFIFO/n658 ), .C(
        \u_inFIFO/n659 ), .D(\u_inFIFO/n660 ), .S0(\u_inFIFO/N40 ), .S1(n15), 
        .Q(\u_inFIFO/n656 ) );
  IMUX40 \u_inFIFO/U604  ( .A(\u_inFIFO/FIFO[80][0] ), .B(
        \u_inFIFO/FIFO[81][0] ), .C(\u_inFIFO/FIFO[82][0] ), .D(
        \u_inFIFO/FIFO[83][0] ), .S0(n1199), .S1(n764), .Q(\u_inFIFO/n595 ) );
  IMUX40 \u_inFIFO/U602  ( .A(\u_inFIFO/FIFO[88][0] ), .B(
        \u_inFIFO/FIFO[89][0] ), .C(\u_inFIFO/FIFO[90][0] ), .D(
        \u_inFIFO/FIFO[91][0] ), .S0(n1199), .S1(n1201), .Q(\u_inFIFO/n596 )
         );
  IMUX40 \u_inFIFO/U603  ( .A(\u_inFIFO/FIFO[84][0] ), .B(
        \u_inFIFO/FIFO[85][0] ), .C(\u_inFIFO/FIFO[86][0] ), .D(
        \u_inFIFO/FIFO[87][0] ), .S0(n1199), .S1(n1201), .Q(\u_inFIFO/n597 )
         );
  IMUX40 \u_inFIFO/U559  ( .A(\u_inFIFO/n595 ), .B(\u_inFIFO/n596 ), .C(
        \u_inFIFO/n597 ), .D(\u_inFIFO/n598 ), .S0(n1202), .S1(n15), .Q(
        \u_inFIFO/n594 ) );
  IMUX40 \u_inFIFO/U621  ( .A(\u_inFIFO/FIFO[16][0] ), .B(
        \u_inFIFO/FIFO[17][0] ), .C(\u_inFIFO/FIFO[18][0] ), .D(
        \u_inFIFO/FIFO[19][0] ), .S0(n1198), .S1(n764), .Q(\u_inFIFO/n615 ) );
  IMUX40 \u_inFIFO/U619  ( .A(\u_inFIFO/FIFO[24][0] ), .B(
        \u_inFIFO/FIFO[25][0] ), .C(\u_inFIFO/FIFO[26][0] ), .D(
        \u_inFIFO/FIFO[27][0] ), .S0(n1198), .S1(n764), .Q(\u_inFIFO/n616 ) );
  IMUX40 \u_inFIFO/U620  ( .A(\u_inFIFO/FIFO[20][0] ), .B(
        \u_inFIFO/FIFO[21][0] ), .C(\u_inFIFO/FIFO[22][0] ), .D(
        \u_inFIFO/FIFO[23][0] ), .S0(n1198), .S1(n764), .Q(\u_inFIFO/n617 ) );
  IMUX40 \u_inFIFO/U563  ( .A(\u_inFIFO/n615 ), .B(\u_inFIFO/n616 ), .C(
        \u_inFIFO/n617 ), .D(\u_inFIFO/n618 ), .S0(n1202), .S1(n15), .Q(
        \u_inFIFO/n614 ) );
  IMUX40 \u_inFIFO/U598  ( .A(\u_inFIFO/FIFO[104][0] ), .B(
        \u_inFIFO/FIFO[105][0] ), .C(\u_inFIFO/FIFO[106][0] ), .D(
        \u_inFIFO/FIFO[107][0] ), .S0(n1199), .S1(n1201), .Q(\u_inFIFO/n591 )
         );
  IMUX40 \u_inFIFO/U597  ( .A(\u_inFIFO/FIFO[108][0] ), .B(
        \u_inFIFO/FIFO[109][0] ), .C(\u_inFIFO/FIFO[110][0] ), .D(
        \u_inFIFO/FIFO[111][0] ), .S0(n1198), .S1(n1201), .Q(\u_inFIFO/n593 )
         );
  IMUX40 \u_inFIFO/U600  ( .A(\u_inFIFO/FIFO[96][0] ), .B(
        \u_inFIFO/FIFO[97][0] ), .C(\u_inFIFO/FIFO[98][0] ), .D(
        \u_inFIFO/FIFO[99][0] ), .S0(n1197), .S1(n1201), .Q(\u_inFIFO/n590 )
         );
  IMUX40 \u_inFIFO/U596  ( .A(\u_inFIFO/FIFO[112][0] ), .B(
        \u_inFIFO/FIFO[113][0] ), .C(\u_inFIFO/FIFO[114][0] ), .D(
        \u_inFIFO/FIFO[115][0] ), .S0(n1196), .S1(n1201), .Q(\u_inFIFO/n585 )
         );
  IMUX40 \u_inFIFO/U721  ( .A(\u_inFIFO/FIFO[24][3] ), .B(
        \u_inFIFO/FIFO[25][3] ), .C(\u_inFIFO/FIFO[26][3] ), .D(
        \u_inFIFO/FIFO[27][3] ), .S0(n13), .S1(\u_inFIFO/N38 ), .Q(
        \u_inFIFO/n742 ) );
  IMUX40 \u_inFIFO/U723  ( .A(\u_inFIFO/FIFO[16][3] ), .B(
        \u_inFIFO/FIFO[17][3] ), .C(\u_inFIFO/FIFO[18][3] ), .D(
        \u_inFIFO/FIFO[19][3] ), .S0(n13), .S1(\u_inFIFO/N38 ), .Q(
        \u_inFIFO/n741 ) );
  IMUX40 \u_inFIFO/U720  ( .A(\u_inFIFO/FIFO[28][3] ), .B(
        \u_inFIFO/FIFO[29][3] ), .C(\u_inFIFO/FIFO[30][3] ), .D(
        \u_inFIFO/FIFO[31][3] ), .S0(n13), .S1(\u_inFIFO/N38 ), .Q(
        \u_inFIFO/n744 ) );
  IMUX40 \u_inFIFO/U713  ( .A(\u_inFIFO/FIFO[56][3] ), .B(
        \u_inFIFO/FIFO[57][3] ), .C(\u_inFIFO/FIFO[58][3] ), .D(
        \u_inFIFO/FIFO[59][3] ), .S0(n13), .S1(n764), .Q(\u_inFIFO/n732 ) );
  IMUX40 \u_inFIFO/U715  ( .A(\u_inFIFO/FIFO[48][3] ), .B(
        \u_inFIFO/FIFO[49][3] ), .C(\u_inFIFO/FIFO[50][3] ), .D(
        \u_inFIFO/FIFO[51][3] ), .S0(n13), .S1(\u_inFIFO/N38 ), .Q(
        \u_inFIFO/n731 ) );
  IMUX40 \u_inFIFO/U712  ( .A(\u_inFIFO/FIFO[60][3] ), .B(
        \u_inFIFO/FIFO[61][3] ), .C(\u_inFIFO/FIFO[62][3] ), .D(
        \u_inFIFO/FIFO[63][3] ), .S0(n13), .S1(n1201), .Q(\u_inFIFO/n734 ) );
  IMUX40 \u_inFIFO/U717  ( .A(\u_inFIFO/FIFO[40][3] ), .B(
        \u_inFIFO/FIFO[41][3] ), .C(\u_inFIFO/FIFO[42][3] ), .D(
        \u_inFIFO/FIFO[43][3] ), .S0(n13), .S1(\u_inFIFO/N38 ), .Q(
        \u_inFIFO/n737 ) );
  IMUX40 \u_inFIFO/U719  ( .A(\u_inFIFO/FIFO[32][3] ), .B(
        \u_inFIFO/FIFO[33][3] ), .C(\u_inFIFO/FIFO[34][3] ), .D(
        \u_inFIFO/FIFO[35][3] ), .S0(n13), .S1(\u_inFIFO/N38 ), .Q(
        \u_inFIFO/n736 ) );
  IMUX40 \u_inFIFO/U716  ( .A(\u_inFIFO/FIFO[44][3] ), .B(
        \u_inFIFO/FIFO[45][3] ), .C(\u_inFIFO/FIFO[46][3] ), .D(
        \u_inFIFO/FIFO[47][3] ), .S0(n13), .S1(\u_inFIFO/N38 ), .Q(
        \u_inFIFO/n739 ) );
  IMUX40 \u_inFIFO/U724  ( .A(\u_inFIFO/FIFO[12][3] ), .B(
        \u_inFIFO/FIFO[13][3] ), .C(\u_inFIFO/FIFO[14][3] ), .D(
        \u_inFIFO/FIFO[15][3] ), .S0(n13), .S1(\u_inFIFO/N38 ), .Q(
        \u_inFIFO/n749 ) );
  IMUX40 \u_inFIFO/U703  ( .A(\u_inFIFO/FIFO[92][3] ), .B(
        \u_inFIFO/FIFO[93][3] ), .C(\u_inFIFO/FIFO[94][3] ), .D(
        \u_inFIFO/FIFO[95][3] ), .S0(n13), .S1(n764), .Q(\u_inFIFO/n724 ) );
  IMUX40 \u_inFIFO/U704  ( .A(\u_inFIFO/FIFO[88][3] ), .B(
        \u_inFIFO/FIFO[89][3] ), .C(\u_inFIFO/FIFO[90][3] ), .D(
        \u_inFIFO/FIFO[91][3] ), .S0(n13), .S1(n1200), .Q(\u_inFIFO/n722 ) );
  IMUX40 \u_inFIFO/U706  ( .A(\u_inFIFO/FIFO[80][3] ), .B(
        \u_inFIFO/FIFO[81][3] ), .C(\u_inFIFO/FIFO[82][3] ), .D(
        \u_inFIFO/FIFO[83][3] ), .S0(n13), .S1(n1200), .Q(\u_inFIFO/n721 ) );
  IMUX40 \u_inFIFO/U707  ( .A(\u_inFIFO/FIFO[76][3] ), .B(
        \u_inFIFO/FIFO[77][3] ), .C(\u_inFIFO/FIFO[78][3] ), .D(
        \u_inFIFO/FIFO[79][3] ), .S0(n13), .S1(\u_inFIFO/N38 ), .Q(
        \u_inFIFO/n729 ) );
  IMUX40 \u_inFIFO/U708  ( .A(\u_inFIFO/FIFO[72][3] ), .B(
        \u_inFIFO/FIFO[73][3] ), .C(\u_inFIFO/FIFO[74][3] ), .D(
        \u_inFIFO/FIFO[75][3] ), .S0(n13), .S1(n764), .Q(\u_inFIFO/n727 ) );
  IMUX40 \u_inFIFO/U710  ( .A(\u_inFIFO/FIFO[64][3] ), .B(
        \u_inFIFO/FIFO[65][3] ), .C(\u_inFIFO/FIFO[66][3] ), .D(
        \u_inFIFO/FIFO[67][3] ), .S0(n13), .S1(\u_inFIFO/N38 ), .Q(
        \u_inFIFO/n726 ) );
  IMUX40 \u_inFIFO/U699  ( .A(\u_inFIFO/FIFO[108][3] ), .B(
        \u_inFIFO/FIFO[109][3] ), .C(\u_inFIFO/FIFO[110][3] ), .D(
        \u_inFIFO/FIFO[111][3] ), .S0(n1199), .S1(n1200), .Q(\u_inFIFO/n719 )
         );
  IMUX40 \u_inFIFO/U700  ( .A(\u_inFIFO/FIFO[104][3] ), .B(
        \u_inFIFO/FIFO[105][3] ), .C(\u_inFIFO/FIFO[106][3] ), .D(
        \u_inFIFO/FIFO[107][3] ), .S0(n1197), .S1(n1200), .Q(\u_inFIFO/n717 )
         );
  IMUX40 \u_inFIFO/U702  ( .A(\u_inFIFO/FIFO[96][3] ), .B(
        \u_inFIFO/FIFO[97][3] ), .C(\u_inFIFO/FIFO[98][3] ), .D(
        \u_inFIFO/FIFO[99][3] ), .S0(n1196), .S1(n764), .Q(\u_inFIFO/n716 ) );
  IMUX40 \u_inFIFO/U698  ( .A(\u_inFIFO/FIFO[112][3] ), .B(
        \u_inFIFO/FIFO[113][3] ), .C(\u_inFIFO/FIFO[114][3] ), .D(
        \u_inFIFO/FIFO[115][3] ), .S0(n1197), .S1(n1201), .Q(\u_inFIFO/n711 )
         );
  IMUX40 \u_inFIFO/U670  ( .A(\u_inFIFO/FIFO[88][2] ), .B(
        \u_inFIFO/FIFO[89][2] ), .C(\u_inFIFO/FIFO[90][2] ), .D(
        \u_inFIFO/FIFO[91][2] ), .S0(n1196), .S1(n764), .Q(\u_inFIFO/n680 ) );
  IMUX40 \u_inFIFO/U672  ( .A(\u_inFIFO/FIFO[80][2] ), .B(
        \u_inFIFO/FIFO[81][2] ), .C(\u_inFIFO/FIFO[82][2] ), .D(
        \u_inFIFO/FIFO[83][2] ), .S0(n1199), .S1(n1200), .Q(\u_inFIFO/n679 )
         );
  IMUX40 \u_inFIFO/U669  ( .A(\u_inFIFO/FIFO[92][2] ), .B(
        \u_inFIFO/FIFO[93][2] ), .C(\u_inFIFO/FIFO[94][2] ), .D(
        \u_inFIFO/FIFO[95][2] ), .S0(n1197), .S1(\u_inFIFO/N38 ), .Q(
        \u_inFIFO/n682 ) );
  IMUX40 \u_inFIFO/U665  ( .A(\u_inFIFO/FIFO[108][2] ), .B(
        \u_inFIFO/FIFO[109][2] ), .C(\u_inFIFO/FIFO[110][2] ), .D(
        \u_inFIFO/FIFO[111][2] ), .S0(n1199), .S1(n1200), .Q(\u_inFIFO/n677 )
         );
  IMUX40 \u_inFIFO/U673  ( .A(\u_inFIFO/FIFO[76][2] ), .B(
        \u_inFIFO/FIFO[77][2] ), .C(\u_inFIFO/FIFO[78][2] ), .D(
        \u_inFIFO/FIFO[79][2] ), .S0(n1197), .S1(\u_inFIFO/N38 ), .Q(
        \u_inFIFO/n687 ) );
  IMUX40 \u_inFIFO/U664  ( .A(\u_inFIFO/FIFO[112][2] ), .B(
        \u_inFIFO/FIFO[113][2] ), .C(\u_inFIFO/FIFO[114][2] ), .D(
        \u_inFIFO/FIFO[115][2] ), .S0(n1196), .S1(n1200), .Q(\u_inFIFO/n669 )
         );
  IMUX40 \u_inFIFO/U686  ( .A(\u_inFIFO/FIFO[28][2] ), .B(
        \u_inFIFO/FIFO[29][2] ), .C(\u_inFIFO/FIFO[30][2] ), .D(
        \u_inFIFO/FIFO[31][2] ), .S0(n1196), .S1(n764), .Q(\u_inFIFO/n702 ) );
  IMUX40 \u_inFIFO/U678  ( .A(\u_inFIFO/FIFO[60][2] ), .B(
        \u_inFIFO/FIFO[61][2] ), .C(\u_inFIFO/FIFO[62][2] ), .D(
        \u_inFIFO/FIFO[63][2] ), .S0(n1196), .S1(n1201), .Q(\u_inFIFO/n692 )
         );
  IMUX40 \u_inFIFO/U682  ( .A(\u_inFIFO/FIFO[44][2] ), .B(
        \u_inFIFO/FIFO[45][2] ), .C(\u_inFIFO/FIFO[46][2] ), .D(
        \u_inFIFO/FIFO[47][2] ), .S0(n1196), .S1(n764), .Q(\u_inFIFO/n697 ) );
  IMUX40 \u_inFIFO/U690  ( .A(\u_inFIFO/FIFO[12][2] ), .B(
        \u_inFIFO/FIFO[13][2] ), .C(\u_inFIFO/FIFO[14][2] ), .D(
        \u_inFIFO/FIFO[15][2] ), .S0(n1198), .S1(n764), .Q(\u_inFIFO/n707 ) );
  IMUX40 \u_inFIFO/U636  ( .A(\u_inFIFO/FIFO[88][1] ), .B(
        \u_inFIFO/FIFO[89][1] ), .C(\u_inFIFO/FIFO[90][1] ), .D(
        \u_inFIFO/FIFO[91][1] ), .S0(n1198), .S1(\u_inFIFO/N38 ), .Q(
        \u_inFIFO/n638 ) );
  IMUX40 \u_inFIFO/U638  ( .A(\u_inFIFO/FIFO[80][1] ), .B(
        \u_inFIFO/FIFO[81][1] ), .C(\u_inFIFO/FIFO[82][1] ), .D(
        \u_inFIFO/FIFO[83][1] ), .S0(n1199), .S1(\u_inFIFO/N38 ), .Q(
        \u_inFIFO/n637 ) );
  IMUX40 \u_inFIFO/U635  ( .A(\u_inFIFO/FIFO[92][1] ), .B(
        \u_inFIFO/FIFO[93][1] ), .C(\u_inFIFO/FIFO[94][1] ), .D(
        \u_inFIFO/FIFO[95][1] ), .S0(n1198), .S1(\u_inFIFO/N38 ), .Q(
        \u_inFIFO/n640 ) );
  IMUX40 \u_inFIFO/U631  ( .A(\u_inFIFO/FIFO[108][1] ), .B(
        \u_inFIFO/FIFO[109][1] ), .C(\u_inFIFO/FIFO[110][1] ), .D(
        \u_inFIFO/FIFO[111][1] ), .S0(n1196), .S1(\u_inFIFO/N38 ), .Q(
        \u_inFIFO/n635 ) );
  IMUX40 \u_inFIFO/U639  ( .A(\u_inFIFO/FIFO[76][1] ), .B(
        \u_inFIFO/FIFO[77][1] ), .C(\u_inFIFO/FIFO[78][1] ), .D(
        \u_inFIFO/FIFO[79][1] ), .S0(n1197), .S1(\u_inFIFO/N38 ), .Q(
        \u_inFIFO/n645 ) );
  IMUX40 \u_inFIFO/U630  ( .A(\u_inFIFO/FIFO[112][1] ), .B(
        \u_inFIFO/FIFO[113][1] ), .C(\u_inFIFO/FIFO[114][1] ), .D(
        \u_inFIFO/FIFO[115][1] ), .S0(n1196), .S1(n1201), .Q(\u_inFIFO/n627 )
         );
  IMUX40 \u_inFIFO/U652  ( .A(\u_inFIFO/FIFO[28][1] ), .B(
        \u_inFIFO/FIFO[29][1] ), .C(\u_inFIFO/FIFO[30][1] ), .D(
        \u_inFIFO/FIFO[31][1] ), .S0(n13), .S1(n1200), .Q(\u_inFIFO/n660 ) );
  IMUX40 \u_inFIFO/U644  ( .A(\u_inFIFO/FIFO[60][1] ), .B(
        \u_inFIFO/FIFO[61][1] ), .C(\u_inFIFO/FIFO[62][1] ), .D(
        \u_inFIFO/FIFO[63][1] ), .S0(n1197), .S1(\u_inFIFO/N38 ), .Q(
        \u_inFIFO/n650 ) );
  IMUX40 \u_inFIFO/U648  ( .A(\u_inFIFO/FIFO[44][1] ), .B(
        \u_inFIFO/FIFO[45][1] ), .C(\u_inFIFO/FIFO[46][1] ), .D(
        \u_inFIFO/FIFO[47][1] ), .S0(n1197), .S1(n1200), .Q(\u_inFIFO/n655 )
         );
  IMUX40 \u_inFIFO/U656  ( .A(\u_inFIFO/FIFO[12][1] ), .B(
        \u_inFIFO/FIFO[13][1] ), .C(\u_inFIFO/FIFO[14][1] ), .D(
        \u_inFIFO/FIFO[15][1] ), .S0(n1198), .S1(n1200), .Q(\u_inFIFO/n665 )
         );
  IMUX40 \u_inFIFO/U601  ( .A(\u_inFIFO/FIFO[92][0] ), .B(
        \u_inFIFO/FIFO[93][0] ), .C(\u_inFIFO/FIFO[94][0] ), .D(
        \u_inFIFO/FIFO[95][0] ), .S0(n1199), .S1(n1201), .Q(\u_inFIFO/n598 )
         );
  IMUX40 \u_inFIFO/U605  ( .A(\u_inFIFO/FIFO[76][0] ), .B(
        \u_inFIFO/FIFO[77][0] ), .C(\u_inFIFO/FIFO[78][0] ), .D(
        \u_inFIFO/FIFO[79][0] ), .S0(n1199), .S1(n1201), .Q(\u_inFIFO/n603 )
         );
  IMUX40 \u_inFIFO/U618  ( .A(\u_inFIFO/FIFO[28][0] ), .B(
        \u_inFIFO/FIFO[29][0] ), .C(\u_inFIFO/FIFO[30][0] ), .D(
        \u_inFIFO/FIFO[31][0] ), .S0(n1198), .S1(\u_inFIFO/N38 ), .Q(
        \u_inFIFO/n618 ) );
  IMUX40 \u_inFIFO/U610  ( .A(\u_inFIFO/FIFO[60][0] ), .B(
        \u_inFIFO/FIFO[61][0] ), .C(\u_inFIFO/FIFO[62][0] ), .D(
        \u_inFIFO/FIFO[63][0] ), .S0(n1199), .S1(n1201), .Q(\u_inFIFO/n608 )
         );
  IMUX40 \u_inFIFO/U614  ( .A(\u_inFIFO/FIFO[44][0] ), .B(
        \u_inFIFO/FIFO[45][0] ), .C(\u_inFIFO/FIFO[46][0] ), .D(
        \u_inFIFO/FIFO[47][0] ), .S0(n1198), .S1(\u_inFIFO/N38 ), .Q(
        \u_inFIFO/n613 ) );
  IMUX40 \u_inFIFO/U622  ( .A(\u_inFIFO/FIFO[12][0] ), .B(
        \u_inFIFO/FIFO[13][0] ), .C(\u_inFIFO/FIFO[14][0] ), .D(
        \u_inFIFO/FIFO[15][0] ), .S0(n1198), .S1(\u_inFIFO/N38 ), .Q(
        \u_inFIFO/n623 ) );
  IMUX40 \u_inFIFO/U727  ( .A(\u_inFIFO/FIFO[0][3] ), .B(\u_inFIFO/FIFO[1][3] ), .C(\u_inFIFO/FIFO[2][3] ), .D(\u_inFIFO/FIFO[3][3] ), .S0(n13), .S1(n1200), 
        .Q(\u_inFIFO/n746 ) );
  IMUX40 \u_inFIFO/U725  ( .A(\u_inFIFO/FIFO[8][3] ), .B(\u_inFIFO/FIFO[9][3] ), .C(\u_inFIFO/FIFO[10][3] ), .D(\u_inFIFO/FIFO[11][3] ), .S0(n13), .S1(
        \u_inFIFO/N38 ), .Q(\u_inFIFO/n747 ) );
  IMUX40 \u_inFIFO/U726  ( .A(\u_inFIFO/FIFO[4][3] ), .B(\u_inFIFO/FIFO[5][3] ), .C(\u_inFIFO/FIFO[6][3] ), .D(\u_inFIFO/FIFO[7][3] ), .S0(n13), .S1(
        \u_inFIFO/N38 ), .Q(\u_inFIFO/n748 ) );
  IMUX40 \u_inFIFO/U591  ( .A(\u_inFIFO/n746 ), .B(\u_inFIFO/n747 ), .C(
        \u_inFIFO/n748 ), .D(\u_inFIFO/n749 ), .S0(\u_inFIFO/N40 ), .S1(n15), 
        .Q(\u_inFIFO/n745 ) );
  IMUX40 \u_inFIFO/U696  ( .A(\u_inFIFO/FIFO[120][3] ), .B(
        \u_inFIFO/FIFO[121][3] ), .C(\u_inFIFO/FIFO[122][3] ), .D(
        \u_inFIFO/FIFO[123][3] ), .S0(n1197), .S1(n764), .Q(\u_inFIFO/n712 )
         );
  IMUX40 \u_inFIFO/U695  ( .A(\u_inFIFO/FIFO[124][3] ), .B(
        \u_inFIFO/FIFO[125][3] ), .C(\u_inFIFO/FIFO[126][3] ), .D(
        \u_inFIFO/FIFO[127][3] ), .S0(n1199), .S1(n1201), .Q(\u_inFIFO/n714 )
         );
  IMUX40 \u_inFIFO/U697  ( .A(\u_inFIFO/FIFO[116][3] ), .B(
        \u_inFIFO/FIFO[117][3] ), .C(\u_inFIFO/FIFO[118][3] ), .D(
        \u_inFIFO/FIFO[119][3] ), .S0(n1198), .S1(n764), .Q(\u_inFIFO/n713 )
         );
  IMUX40 \u_inFIFO/U584  ( .A(\u_inFIFO/n711 ), .B(\u_inFIFO/n712 ), .C(
        \u_inFIFO/n713 ), .D(\u_inFIFO/n714 ), .S0(\u_inFIFO/N40 ), .S1(n15), 
        .Q(\u_inFIFO/n710 ) );
  IMUX40 \u_inFIFO/U668  ( .A(\u_inFIFO/FIFO[96][2] ), .B(
        \u_inFIFO/FIFO[97][2] ), .C(\u_inFIFO/FIFO[98][2] ), .D(
        \u_inFIFO/FIFO[99][2] ), .S0(n1197), .S1(n1201), .Q(\u_inFIFO/n674 )
         );
  IMUX40 \u_inFIFO/U666  ( .A(\u_inFIFO/FIFO[104][2] ), .B(
        \u_inFIFO/FIFO[105][2] ), .C(\u_inFIFO/FIFO[106][2] ), .D(
        \u_inFIFO/FIFO[107][2] ), .S0(n1198), .S1(n1201), .Q(\u_inFIFO/n675 )
         );
  IMUX40 \u_inFIFO/U667  ( .A(\u_inFIFO/FIFO[100][2] ), .B(
        \u_inFIFO/FIFO[101][2] ), .C(\u_inFIFO/FIFO[102][2] ), .D(
        \u_inFIFO/FIFO[103][2] ), .S0(n1196), .S1(\u_inFIFO/N38 ), .Q(
        \u_inFIFO/n676 ) );
  IMUX40 \u_inFIFO/U576  ( .A(\u_inFIFO/n674 ), .B(\u_inFIFO/n675 ), .C(
        \u_inFIFO/n676 ), .D(\u_inFIFO/n677 ), .S0(\u_inFIFO/N40 ), .S1(n15), 
        .Q(\u_inFIFO/n673 ) );
  IMUX40 \u_inFIFO/U676  ( .A(\u_inFIFO/FIFO[64][2] ), .B(
        \u_inFIFO/FIFO[65][2] ), .C(\u_inFIFO/FIFO[66][2] ), .D(
        \u_inFIFO/FIFO[67][2] ), .S0(n1199), .S1(n1201), .Q(\u_inFIFO/n684 )
         );
  IMUX40 \u_inFIFO/U674  ( .A(\u_inFIFO/FIFO[72][2] ), .B(
        \u_inFIFO/FIFO[73][2] ), .C(\u_inFIFO/FIFO[74][2] ), .D(
        \u_inFIFO/FIFO[75][2] ), .S0(n1199), .S1(\u_inFIFO/N38 ), .Q(
        \u_inFIFO/n685 ) );
  IMUX40 \u_inFIFO/U675  ( .A(\u_inFIFO/FIFO[68][2] ), .B(
        \u_inFIFO/FIFO[69][2] ), .C(\u_inFIFO/FIFO[70][2] ), .D(
        \u_inFIFO/FIFO[71][2] ), .S0(n1199), .S1(n1200), .Q(\u_inFIFO/n686 )
         );
  IMUX40 \u_inFIFO/U578  ( .A(\u_inFIFO/n684 ), .B(\u_inFIFO/n685 ), .C(
        \u_inFIFO/n686 ), .D(\u_inFIFO/n687 ), .S0(\u_inFIFO/N40 ), .S1(n15), 
        .Q(\u_inFIFO/n683 ) );
  IMUX40 \u_inFIFO/U662  ( .A(\u_inFIFO/FIFO[120][2] ), .B(
        \u_inFIFO/FIFO[121][2] ), .C(\u_inFIFO/FIFO[122][2] ), .D(
        \u_inFIFO/FIFO[123][2] ), .S0(n1196), .S1(n1200), .Q(\u_inFIFO/n670 )
         );
  IMUX40 \u_inFIFO/U661  ( .A(\u_inFIFO/FIFO[124][2] ), .B(
        \u_inFIFO/FIFO[125][2] ), .C(\u_inFIFO/FIFO[126][2] ), .D(
        \u_inFIFO/FIFO[127][2] ), .S0(n1196), .S1(n1200), .Q(\u_inFIFO/n672 )
         );
  IMUX40 \u_inFIFO/U663  ( .A(\u_inFIFO/FIFO[116][2] ), .B(
        \u_inFIFO/FIFO[117][2] ), .C(\u_inFIFO/FIFO[118][2] ), .D(
        \u_inFIFO/FIFO[119][2] ), .S0(n1199), .S1(n1200), .Q(\u_inFIFO/n671 )
         );
  IMUX40 \u_inFIFO/U575  ( .A(\u_inFIFO/n669 ), .B(\u_inFIFO/n670 ), .C(
        \u_inFIFO/n671 ), .D(\u_inFIFO/n672 ), .S0(n1202), .S1(n15), .Q(
        \u_inFIFO/n668 ) );
  IMUX40 \u_inFIFO/U681  ( .A(\u_inFIFO/FIFO[48][2] ), .B(
        \u_inFIFO/FIFO[49][2] ), .C(\u_inFIFO/FIFO[50][2] ), .D(
        \u_inFIFO/FIFO[51][2] ), .S0(n1196), .S1(n764), .Q(\u_inFIFO/n689 ) );
  IMUX40 \u_inFIFO/U679  ( .A(\u_inFIFO/FIFO[56][2] ), .B(
        \u_inFIFO/FIFO[57][2] ), .C(\u_inFIFO/FIFO[58][2] ), .D(
        \u_inFIFO/FIFO[59][2] ), .S0(n1196), .S1(\u_inFIFO/N38 ), .Q(
        \u_inFIFO/n690 ) );
  IMUX40 \u_inFIFO/U680  ( .A(\u_inFIFO/FIFO[52][2] ), .B(
        \u_inFIFO/FIFO[53][2] ), .C(\u_inFIFO/FIFO[54][2] ), .D(
        \u_inFIFO/FIFO[55][2] ), .S0(n1196), .S1(n1200), .Q(\u_inFIFO/n691 )
         );
  IMUX40 \u_inFIFO/U579  ( .A(\u_inFIFO/n689 ), .B(\u_inFIFO/n690 ), .C(
        \u_inFIFO/n691 ), .D(\u_inFIFO/n692 ), .S0(\u_inFIFO/N40 ), .S1(n15), 
        .Q(\u_inFIFO/n688 ) );
  IMUX40 \u_inFIFO/U685  ( .A(\u_inFIFO/FIFO[32][2] ), .B(
        \u_inFIFO/FIFO[33][2] ), .C(\u_inFIFO/FIFO[34][2] ), .D(
        \u_inFIFO/FIFO[35][2] ), .S0(n1196), .S1(n764), .Q(\u_inFIFO/n694 ) );
  IMUX40 \u_inFIFO/U683  ( .A(\u_inFIFO/FIFO[40][2] ), .B(
        \u_inFIFO/FIFO[41][2] ), .C(\u_inFIFO/FIFO[42][2] ), .D(
        \u_inFIFO/FIFO[43][2] ), .S0(n1196), .S1(n764), .Q(\u_inFIFO/n695 ) );
  IMUX40 \u_inFIFO/U684  ( .A(\u_inFIFO/FIFO[36][2] ), .B(
        \u_inFIFO/FIFO[37][2] ), .C(\u_inFIFO/FIFO[38][2] ), .D(
        \u_inFIFO/FIFO[39][2] ), .S0(n1196), .S1(n764), .Q(\u_inFIFO/n696 ) );
  IMUX40 \u_inFIFO/U580  ( .A(\u_inFIFO/n694 ), .B(\u_inFIFO/n695 ), .C(
        \u_inFIFO/n696 ), .D(\u_inFIFO/n697 ), .S0(\u_inFIFO/N40 ), .S1(n15), 
        .Q(\u_inFIFO/n693 ) );
  IMUX40 \u_inFIFO/U693  ( .A(\u_inFIFO/FIFO[0][2] ), .B(\u_inFIFO/FIFO[1][2] ), .C(\u_inFIFO/FIFO[2][2] ), .D(\u_inFIFO/FIFO[3][2] ), .S0(n13), .S1(n764), 
        .Q(\u_inFIFO/n704 ) );
  IMUX40 \u_inFIFO/U691  ( .A(\u_inFIFO/FIFO[8][2] ), .B(\u_inFIFO/FIFO[9][2] ), .C(\u_inFIFO/FIFO[10][2] ), .D(\u_inFIFO/FIFO[11][2] ), .S0(n1199), .S1(n764), .Q(\u_inFIFO/n705 ) );
  IMUX40 \u_inFIFO/U692  ( .A(\u_inFIFO/FIFO[4][2] ), .B(\u_inFIFO/FIFO[5][2] ), .C(\u_inFIFO/FIFO[6][2] ), .D(\u_inFIFO/FIFO[7][2] ), .S0(n1198), .S1(n764), 
        .Q(\u_inFIFO/n706 ) );
  IMUX40 \u_inFIFO/U582  ( .A(\u_inFIFO/n704 ), .B(\u_inFIFO/n705 ), .C(
        \u_inFIFO/n706 ), .D(\u_inFIFO/n707 ), .S0(\u_inFIFO/N40 ), .S1(n15), 
        .Q(\u_inFIFO/n703 ) );
  IMUX40 \u_inFIFO/U634  ( .A(\u_inFIFO/FIFO[96][1] ), .B(
        \u_inFIFO/FIFO[97][1] ), .C(\u_inFIFO/FIFO[98][1] ), .D(
        \u_inFIFO/FIFO[99][1] ), .S0(n1197), .S1(\u_inFIFO/N38 ), .Q(
        \u_inFIFO/n632 ) );
  IMUX40 \u_inFIFO/U632  ( .A(\u_inFIFO/FIFO[104][1] ), .B(
        \u_inFIFO/FIFO[105][1] ), .C(\u_inFIFO/FIFO[106][1] ), .D(
        \u_inFIFO/FIFO[107][1] ), .S0(n1198), .S1(\u_inFIFO/N38 ), .Q(
        \u_inFIFO/n633 ) );
  IMUX40 \u_inFIFO/U633  ( .A(\u_inFIFO/FIFO[100][1] ), .B(
        \u_inFIFO/FIFO[101][1] ), .C(\u_inFIFO/FIFO[102][1] ), .D(
        \u_inFIFO/FIFO[103][1] ), .S0(n1198), .S1(\u_inFIFO/N38 ), .Q(
        \u_inFIFO/n634 ) );
  IMUX40 \u_inFIFO/U567  ( .A(\u_inFIFO/n632 ), .B(\u_inFIFO/n633 ), .C(
        \u_inFIFO/n634 ), .D(\u_inFIFO/n635 ), .S0(\u_inFIFO/N40 ), .S1(n15), 
        .Q(\u_inFIFO/n631 ) );
  IMUX40 \u_inFIFO/U642  ( .A(\u_inFIFO/FIFO[64][1] ), .B(
        \u_inFIFO/FIFO[65][1] ), .C(\u_inFIFO/FIFO[66][1] ), .D(
        \u_inFIFO/FIFO[67][1] ), .S0(n1197), .S1(\u_inFIFO/N38 ), .Q(
        \u_inFIFO/n642 ) );
  IMUX40 \u_inFIFO/U640  ( .A(\u_inFIFO/FIFO[72][1] ), .B(
        \u_inFIFO/FIFO[73][1] ), .C(\u_inFIFO/FIFO[74][1] ), .D(
        \u_inFIFO/FIFO[75][1] ), .S0(n1197), .S1(\u_inFIFO/N38 ), .Q(
        \u_inFIFO/n643 ) );
  IMUX40 \u_inFIFO/U641  ( .A(\u_inFIFO/FIFO[68][1] ), .B(
        \u_inFIFO/FIFO[69][1] ), .C(\u_inFIFO/FIFO[70][1] ), .D(
        \u_inFIFO/FIFO[71][1] ), .S0(n1197), .S1(\u_inFIFO/N38 ), .Q(
        \u_inFIFO/n644 ) );
  IMUX40 \u_inFIFO/U569  ( .A(\u_inFIFO/n642 ), .B(\u_inFIFO/n643 ), .C(
        \u_inFIFO/n644 ), .D(\u_inFIFO/n645 ), .S0(\u_inFIFO/N40 ), .S1(n15), 
        .Q(\u_inFIFO/n641 ) );
  IMUX40 \u_inFIFO/U628  ( .A(\u_inFIFO/FIFO[120][1] ), .B(
        \u_inFIFO/FIFO[121][1] ), .C(\u_inFIFO/FIFO[122][1] ), .D(
        \u_inFIFO/FIFO[123][1] ), .S0(n1196), .S1(\u_inFIFO/N38 ), .Q(
        \u_inFIFO/n628 ) );
  IMUX40 \u_inFIFO/U627  ( .A(\u_inFIFO/FIFO[124][1] ), .B(
        \u_inFIFO/FIFO[125][1] ), .C(\u_inFIFO/FIFO[126][1] ), .D(
        \u_inFIFO/FIFO[127][1] ), .S0(n1197), .S1(\u_inFIFO/N38 ), .Q(
        \u_inFIFO/n630 ) );
  IMUX40 \u_inFIFO/U629  ( .A(\u_inFIFO/FIFO[116][1] ), .B(
        \u_inFIFO/FIFO[117][1] ), .C(\u_inFIFO/FIFO[118][1] ), .D(
        \u_inFIFO/FIFO[119][1] ), .S0(n1197), .S1(\u_inFIFO/N38 ), .Q(
        \u_inFIFO/n629 ) );
  IMUX40 \u_inFIFO/U566  ( .A(\u_inFIFO/n627 ), .B(\u_inFIFO/n628 ), .C(
        \u_inFIFO/n629 ), .D(\u_inFIFO/n630 ), .S0(n1202), .S1(n15), .Q(
        \u_inFIFO/n626 ) );
  IMUX40 \u_inFIFO/U647  ( .A(\u_inFIFO/FIFO[48][1] ), .B(
        \u_inFIFO/FIFO[49][1] ), .C(\u_inFIFO/FIFO[50][1] ), .D(
        \u_inFIFO/FIFO[51][1] ), .S0(n1197), .S1(\u_inFIFO/N38 ), .Q(
        \u_inFIFO/n647 ) );
  IMUX40 \u_inFIFO/U645  ( .A(\u_inFIFO/FIFO[56][1] ), .B(
        \u_inFIFO/FIFO[57][1] ), .C(\u_inFIFO/FIFO[58][1] ), .D(
        \u_inFIFO/FIFO[59][1] ), .S0(n1197), .S1(\u_inFIFO/N38 ), .Q(
        \u_inFIFO/n648 ) );
  IMUX40 \u_inFIFO/U646  ( .A(\u_inFIFO/FIFO[52][1] ), .B(
        \u_inFIFO/FIFO[53][1] ), .C(\u_inFIFO/FIFO[54][1] ), .D(
        \u_inFIFO/FIFO[55][1] ), .S0(n1197), .S1(\u_inFIFO/N38 ), .Q(
        \u_inFIFO/n649 ) );
  IMUX40 \u_inFIFO/U570  ( .A(\u_inFIFO/n647 ), .B(\u_inFIFO/n648 ), .C(
        \u_inFIFO/n649 ), .D(\u_inFIFO/n650 ), .S0(n1202), .S1(n15), .Q(
        \u_inFIFO/n646 ) );
  IMUX40 \u_inFIFO/U651  ( .A(\u_inFIFO/FIFO[32][1] ), .B(
        \u_inFIFO/FIFO[33][1] ), .C(\u_inFIFO/FIFO[34][1] ), .D(
        \u_inFIFO/FIFO[35][1] ), .S0(n1197), .S1(n1200), .Q(\u_inFIFO/n652 )
         );
  IMUX40 \u_inFIFO/U649  ( .A(\u_inFIFO/FIFO[40][1] ), .B(
        \u_inFIFO/FIFO[41][1] ), .C(\u_inFIFO/FIFO[42][1] ), .D(
        \u_inFIFO/FIFO[43][1] ), .S0(n1197), .S1(n1200), .Q(\u_inFIFO/n653 )
         );
  IMUX40 \u_inFIFO/U650  ( .A(\u_inFIFO/FIFO[36][1] ), .B(
        \u_inFIFO/FIFO[37][1] ), .C(\u_inFIFO/FIFO[38][1] ), .D(
        \u_inFIFO/FIFO[39][1] ), .S0(n1197), .S1(n1200), .Q(\u_inFIFO/n654 )
         );
  IMUX40 \u_inFIFO/U571  ( .A(\u_inFIFO/n652 ), .B(\u_inFIFO/n653 ), .C(
        \u_inFIFO/n654 ), .D(\u_inFIFO/n655 ), .S0(\u_inFIFO/N40 ), .S1(n15), 
        .Q(\u_inFIFO/n651 ) );
  IMUX40 \u_inFIFO/U659  ( .A(\u_inFIFO/FIFO[0][1] ), .B(\u_inFIFO/FIFO[1][1] ), .C(\u_inFIFO/FIFO[2][1] ), .D(\u_inFIFO/FIFO[3][1] ), .S0(n13), .S1(n1200), 
        .Q(\u_inFIFO/n662 ) );
  IMUX40 \u_inFIFO/U657  ( .A(\u_inFIFO/FIFO[8][1] ), .B(\u_inFIFO/FIFO[9][1] ), .C(\u_inFIFO/FIFO[10][1] ), .D(\u_inFIFO/FIFO[11][1] ), .S0(n1196), .S1(
        n1200), .Q(\u_inFIFO/n663 ) );
  IMUX40 \u_inFIFO/U658  ( .A(\u_inFIFO/FIFO[4][1] ), .B(\u_inFIFO/FIFO[5][1] ), .C(\u_inFIFO/FIFO[6][1] ), .D(\u_inFIFO/FIFO[7][1] ), .S0(n13), .S1(n1200), 
        .Q(\u_inFIFO/n664 ) );
  IMUX40 \u_inFIFO/U573  ( .A(\u_inFIFO/n662 ), .B(\u_inFIFO/n663 ), .C(
        \u_inFIFO/n664 ), .D(\u_inFIFO/n665 ), .S0(\u_inFIFO/N40 ), .S1(n15), 
        .Q(\u_inFIFO/n661 ) );
  IMUX40 \u_inFIFO/U594  ( .A(\u_inFIFO/FIFO[120][0] ), .B(
        \u_inFIFO/FIFO[121][0] ), .C(\u_inFIFO/FIFO[122][0] ), .D(
        \u_inFIFO/FIFO[123][0] ), .S0(n1198), .S1(n1201), .Q(\u_inFIFO/n586 )
         );
  IMUX40 \u_inFIFO/U593  ( .A(\u_inFIFO/FIFO[124][0] ), .B(
        \u_inFIFO/FIFO[125][0] ), .C(\u_inFIFO/FIFO[126][0] ), .D(
        \u_inFIFO/FIFO[127][0] ), .S0(n1197), .S1(\u_inFIFO/N38 ), .Q(
        \u_inFIFO/n588 ) );
  IMUX40 \u_inFIFO/U595  ( .A(\u_inFIFO/FIFO[116][0] ), .B(
        \u_inFIFO/FIFO[117][0] ), .C(\u_inFIFO/FIFO[118][0] ), .D(
        \u_inFIFO/FIFO[119][0] ), .S0(n1198), .S1(n1201), .Q(\u_inFIFO/n587 )
         );
  IMUX40 \u_inFIFO/U557  ( .A(\u_inFIFO/n585 ), .B(\u_inFIFO/n586 ), .C(
        \u_inFIFO/n587 ), .D(\u_inFIFO/n588 ), .S0(n1202), .S1(n15), .Q(
        \u_inFIFO/n584 ) );
  IMUX40 \u_inFIFO/U608  ( .A(\u_inFIFO/FIFO[64][0] ), .B(
        \u_inFIFO/FIFO[65][0] ), .C(\u_inFIFO/FIFO[66][0] ), .D(
        \u_inFIFO/FIFO[67][0] ), .S0(n1199), .S1(n764), .Q(\u_inFIFO/n600 ) );
  IMUX40 \u_inFIFO/U606  ( .A(\u_inFIFO/FIFO[72][0] ), .B(
        \u_inFIFO/FIFO[73][0] ), .C(\u_inFIFO/FIFO[74][0] ), .D(
        \u_inFIFO/FIFO[75][0] ), .S0(n1199), .S1(n1201), .Q(\u_inFIFO/n601 )
         );
  IMUX40 \u_inFIFO/U607  ( .A(\u_inFIFO/FIFO[68][0] ), .B(
        \u_inFIFO/FIFO[69][0] ), .C(\u_inFIFO/FIFO[70][0] ), .D(
        \u_inFIFO/FIFO[71][0] ), .S0(n1199), .S1(n1201), .Q(\u_inFIFO/n602 )
         );
  IMUX40 \u_inFIFO/U560  ( .A(\u_inFIFO/n600 ), .B(\u_inFIFO/n601 ), .C(
        \u_inFIFO/n602 ), .D(\u_inFIFO/n603 ), .S0(n1202), .S1(n15), .Q(
        \u_inFIFO/n599 ) );
  IMUX40 \u_inFIFO/U613  ( .A(\u_inFIFO/FIFO[48][0] ), .B(
        \u_inFIFO/FIFO[49][0] ), .C(\u_inFIFO/FIFO[50][0] ), .D(
        \u_inFIFO/FIFO[51][0] ), .S0(n1199), .S1(\u_inFIFO/N38 ), .Q(
        \u_inFIFO/n605 ) );
  IMUX40 \u_inFIFO/U611  ( .A(\u_inFIFO/FIFO[56][0] ), .B(
        \u_inFIFO/FIFO[57][0] ), .C(\u_inFIFO/FIFO[58][0] ), .D(
        \u_inFIFO/FIFO[59][0] ), .S0(n1199), .S1(n1201), .Q(\u_inFIFO/n606 )
         );
  IMUX40 \u_inFIFO/U612  ( .A(\u_inFIFO/FIFO[52][0] ), .B(
        \u_inFIFO/FIFO[53][0] ), .C(\u_inFIFO/FIFO[54][0] ), .D(
        \u_inFIFO/FIFO[55][0] ), .S0(n1199), .S1(n1201), .Q(\u_inFIFO/n607 )
         );
  IMUX40 \u_inFIFO/U561  ( .A(\u_inFIFO/n605 ), .B(\u_inFIFO/n606 ), .C(
        \u_inFIFO/n607 ), .D(\u_inFIFO/n608 ), .S0(n1202), .S1(n15), .Q(
        \u_inFIFO/n604 ) );
  IMUX40 \u_inFIFO/U617  ( .A(\u_inFIFO/FIFO[32][0] ), .B(
        \u_inFIFO/FIFO[33][0] ), .C(\u_inFIFO/FIFO[34][0] ), .D(
        \u_inFIFO/FIFO[35][0] ), .S0(n1198), .S1(n764), .Q(\u_inFIFO/n610 ) );
  IMUX40 \u_inFIFO/U615  ( .A(\u_inFIFO/FIFO[40][0] ), .B(
        \u_inFIFO/FIFO[41][0] ), .C(\u_inFIFO/FIFO[42][0] ), .D(
        \u_inFIFO/FIFO[43][0] ), .S0(n1198), .S1(\u_inFIFO/N38 ), .Q(
        \u_inFIFO/n611 ) );
  IMUX40 \u_inFIFO/U616  ( .A(\u_inFIFO/FIFO[36][0] ), .B(
        \u_inFIFO/FIFO[37][0] ), .C(\u_inFIFO/FIFO[38][0] ), .D(
        \u_inFIFO/FIFO[39][0] ), .S0(n1198), .S1(\u_inFIFO/N38 ), .Q(
        \u_inFIFO/n612 ) );
  IMUX40 \u_inFIFO/U562  ( .A(\u_inFIFO/n610 ), .B(\u_inFIFO/n611 ), .C(
        \u_inFIFO/n612 ), .D(\u_inFIFO/n613 ), .S0(n1202), .S1(n15), .Q(
        \u_inFIFO/n609 ) );
  IMUX40 \u_inFIFO/U625  ( .A(\u_inFIFO/FIFO[0][0] ), .B(\u_inFIFO/FIFO[1][0] ), .C(\u_inFIFO/FIFO[2][0] ), .D(\u_inFIFO/FIFO[3][0] ), .S0(n1198), .S1(n764), 
        .Q(\u_inFIFO/n620 ) );
  IMUX40 \u_inFIFO/U623  ( .A(\u_inFIFO/FIFO[8][0] ), .B(\u_inFIFO/FIFO[9][0] ), .C(\u_inFIFO/FIFO[10][0] ), .D(\u_inFIFO/FIFO[11][0] ), .S0(n1198), .S1(n764), .Q(\u_inFIFO/n621 ) );
  IMUX40 \u_inFIFO/U624  ( .A(\u_inFIFO/FIFO[4][0] ), .B(\u_inFIFO/FIFO[5][0] ), .C(\u_inFIFO/FIFO[6][0] ), .D(\u_inFIFO/FIFO[7][0] ), .S0(n1198), .S1(n764), 
        .Q(\u_inFIFO/n622 ) );
  IMUX40 \u_inFIFO/U564  ( .A(\u_inFIFO/n620 ), .B(\u_inFIFO/n621 ), .C(
        \u_inFIFO/n622 ), .D(\u_inFIFO/n623 ), .S0(n1202), .S1(n15), .Q(
        \u_inFIFO/n619 ) );
  IMUX21 \u_cordic/mycordic/U553  ( .A(\u_cordic/mycordic/n586 ), .B(n95), .S(
        n766), .Q(\u_cordic/mycordic/n585 ) );
  MUX22 \u_cordic/mycordic/U554  ( .A(
        \u_cordic/mycordic/present_ANGLE_table[6][15] ), .B(
        \u_cordic/mycordic/n585 ), .S(n384), .Q(
        \u_cordic/mycordic/next_ANGLE_table[6][15] ) );
  IMUX21 \u_cordic/mycordic/U549  ( .A(\u_cordic/mycordic/n582 ), .B(n375), 
        .S(n766), .Q(\u_cordic/mycordic/n581 ) );
  MUX22 \u_cordic/mycordic/U550  ( .A(
        \u_cordic/mycordic/present_ANGLE_table[6][13] ), .B(
        \u_cordic/mycordic/n581 ), .S(n384), .Q(
        \u_cordic/mycordic/next_ANGLE_table[6][13] ) );
  XOR31 \u_cordic/mycordic/sub_194/U2_7  ( .A(
        \u_cordic/mycordic/present_I_table[2][7] ), .B(n287), .C(
        \u_cordic/mycordic/sub_194/carry [7]), .Q(\u_cordic/mycordic/N355 ) );
  XOR31 \u_cordic/mycordic/add_189/U1_7  ( .A(
        \u_cordic/mycordic/present_I_table[2][7] ), .B(
        \u_cordic/mycordic/present_Q_table[2][7] ), .C(
        \u_cordic/mycordic/add_189/carry [7]), .Q(\u_cordic/mycordic/N323 ) );
  XOR31 \u_cordic/mycordic/sub_205/U2_7  ( .A(
        \u_cordic/mycordic/present_I_table[3][7] ), .B(n245), .C(
        \u_cordic/mycordic/sub_205/carry [7]), .Q(\u_cordic/mycordic/N419 ) );
  XOR31 \u_cordic/mycordic/add_200/U1_7  ( .A(
        \u_cordic/mycordic/present_I_table[3][7] ), .B(
        \u_cordic/mycordic/present_Q_table[3][7] ), .C(
        \u_cordic/mycordic/add_200/carry [7]), .Q(\u_cordic/mycordic/N387 ) );
  IMUX21 \u_cordic/mycordic/U551  ( .A(\u_cordic/mycordic/n584 ), .B(n374), 
        .S(n766), .Q(\u_cordic/mycordic/n583 ) );
  MUX22 \u_cordic/mycordic/U552  ( .A(
        \u_cordic/mycordic/present_ANGLE_table[6][14] ), .B(
        \u_cordic/mycordic/n583 ), .S(n384), .Q(
        \u_cordic/mycordic/next_ANGLE_table[6][14] ) );
  NAND22 \u_cordic/mycordic/U571  ( .A(\u_cordic/mycordic/N629 ), .B(n758), 
        .Q(\u_cordic/mycordic/n584 ) );
  NAND22 \u_cordic/mycordic/U572  ( .A(\u_cordic/mycordic/N630 ), .B(n757), 
        .Q(\u_cordic/mycordic/n586 ) );
  XOR31 \u_cordic/mycordic/sub_223/U2_7  ( .A(
        \u_cordic/mycordic/present_Q_table[5][7] ), .B(n199), .C(
        \u_cordic/mycordic/sub_223/carry[7] ), .Q(\u_cordic/mycordic/N500 ) );
  XOR31 \u_cordic/mycordic/add_228/U1_7  ( .A(
        \u_cordic/mycordic/present_Q_table[5][7] ), .B(
        \u_cordic/mycordic/present_I_table[5][7] ), .C(
        \u_cordic/mycordic/add_228/carry[7] ), .Q(\u_cordic/mycordic/N517 ) );
  XOR31 \u_cordic/mycordic/sub_212/U2_7  ( .A(
        \u_cordic/mycordic/present_Q_table[4][7] ), .B(n47), .C(
        \u_cordic/mycordic/sub_212/carry [7]), .Q(\u_cordic/mycordic/N455 ) );
  XOR31 \u_cordic/mycordic/add_217/U1_7  ( .A(
        \u_cordic/mycordic/present_Q_table[4][7] ), .B(
        \u_cordic/mycordic/present_I_table[4][7] ), .C(
        \u_cordic/mycordic/add_217/carry [7]), .Q(\u_cordic/mycordic/N483 ) );
  XOR31 \u_cordic/mycordic/add_211/U1_7  ( .A(
        \u_cordic/mycordic/present_I_table[4][7] ), .B(
        \u_cordic/mycordic/present_Q_table[4][7] ), .C(
        \u_cordic/mycordic/add_211/carry [7]), .Q(\u_cordic/mycordic/N447 ) );
  XOR31 \u_cordic/mycordic/sub_216/U2_7  ( .A(
        \u_cordic/mycordic/present_I_table[4][7] ), .B(n48), .C(
        \u_cordic/mycordic/sub_216/carry [7]), .Q(\u_cordic/mycordic/N475 ) );
  XOR31 \u_cordic/mycordic/sub_190/U2_7  ( .A(
        \u_cordic/mycordic/present_Q_table[2][7] ), .B(n288), .C(
        \u_cordic/mycordic/sub_190/carry [7]), .Q(\u_cordic/mycordic/N331 ) );
  XOR31 \u_cordic/mycordic/add_195/U1_7  ( .A(
        \u_cordic/mycordic/present_Q_table[2][7] ), .B(
        \u_cordic/mycordic/present_I_table[2][7] ), .C(
        \u_cordic/mycordic/add_195/carry [7]), .Q(\u_cordic/mycordic/N363 ) );
  XOR31 \u_cordic/mycordic/sub_201/U2_7  ( .A(
        \u_cordic/mycordic/present_Q_table[3][7] ), .B(n246), .C(
        \u_cordic/mycordic/sub_201/carry [7]), .Q(\u_cordic/mycordic/N395 ) );
  XOR31 \u_cordic/mycordic/add_206/U1_7  ( .A(
        \u_cordic/mycordic/present_Q_table[3][7] ), .B(
        \u_cordic/mycordic/present_I_table[3][7] ), .C(
        \u_cordic/mycordic/add_206/carry [7]), .Q(\u_cordic/mycordic/N427 ) );
  XOR31 \u_decoder/fir_filter/add_326/U1_14  ( .A(
        \u_decoder/fir_filter/Q_data_mult_0_buff [14]), .B(
        \u_decoder/fir_filter/Q_data_add_1_buff [14]), .C(
        \u_decoder/fir_filter/add_326/carry [14]), .Q(
        \u_decoder/fir_filter/Q_data_add_0 [14]) );
  XOR31 \u_decoder/fir_filter/add_327/U1_14  ( .A(
        \u_decoder/fir_filter/Q_data_mult_1_buff [14]), .B(
        \u_decoder/fir_filter/Q_data_add_2_buff [14]), .C(
        \u_decoder/fir_filter/add_327/carry [14]), .Q(
        \u_decoder/fir_filter/Q_data_add_1 [14]) );
  XOR31 \u_decoder/fir_filter/add_328/U1_14  ( .A(
        \u_decoder/fir_filter/Q_data_mult_2_buff [14]), .B(
        \u_decoder/fir_filter/Q_data_add_3_buff [14]), .C(
        \u_decoder/fir_filter/add_328/carry [14]), .Q(
        \u_decoder/fir_filter/Q_data_add_2 [14]) );
  XOR31 \u_decoder/fir_filter/add_329/U1_14  ( .A(
        \u_decoder/fir_filter/Q_data_mult_3_buff [14]), .B(
        \u_decoder/fir_filter/Q_data_add_4_buff [14]), .C(
        \u_decoder/fir_filter/add_329/carry [14]), .Q(
        \u_decoder/fir_filter/Q_data_add_3 [14]) );
  XOR31 \u_decoder/fir_filter/add_331/U1_14  ( .A(
        \u_decoder/fir_filter/Q_data_mult_5_buff [14]), .B(
        \u_decoder/fir_filter/Q_data_add_6_buff [14]), .C(
        \u_decoder/fir_filter/add_331/carry [14]), .Q(
        \u_decoder/fir_filter/Q_data_add_5 [14]) );
  XOR31 \u_decoder/fir_filter/add_332/U1_14  ( .A(
        \u_decoder/fir_filter/Q_data_mult_6_buff [14]), .B(
        \u_decoder/fir_filter/Q_data_add_7_buff [14]), .C(
        \u_decoder/fir_filter/add_332/carry [14]), .Q(
        \u_decoder/fir_filter/Q_data_add_6 [14]) );
  XOR31 \u_decoder/fir_filter/add_333/U1_14  ( .A(
        \u_decoder/fir_filter/Q_data_mult_7_buff [14]), .B(
        \u_decoder/fir_filter/Q_data_mult_8_buff [14]), .C(
        \u_decoder/fir_filter/add_333/carry [14]), .Q(
        \u_decoder/fir_filter/Q_data_add_7 [14]) );
  XOR31 \u_decoder/fir_filter/add_294/U1_14  ( .A(
        \u_decoder/fir_filter/I_data_mult_0_buff [14]), .B(
        \u_decoder/fir_filter/I_data_add_1_buff [14]), .C(
        \u_decoder/fir_filter/add_294/carry [14]), .Q(
        \u_decoder/fir_filter/I_data_add_0 [14]) );
  XOR31 \u_decoder/fir_filter/add_295/U1_14  ( .A(
        \u_decoder/fir_filter/I_data_mult_1_buff [14]), .B(
        \u_decoder/fir_filter/I_data_add_2_buff [14]), .C(
        \u_decoder/fir_filter/add_295/carry [14]), .Q(
        \u_decoder/fir_filter/I_data_add_1 [14]) );
  XOR31 \u_decoder/fir_filter/add_296/U1_14  ( .A(
        \u_decoder/fir_filter/I_data_mult_2_buff [14]), .B(
        \u_decoder/fir_filter/I_data_add_3_buff [14]), .C(
        \u_decoder/fir_filter/add_296/carry [14]), .Q(
        \u_decoder/fir_filter/I_data_add_2 [14]) );
  XOR31 \u_decoder/fir_filter/add_297/U1_14  ( .A(
        \u_decoder/fir_filter/I_data_mult_3_buff [14]), .B(
        \u_decoder/fir_filter/I_data_add_4_buff [14]), .C(
        \u_decoder/fir_filter/add_297/carry [14]), .Q(
        \u_decoder/fir_filter/I_data_add_3 [14]) );
  XOR31 \u_decoder/fir_filter/add_299/U1_14  ( .A(
        \u_decoder/fir_filter/I_data_mult_5_buff [14]), .B(
        \u_decoder/fir_filter/I_data_add_6_buff [14]), .C(
        \u_decoder/fir_filter/add_299/carry [14]), .Q(
        \u_decoder/fir_filter/I_data_add_5 [14]) );
  XOR31 \u_decoder/fir_filter/add_300/U1_14  ( .A(
        \u_decoder/fir_filter/I_data_mult_6_buff [14]), .B(
        \u_decoder/fir_filter/I_data_add_7_buff [14]), .C(
        \u_decoder/fir_filter/add_300/carry [14]), .Q(
        \u_decoder/fir_filter/I_data_add_6 [14]) );
  XOR31 \u_decoder/fir_filter/add_301/U1_14  ( .A(
        \u_decoder/fir_filter/I_data_mult_7_buff [14]), .B(
        \u_decoder/fir_filter/I_data_mult_8_buff [14]), .C(
        \u_decoder/fir_filter/add_301/carry [14]), .Q(
        \u_decoder/fir_filter/I_data_add_7 [14]) );
  XOR31 \u_decoder/fir_filter/add_330/U1_14  ( .A(
        \u_decoder/fir_filter/Q_data_mult_4_buff [14]), .B(
        \u_decoder/fir_filter/Q_data_add_5_buff [14]), .C(
        \u_decoder/fir_filter/add_330/carry [14]), .Q(
        \u_decoder/fir_filter/Q_data_add_4 [14]) );
  XOR31 \u_decoder/fir_filter/add_298/U1_14  ( .A(
        \u_decoder/fir_filter/I_data_mult_4_buff [14]), .B(
        \u_decoder/fir_filter/I_data_add_5_buff [14]), .C(
        \u_decoder/fir_filter/add_298/carry [14]), .Q(
        \u_decoder/fir_filter/I_data_add_4 [14]) );
  XOR31 \u_cordic/my_rotation/sub_35/U2_15  ( .A(
        \u_cordic/my_rotation/present_angle[0][15] ), .B(n193), .C(
        \u_cordic/my_rotation/sub_35/carry [15]), .Q(
        \u_cordic/my_rotation/N23 ) );
  IMUX40 \u_inFIFO/U585  ( .A(\u_inFIFO/n716 ), .B(\u_inFIFO/n717 ), .C(
        \u_inFIFO/n718 ), .D(\u_inFIFO/n719 ), .S0(\u_inFIFO/N40 ), .S1(n15), 
        .Q(\u_inFIFO/n715 ) );
  IMUX40 \u_inFIFO/U587  ( .A(\u_inFIFO/n726 ), .B(\u_inFIFO/n727 ), .C(
        \u_inFIFO/n728 ), .D(\u_inFIFO/n729 ), .S0(\u_inFIFO/N40 ), .S1(n15), 
        .Q(\u_inFIFO/n725 ) );
  IMUX40 \u_inFIFO/U586  ( .A(\u_inFIFO/n721 ), .B(\u_inFIFO/n722 ), .C(
        \u_inFIFO/n723 ), .D(\u_inFIFO/n724 ), .S0(\u_inFIFO/N40 ), .S1(n15), 
        .Q(\u_inFIFO/n720 ) );
  IMUX40 \u_inFIFO/U711  ( .A(\u_inFIFO/n725 ), .B(\u_inFIFO/n715 ), .C(
        \u_inFIFO/n720 ), .D(\u_inFIFO/n710 ), .S0(n49), .S1(n765), .Q(
        \u_inFIFO/n751 ) );
  IMUX40 \u_inFIFO/U589  ( .A(\u_inFIFO/n736 ), .B(\u_inFIFO/n737 ), .C(
        \u_inFIFO/n738 ), .D(\u_inFIFO/n739 ), .S0(\u_inFIFO/N40 ), .S1(n15), 
        .Q(\u_inFIFO/n735 ) );
  IMUX40 \u_inFIFO/U588  ( .A(\u_inFIFO/n731 ), .B(\u_inFIFO/n732 ), .C(
        \u_inFIFO/n733 ), .D(\u_inFIFO/n734 ), .S0(\u_inFIFO/N40 ), .S1(n15), 
        .Q(\u_inFIFO/n730 ) );
  IMUX40 \u_inFIFO/U590  ( .A(\u_inFIFO/n741 ), .B(\u_inFIFO/n742 ), .C(
        \u_inFIFO/n743 ), .D(\u_inFIFO/n744 ), .S0(\u_inFIFO/N40 ), .S1(n15), 
        .Q(\u_inFIFO/n740 ) );
  IMUX40 \u_inFIFO/U728  ( .A(\u_inFIFO/n745 ), .B(\u_inFIFO/n735 ), .C(
        \u_inFIFO/n740 ), .D(\u_inFIFO/n730 ), .S0(n49), .S1(n765), .Q(
        \u_inFIFO/n750 ) );
  XOR31 \u_decoder/iq_demod/dp_cluster_0/sub_153/U2_7  ( .A(
        \u_decoder/iq_demod/dp_cluster_0/mult_I_cos_out [7]), .B(n350), .C(
        \u_decoder/iq_demod/dp_cluster_0/sub_153/carry [7]), .Q(
        \u_decoder/iq_demod/add_I_out [7]) );
  XOR31 \u_decoder/iq_demod/dp_cluster_1/add_154/U1_7  ( .A(
        \u_decoder/iq_demod/dp_cluster_1/mult_I_sin_out [7]), .B(
        \u_decoder/iq_demod/dp_cluster_1/mult_Q_cos_out [7]), .C(
        \u_decoder/iq_demod/dp_cluster_1/add_154/carry [7]), .Q(
        \u_decoder/iq_demod/add_Q_out [7]) );
  IMUX21 \u_inFIFO/U592  ( .A(\u_inFIFO/n750 ), .B(\u_inFIFO/n751 ), .S(
        \u_inFIFO/N43 ), .Q(\u_inFIFO/N200 ) );
  ADD32 \u_cordic/mycordic/r144/U1_3  ( .A(
        \u_cordic/mycordic/present_I_table[1][3] ), .B(
        \u_cordic/mycordic/present_Q_table[1][3] ), .CI(n2), .CO(
        \u_cordic/mycordic/r144/carry [4]), .S(\u_cordic/mycordic/N255 ) );
  ADD32 \u_cordic/mycordic/sub_182/U2_3  ( .A(
        \u_cordic/mycordic/present_I_table[1][3] ), .B(n216), .CI(n1), .CO(
        \u_cordic/mycordic/sub_182/carry [4]), .S(\u_cordic/mycordic/N287 ) );
  ADD32 \u_cordic/mycordic/sub_178/U2_3  ( .A(
        \u_cordic/mycordic/present_Q_table[1][3] ), .B(n215), .CI(n1), .CO(
        \u_cordic/mycordic/sub_178/carry [4]), .S(\u_cordic/mycordic/N263 ) );
  LOGIC1 U2 ( .Q(n1) );
  LOGIC0 U3 ( .Q(n2) );
  NOR21 U4 ( .A(n692), .B(n693), .Q(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/A2[5] ) );
  INV3 U5 ( .A(\u_cordic/mycordic/n353 ), .Q(n1436) );
  INV3 U6 ( .A(\u_decoder/fir_filter/n1084 ), .Q(n2259) );
  INV3 U7 ( .A(\u_decoder/fir_filter/n787 ), .Q(n2330) );
  NOR21 U8 ( .A(\u_coder/n315 ), .B(n373), .Q(\u_coder/N522 ) );
  INV2 U9 ( .A(\u_inFIFO/n225 ), .Q(n1211) );
  CLKIN3 U10 ( .A(n1211), .Q(n1210) );
  XNR21 U11 ( .A(n303), .B(\u_cordic/mycordic/sub_add_150_b0/carry [7]), .Q(
        n51) );
  XOR21 U12 ( .A(\u_cdr/phd1/cnt_phd/cnt [1]), .B(n1363), .Q(n61) );
  XNR21 U13 ( .A(n1195), .B(n2347), .Q(n67) );
  XNR21 U14 ( .A(n1193), .B(n2276), .Q(n68) );
  XNR21 U15 ( .A(n2854), .B(n2855), .Q(n69) );
  XNR21 U16 ( .A(n2940), .B(n2941), .Q(n70) );
  XOR21 U17 ( .A(n2835), .B(n2836), .Q(n76) );
  XOR21 U18 ( .A(n2921), .B(n2922), .Q(n77) );
  XNR31 U19 ( .A(\u_decoder/fir_filter/dp_cluster_0/r177/A2[7] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r177/A1[7] ), .C(n2795), .Q(n78) );
  XNR31 U20 ( .A(\u_decoder/fir_filter/dp_cluster_0/r164/A2[7] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r164/A1[7] ), .C(n2881), .Q(n79) );
  XOR21 U21 ( .A(n2791), .B(n2792), .Q(n82) );
  XOR21 U22 ( .A(\u_decoder/iq_demod/dp_cluster_0/mult_151/A1[2] ), .B(n2386), 
        .Q(n83) );
  XNR21 U23 ( .A(\u_cordic/mycordic/present_ANGLE_table[6][15] ), .B(
        \u_cordic/mycordic/r173/carry [15]), .Q(n95) );
  XNR21 U24 ( .A(n2814), .B(n2815), .Q(n127) );
  XNR21 U25 ( .A(n2900), .B(n2901), .Q(n128) );
  XOR21 U26 ( .A(n2365), .B(n2803), .Q(n131) );
  XOR21 U27 ( .A(n2294), .B(n2889), .Q(n132) );
  XNR21 U28 ( .A(\u_decoder/iq_demod/dp_cluster_0/mult_151/ab[0][1] ), .B(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/ab[1][0] ), .Q(n170) );
  NOR21 U29 ( .A(n1237), .B(\u_outFIFO/n1117 ), .Q(\u_outFIFO/n660 ) );
  AOI221 U30 ( .A(\u_decoder/fir_filter/I_data_mult_4 [14]), .B(n1083), .C(
        \u_decoder/fir_filter/I_data_mult_4_buff [14]), .D(n1162), .Q(
        \u_decoder/fir_filter/n1084 ) );
  AOI221 U31 ( .A(\u_decoder/fir_filter/Q_data_mult_4 [14]), .B(n1083), .C(
        \u_decoder/fir_filter/Q_data_mult_4_buff [14]), .D(n1160), .Q(
        \u_decoder/fir_filter/n787 ) );
  BUF2 U32 ( .A(\u_decoder/I_prefilter [7]), .Q(n1193) );
  BUF2 U33 ( .A(\u_decoder/Q_prefilter [7]), .Q(n1195) );
  BUF2 U34 ( .A(\u_decoder/I_prefilter [7]), .Q(n1192) );
  BUF2 U35 ( .A(\u_decoder/Q_prefilter [7]), .Q(n1194) );
  NOR21 U36 ( .A(\u_outFIFO/n285 ), .B(\u_outFIFO/k_FIFO [1]), .Q(
        \u_outFIFO/n666 ) );
  NOR21 U37 ( .A(\u_outFIFO/n284 ), .B(\u_outFIFO/k_FIFO [0]), .Q(
        \u_outFIFO/n664 ) );
  NOR21 U38 ( .A(\u_outFIFO/i_FIFO [3]), .B(\u_outFIFO/i_FIFO [2]), .Q(
        \u_outFIFO/n983 ) );
  AOI221 U39 ( .A(n1901), .B(\u_cordic/mycordic/N247 ), .C(
        \u_cordic/mycordic/n354 ), .D(
        \u_cordic/mycordic/present_Q_table[0][7] ), .Q(
        \u_cordic/mycordic/n353 ) );
  INV3 U40 ( .A(\u_cordic/mycordic/n520 ), .Q(n1904) );
  INV3 U41 ( .A(n1103), .Q(n1083) );
  INV3 U42 ( .A(n1100), .Q(n1091) );
  INV3 U43 ( .A(n1100), .Q(n1092) );
  INV3 U44 ( .A(n1099), .Q(n1093) );
  INV3 U45 ( .A(n1099), .Q(n1094) );
  INV3 U46 ( .A(n1099), .Q(n1095) );
  INV3 U47 ( .A(n1102), .Q(n1084) );
  INV3 U48 ( .A(n1102), .Q(n1085) );
  INV3 U49 ( .A(n1102), .Q(n1086) );
  INV3 U50 ( .A(n1101), .Q(n1087) );
  INV3 U51 ( .A(n1101), .Q(n1088) );
  INV3 U52 ( .A(n1101), .Q(n1089) );
  INV3 U53 ( .A(n1100), .Q(n1090) );
  INV3 U54 ( .A(n1098), .Q(n1096) );
  INV3 U55 ( .A(n1098), .Q(n1097) );
  BUF2 U56 ( .A(n913), .Q(n926) );
  BUF2 U57 ( .A(n925), .Q(n951) );
  BUF2 U58 ( .A(n925), .Q(n950) );
  BUF2 U59 ( .A(n924), .Q(n949) );
  BUF2 U60 ( .A(n924), .Q(n948) );
  BUF2 U61 ( .A(n923), .Q(n947) );
  BUF2 U62 ( .A(n923), .Q(n946) );
  BUF2 U63 ( .A(n922), .Q(n945) );
  BUF2 U64 ( .A(n922), .Q(n944) );
  BUF2 U65 ( .A(n921), .Q(n943) );
  BUF2 U66 ( .A(n921), .Q(n942) );
  BUF2 U67 ( .A(n920), .Q(n941) );
  BUF2 U68 ( .A(n920), .Q(n940) );
  BUF2 U69 ( .A(n919), .Q(n939) );
  BUF2 U70 ( .A(n919), .Q(n938) );
  BUF2 U71 ( .A(n918), .Q(n937) );
  BUF2 U72 ( .A(n918), .Q(n936) );
  BUF2 U73 ( .A(n917), .Q(n935) );
  BUF2 U74 ( .A(n917), .Q(n934) );
  BUF2 U75 ( .A(n916), .Q(n933) );
  BUF2 U76 ( .A(n916), .Q(n932) );
  BUF2 U77 ( .A(n915), .Q(n931) );
  BUF2 U78 ( .A(n915), .Q(n930) );
  BUF2 U79 ( .A(n914), .Q(n929) );
  BUF2 U80 ( .A(n914), .Q(n928) );
  BUF2 U81 ( .A(n913), .Q(n927) );
  AOI211 U82 ( .A(n2921), .B(n2278), .C(n2280), .Q(n2940) );
  INV3 U83 ( .A(n2923), .Q(n2280) );
  AOI211 U84 ( .A(n2835), .B(n2349), .C(n2351), .Q(n2854) );
  INV3 U85 ( .A(n2837), .Q(n2351) );
  AOI211 U86 ( .A(n2943), .B(n2262), .C(n2264), .Q(n2962) );
  INV3 U87 ( .A(n2945), .Q(n2264) );
  AOI211 U88 ( .A(n2857), .B(n2333), .C(n2335), .Q(n2876) );
  INV3 U89 ( .A(n2859), .Q(n2335) );
  INV3 U90 ( .A(n2960), .Q(n2263) );
  INV3 U91 ( .A(n2874), .Q(n2334) );
  INV3 U92 ( .A(n2924), .Q(n2282) );
  INV3 U93 ( .A(n2838), .Q(n2353) );
  XNR21 U94 ( .A(\u_decoder/fir_filter/dp_cluster_0/r167/SUMB[7][1] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[7][0] ), .Q(n321) );
  XNR21 U95 ( .A(\u_decoder/fir_filter/dp_cluster_0/r180/SUMB[7][1] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[7][0] ), .Q(n322) );
  NAND22 U96 ( .A(n2275), .B(n2937), .Q(n2941) );
  INV3 U97 ( .A(n2934), .Q(n2275) );
  NAND22 U98 ( .A(n2346), .B(n2851), .Q(n2855) );
  INV3 U99 ( .A(n2848), .Q(n2346) );
  NAND22 U100 ( .A(n2278), .B(n2923), .Q(n2922) );
  NAND22 U101 ( .A(n2349), .B(n2837), .Q(n2836) );
  NOR21 U102 ( .A(n586), .B(n587), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r167/A2[7] ) );
  INV3 U103 ( .A(\u_decoder/fir_filter/dp_cluster_0/r167/SUMB[7][1] ), .Q(n587) );
  INV3 U104 ( .A(\u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[7][0] ), .Q(
        n586) );
  NOR21 U105 ( .A(n647), .B(n648), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r180/A2[7] ) );
  INV3 U106 ( .A(\u_decoder/fir_filter/dp_cluster_0/r180/SUMB[7][1] ), .Q(n648) );
  INV3 U107 ( .A(\u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[7][0] ), .Q(
        n647) );
  INV3 U108 ( .A(n2938), .Q(n2279) );
  INV3 U109 ( .A(n2852), .Q(n2350) );
  INV3 U110 ( .A(n2955), .Q(n2262) );
  INV3 U111 ( .A(n2869), .Q(n2333) );
  INV3 U112 ( .A(n2956), .Q(n2257) );
  INV3 U113 ( .A(n2870), .Q(n2328) );
  INV3 U114 ( .A(n2933), .Q(n2278) );
  INV3 U115 ( .A(n2847), .Q(n2349) );
  BUF2 U116 ( .A(n1141), .Q(n1099) );
  BUF2 U117 ( .A(n1144), .Q(n1102) );
  BUF2 U118 ( .A(n1142), .Q(n1101) );
  BUF2 U119 ( .A(n1139), .Q(n1100) );
  BUF2 U120 ( .A(n1144), .Q(n1103) );
  BUF2 U121 ( .A(n1138), .Q(n1098) );
  BUF2 U122 ( .A(n1143), .Q(n1105) );
  BUF2 U123 ( .A(n1143), .Q(n1104) );
  BUF2 U124 ( .A(n1143), .Q(n1106) );
  BUF2 U125 ( .A(n1140), .Q(n1122) );
  BUF2 U126 ( .A(n1140), .Q(n1123) );
  BUF2 U127 ( .A(n1140), .Q(n1124) );
  BUF2 U128 ( .A(n1140), .Q(n1125) );
  BUF2 U129 ( .A(n1140), .Q(n1126) );
  BUF2 U130 ( .A(n1140), .Q(n1127) );
  BUF2 U131 ( .A(n1139), .Q(n1128) );
  BUF2 U132 ( .A(n1139), .Q(n1129) );
  BUF2 U133 ( .A(n1139), .Q(n1130) );
  BUF2 U134 ( .A(n1139), .Q(n1131) );
  BUF2 U135 ( .A(n1139), .Q(n1132) );
  BUF2 U136 ( .A(n1139), .Q(n1133) );
  BUF2 U137 ( .A(n1142), .Q(n1107) );
  BUF2 U138 ( .A(n1143), .Q(n1108) );
  BUF2 U139 ( .A(n1143), .Q(n1109) );
  BUF2 U140 ( .A(n1142), .Q(n1110) );
  BUF2 U141 ( .A(n1142), .Q(n1111) );
  BUF2 U142 ( .A(n1142), .Q(n1112) );
  BUF2 U143 ( .A(n1142), .Q(n1113) );
  BUF2 U144 ( .A(n1142), .Q(n1114) );
  BUF2 U145 ( .A(n1141), .Q(n1115) );
  BUF2 U146 ( .A(n1141), .Q(n1116) );
  BUF2 U147 ( .A(n1141), .Q(n1117) );
  BUF2 U148 ( .A(n1141), .Q(n1118) );
  BUF2 U149 ( .A(n1141), .Q(n1119) );
  BUF2 U150 ( .A(n1141), .Q(n1120) );
  BUF2 U151 ( .A(n1141), .Q(n1121) );
  BUF2 U152 ( .A(n1138), .Q(n1134) );
  BUF2 U153 ( .A(n1138), .Q(n1135) );
  BUF2 U154 ( .A(n1138), .Q(n1136) );
  BUF2 U155 ( .A(n1794), .Q(n925) );
  BUF2 U156 ( .A(n1794), .Q(n924) );
  BUF2 U157 ( .A(n1794), .Q(n923) );
  BUF2 U158 ( .A(n1794), .Q(n922) );
  BUF2 U159 ( .A(n1794), .Q(n921) );
  BUF2 U160 ( .A(n1794), .Q(n920) );
  BUF2 U161 ( .A(n1794), .Q(n919) );
  BUF2 U162 ( .A(n1794), .Q(n918) );
  BUF2 U163 ( .A(n1794), .Q(n917) );
  BUF2 U164 ( .A(n1794), .Q(n916) );
  BUF2 U165 ( .A(n1794), .Q(n915) );
  BUF2 U166 ( .A(n1794), .Q(n914) );
  BUF2 U167 ( .A(n1794), .Q(n913) );
  BUF2 U168 ( .A(n1138), .Q(n1137) );
  NAND31 U169 ( .A(n1378), .B(n1291), .C(n1379), .Q(n1295) );
  INV3 U170 ( .A(n2898), .Q(n2241) );
  INV3 U171 ( .A(n2812), .Q(n2312) );
  AOI211 U172 ( .A(n2899), .B(\u_decoder/fir_filter/dp_cluster_0/r165/A1[7] ), 
        .C(n2242), .Q(n2898) );
  INV3 U173 ( .A(n2910), .Q(n2242) );
  AOI211 U174 ( .A(n2813), .B(\u_decoder/fir_filter/dp_cluster_0/r178/A1[7] ), 
        .C(n2313), .Q(n2812) );
  INV3 U175 ( .A(n2824), .Q(n2313) );
  NOR21 U176 ( .A(\u_decoder/fir_filter/dp_cluster_0/r167/A1[8] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r167/A2[8] ), .Q(n2942) );
  NOR21 U177 ( .A(\u_decoder/fir_filter/dp_cluster_0/r180/A1[8] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r180/A2[8] ), .Q(n2856) );
  NOR21 U178 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_276/A1[8] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/A2[8] ), .Q(n2964) );
  NOR21 U179 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_308/A1[8] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/A2[8] ), .Q(n2878) );
  INV3 U180 ( .A(n2880), .Q(n2290) );
  INV3 U181 ( .A(n2794), .Q(n2361) );
  INV3 U182 ( .A(\u_decoder/fir_filter/dp_cluster_0/r165/A1[9] ), .Q(n2238) );
  INV3 U183 ( .A(n2897), .Q(n2239) );
  INV3 U184 ( .A(\u_decoder/fir_filter/dp_cluster_0/r178/A1[9] ), .Q(n2309) );
  INV3 U185 ( .A(n2811), .Q(n2310) );
  XOR21 U186 ( .A(\u_decoder/fir_filter/dp_cluster_0/r167/SUMB[6][1] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[6][0] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r167/SUMB[7][0] ) );
  XOR21 U187 ( .A(\u_decoder/fir_filter/dp_cluster_0/r180/SUMB[6][1] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[6][0] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r180/SUMB[7][0] ) );
  XOR21 U188 ( .A(\u_decoder/fir_filter/dp_cluster_0/r164/SUMB[5][2] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r164/CARRYB[6][0] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r164/SUMB[7][0] ) );
  XOR21 U189 ( .A(\u_decoder/fir_filter/dp_cluster_0/r177/SUMB[5][2] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r177/CARRYB[6][0] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r177/SUMB[7][0] ) );
  XOR21 U190 ( .A(\u_decoder/fir_filter/dp_cluster_0/r165/SUMB[4][3] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r165/CARRYB[6][0] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r165/SUMB[7][0] ) );
  XOR21 U191 ( .A(\u_decoder/fir_filter/dp_cluster_0/r178/SUMB[4][3] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r178/CARRYB[6][0] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r178/SUMB[7][0] ) );
  XOR21 U192 ( .A(\u_decoder/fir_filter/dp_cluster_0/r166/SUMB[5][3] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r166/CARRYB[6][1] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r166/SUMB[7][1] ) );
  XOR21 U193 ( .A(\u_decoder/fir_filter/dp_cluster_0/r179/SUMB[5][3] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r179/CARRYB[6][1] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r179/SUMB[7][1] ) );
  XOR21 U194 ( .A(\u_decoder/fir_filter/dp_cluster_0/r167/SUMB[5][3] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[6][1] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r167/SUMB[7][1] ) );
  XOR21 U195 ( .A(\u_decoder/fir_filter/dp_cluster_0/r180/SUMB[5][3] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[6][1] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r180/SUMB[7][1] ) );
  XOR21 U196 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_276/SUMB[5][5] ), 
        .B(\u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[6][3] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/SUMB[7][3] ) );
  XOR21 U197 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_308/SUMB[5][5] ), 
        .B(\u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[6][3] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/SUMB[7][3] ) );
  XNR31 U198 ( .A(\u_decoder/fir_filter/dp_cluster_0/r166/A2[9] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r166/CARRYB[7][3] ), .C(n2912), .Q(
        n323) );
  XNR31 U199 ( .A(\u_decoder/fir_filter/dp_cluster_0/r165/A2[10] ), .B(n2305), 
        .C(n2906), .Q(n324) );
  XNR31 U200 ( .A(\u_decoder/fir_filter/dp_cluster_0/r164/A2[9] ), .B(n2305), 
        .C(n2879), .Q(n325) );
  XNR31 U201 ( .A(\u_decoder/fir_filter/dp_cluster_0/r179/A2[9] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r179/CARRYB[7][3] ), .C(n2826), .Q(
        n326) );
  XNR31 U202 ( .A(\u_decoder/fir_filter/dp_cluster_0/r178/A2[10] ), .B(n2376), 
        .C(n2820), .Q(n327) );
  XNR31 U203 ( .A(\u_decoder/fir_filter/dp_cluster_0/r177/A2[9] ), .B(n2376), 
        .C(n2793), .Q(n328) );
  XOR21 U204 ( .A(n16), .B(
        \u_decoder/fir_filter/dp_cluster_0/r164/CARRYB[6][2] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r164/SUMB[7][2] ) );
  XOR21 U205 ( .A(n17), .B(
        \u_decoder/fir_filter/dp_cluster_0/r177/CARRYB[6][2] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r177/SUMB[7][2] ) );
  INV3 U206 ( .A(\u_decoder/fir_filter/dp_cluster_0/r166/CARRYB[7][3] ), .Q(
        n2245) );
  INV3 U207 ( .A(n2912), .Q(n2246) );
  INV3 U208 ( .A(\u_decoder/fir_filter/dp_cluster_0/r179/CARRYB[7][3] ), .Q(
        n2316) );
  INV3 U209 ( .A(n2826), .Q(n2317) );
  AOI2111 U210 ( .A(n2953), .B(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[7][5] ), .C(n2260), 
        .D(n2954), .Q(n2952) );
  INV3 U211 ( .A(n2958), .Q(n2260) );
  NOR40 U212 ( .A(n2955), .B(n2946), .C(n2956), .D(n2957), .Q(n2954) );
  AOI2111 U213 ( .A(n2867), .B(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[7][5] ), .C(n2331), 
        .D(n2868), .Q(n2866) );
  INV3 U214 ( .A(n2872), .Q(n2331) );
  NOR40 U215 ( .A(n2869), .B(n2860), .C(n2870), .D(n2871), .Q(n2868) );
  NAND22 U216 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_276/A2[9] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/A1[9] ), .Q(n2945) );
  NAND22 U217 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_308/A2[9] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/A1[9] ), .Q(n2859) );
  NOR21 U218 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_276/A2[9] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/A1[9] ), .Q(n2955) );
  NOR21 U219 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_308/A2[9] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/A1[9] ), .Q(n2869) );
  NAND22 U220 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_276/A2[8] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/A1[8] ), .Q(n2947) );
  NAND22 U221 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_308/A2[8] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/A1[8] ), .Q(n2861) );
  XNR21 U222 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_276/A1[8] ), .B(
        n2946), .Q(n2949) );
  XNR21 U223 ( .A(\u_decoder/fir_filter/dp_cluster_0/r167/A1[8] ), .B(n2924), 
        .Q(n2927) );
  XNR21 U224 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_308/A1[8] ), .B(
        n2860), .Q(n2863) );
  XNR21 U225 ( .A(\u_decoder/fir_filter/dp_cluster_0/r180/A1[8] ), .B(n2838), 
        .Q(n2841) );
  INV3 U226 ( .A(n2913), .Q(n2248) );
  INV3 U227 ( .A(n2827), .Q(n2319) );
  NOR21 U228 ( .A(n606), .B(n607), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r165/CARRYB[7][0] ) );
  INV3 U229 ( .A(\u_decoder/fir_filter/dp_cluster_0/r165/SUMB[4][3] ), .Q(n606) );
  INV3 U230 ( .A(\u_decoder/fir_filter/dp_cluster_0/r165/CARRYB[6][0] ), .Q(
        n607) );
  NOR21 U231 ( .A(n667), .B(n668), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r178/CARRYB[7][0] ) );
  INV3 U232 ( .A(\u_decoder/fir_filter/dp_cluster_0/r178/SUMB[4][3] ), .Q(n667) );
  INV3 U233 ( .A(\u_decoder/fir_filter/dp_cluster_0/r178/CARRYB[6][0] ), .Q(
        n668) );
  NOR21 U234 ( .A(n596), .B(n597), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r166/CARRYB[7][1] ) );
  INV3 U235 ( .A(\u_decoder/fir_filter/dp_cluster_0/r166/CARRYB[6][1] ), .Q(
        n597) );
  INV3 U236 ( .A(\u_decoder/fir_filter/dp_cluster_0/r166/SUMB[5][3] ), .Q(n596) );
  NOR21 U237 ( .A(n657), .B(n658), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r179/CARRYB[7][1] ) );
  INV3 U238 ( .A(\u_decoder/fir_filter/dp_cluster_0/r179/CARRYB[6][1] ), .Q(
        n658) );
  INV3 U239 ( .A(\u_decoder/fir_filter/dp_cluster_0/r179/SUMB[5][3] ), .Q(n657) );
  INV3 U240 ( .A(\u_decoder/fir_filter/I_data_mult_3 [10]), .Q(n2281) );
  IMUX21 U241 ( .A(n2927), .B(n2928), .S(
        \u_decoder/fir_filter/dp_cluster_0/r167/A2[8] ), .Q(n2926) );
  NOR21 U242 ( .A(\u_decoder/fir_filter/dp_cluster_0/r167/A1[8] ), .B(n2282), 
        .Q(n2928) );
  INV3 U243 ( .A(\u_decoder/fir_filter/Q_data_mult_3 [10]), .Q(n2352) );
  IMUX21 U244 ( .A(n2841), .B(n2842), .S(
        \u_decoder/fir_filter/dp_cluster_0/r180/A2[8] ), .Q(n2840) );
  NOR21 U245 ( .A(\u_decoder/fir_filter/dp_cluster_0/r180/A1[8] ), .B(n2353), 
        .Q(n2842) );
  INV3 U246 ( .A(n2882), .Q(n2292) );
  INV3 U247 ( .A(n2796), .Q(n2363) );
  NOR21 U248 ( .A(n581), .B(n582), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[7][0] ) );
  INV3 U249 ( .A(\u_decoder/fir_filter/dp_cluster_0/r167/SUMB[6][1] ), .Q(n581) );
  INV3 U250 ( .A(\u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[6][0] ), .Q(
        n582) );
  NOR21 U251 ( .A(n642), .B(n643), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[7][0] ) );
  INV3 U252 ( .A(\u_decoder/fir_filter/dp_cluster_0/r180/SUMB[6][1] ), .Q(n642) );
  INV3 U253 ( .A(\u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[6][0] ), .Q(
        n643) );
  NOR21 U254 ( .A(n618), .B(n619), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r164/CARRYB[7][0] ) );
  INV3 U255 ( .A(\u_decoder/fir_filter/dp_cluster_0/r164/SUMB[5][2] ), .Q(n618) );
  INV3 U256 ( .A(\u_decoder/fir_filter/dp_cluster_0/r164/CARRYB[6][0] ), .Q(
        n619) );
  NOR21 U257 ( .A(n679), .B(n680), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r177/CARRYB[7][0] ) );
  INV3 U258 ( .A(\u_decoder/fir_filter/dp_cluster_0/r177/SUMB[5][2] ), .Q(n679) );
  INV3 U259 ( .A(\u_decoder/fir_filter/dp_cluster_0/r177/CARRYB[6][0] ), .Q(
        n680) );
  AOI211 U260 ( .A(n2251), .B(\u_decoder/fir_filter/dp_cluster_0/r166/A1[7] ), 
        .C(n2249), .Q(n2913) );
  INV3 U261 ( .A(n2919), .Q(n2249) );
  AOI211 U262 ( .A(n2322), .B(\u_decoder/fir_filter/dp_cluster_0/r179/A1[7] ), 
        .C(n2320), .Q(n2827) );
  INV3 U263 ( .A(n2833), .Q(n2320) );
  NAND22 U264 ( .A(\u_decoder/fir_filter/dp_cluster_0/r164/PROD1[4] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r164/A1[3] ), .Q(n2888) );
  NAND22 U265 ( .A(\u_decoder/fir_filter/dp_cluster_0/r177/PROD1[4] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r177/A1[3] ), .Q(n2802) );
  XOR21 U266 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_276/SUMB[4][3] ), 
        .B(\u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[6][0] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/SUMB[7][0] ) );
  XOR21 U267 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_308/SUMB[4][3] ), 
        .B(\u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[6][0] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/SUMB[7][0] ) );
  XNR31 U268 ( .A(\u_decoder/fir_filter/dp_cluster_0/r166/A2[8] ), .B(n2247), 
        .C(n2913), .Q(n329) );
  XNR31 U269 ( .A(\u_decoder/fir_filter/dp_cluster_0/r165/A2[9] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r165/A1[9] ), .C(n2897), .Q(n330)
         );
  XNR31 U270 ( .A(\u_decoder/fir_filter/dp_cluster_0/r165/A2[8] ), .B(n2240), 
        .C(n2898), .Q(n331) );
  XNR31 U271 ( .A(\u_decoder/fir_filter/dp_cluster_0/r165/A2[7] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r165/A1[7] ), .C(n2899), .Q(n332)
         );
  XNR31 U272 ( .A(\u_decoder/fir_filter/dp_cluster_0/r179/A2[8] ), .B(n2318), 
        .C(n2827), .Q(n333) );
  XNR31 U273 ( .A(\u_decoder/fir_filter/dp_cluster_0/r178/A2[9] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r178/A1[9] ), .C(n2811), .Q(n334)
         );
  XNR31 U274 ( .A(\u_decoder/fir_filter/dp_cluster_0/r178/A2[8] ), .B(n2311), 
        .C(n2812), .Q(n335) );
  XNR31 U275 ( .A(\u_decoder/fir_filter/dp_cluster_0/r178/A2[7] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r178/A1[7] ), .C(n2813), .Q(n336)
         );
  XOR21 U276 ( .A(n16), .B(
        \u_decoder/fir_filter/dp_cluster_0/r165/CARRYB[6][3] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r165/SUMB[7][3] ) );
  XOR21 U277 ( .A(n17), .B(
        \u_decoder/fir_filter/dp_cluster_0/r178/CARRYB[6][3] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r178/SUMB[7][3] ) );
  NOR31 U278 ( .A(n2295), .B(n2888), .C(n2294), .Q(n2884) );
  NOR31 U279 ( .A(n2366), .B(n2802), .C(n2365), .Q(n2798) );
  NAND22 U280 ( .A(\u_decoder/fir_filter/dp_cluster_0/r165/PROD1[5] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r165/A1[4] ), .Q(n2902) );
  NAND22 U281 ( .A(\u_decoder/fir_filter/dp_cluster_0/r178/PROD1[5] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r178/A1[4] ), .Q(n2816) );
  NOR21 U282 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_276/A2[10] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/A1[10] ), .Q(n2956) );
  NOR21 U283 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_308/A2[10] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/A1[10] ), .Q(n2870) );
  NOR21 U284 ( .A(\u_decoder/fir_filter/dp_cluster_0/r167/A2[9] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r167/A1[9] ), .Q(n2933) );
  NOR21 U285 ( .A(\u_decoder/fir_filter/dp_cluster_0/r180/A2[9] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r180/A1[9] ), .Q(n2847) );
  NOR21 U286 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_276/A1[8] ), .B(
        n2266), .Q(n2950) );
  INV3 U287 ( .A(n2946), .Q(n2266) );
  NOR21 U288 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_308/A1[8] ), .B(
        n2337), .Q(n2864) );
  INV3 U289 ( .A(n2860), .Q(n2337) );
  NAND22 U290 ( .A(\u_decoder/fir_filter/dp_cluster_0/r167/A2[8] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r167/A1[8] ), .Q(n2925) );
  NAND22 U291 ( .A(\u_decoder/fir_filter/dp_cluster_0/r180/A2[8] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r180/A1[8] ), .Q(n2839) );
  NAND22 U292 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_276/A2[10] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/A1[10] ), .Q(n2959) );
  NAND22 U293 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_308/A2[10] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/A1[10] ), .Q(n2873) );
  NOR21 U294 ( .A(n583), .B(n584), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[7][1] ) );
  INV3 U295 ( .A(\u_decoder/fir_filter/dp_cluster_0/r167/SUMB[5][3] ), .Q(n583) );
  INV3 U296 ( .A(\u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[6][1] ), .Q(
        n584) );
  NOR21 U297 ( .A(n644), .B(n645), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[7][1] ) );
  INV3 U298 ( .A(\u_decoder/fir_filter/dp_cluster_0/r180/SUMB[5][3] ), .Q(n644) );
  INV3 U299 ( .A(\u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[6][1] ), .Q(
        n645) );
  NOR21 U300 ( .A(n568), .B(n569), .Q(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[7][3] ) );
  INV3 U301 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[6][3] ), 
        .Q(n569) );
  INV3 U302 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_276/SUMB[5][5] ), .Q(
        n568) );
  NOR21 U303 ( .A(n629), .B(n630), .Q(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[7][3] ) );
  INV3 U304 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[6][3] ), 
        .Q(n630) );
  INV3 U305 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_308/SUMB[5][5] ), .Q(
        n629) );
  NOR21 U306 ( .A(n566), .B(n567), .Q(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[7][0] ) );
  INV3 U307 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_276/SUMB[4][3] ), .Q(
        n566) );
  INV3 U308 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[6][0] ), 
        .Q(n567) );
  NOR21 U309 ( .A(n10), .B(n608), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r165/CARRYB[7][3] ) );
  INV3 U310 ( .A(\u_decoder/fir_filter/dp_cluster_0/r165/CARRYB[6][3] ), .Q(
        n608) );
  NOR21 U311 ( .A(n10), .B(n620), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r164/CARRYB[7][2] ) );
  INV3 U312 ( .A(\u_decoder/fir_filter/dp_cluster_0/r164/CARRYB[6][2] ), .Q(
        n620) );
  NOR21 U313 ( .A(n9), .B(n669), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r178/CARRYB[7][3] ) );
  INV3 U314 ( .A(\u_decoder/fir_filter/dp_cluster_0/r178/CARRYB[6][3] ), .Q(
        n669) );
  NOR21 U315 ( .A(n9), .B(n681), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r177/CARRYB[7][2] ) );
  INV3 U316 ( .A(\u_decoder/fir_filter/dp_cluster_0/r177/CARRYB[6][2] ), .Q(
        n681) );
  XNR31 U317 ( .A(\u_decoder/fir_filter/dp_cluster_0/r166/A2[7] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r166/A1[7] ), .C(n2251), .Q(n337)
         );
  XNR31 U318 ( .A(\u_decoder/fir_filter/dp_cluster_0/r179/A2[7] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r179/A1[7] ), .C(n2322), .Q(n338)
         );
  XNR31 U319 ( .A(\u_decoder/fir_filter/dp_cluster_0/r164/A2[8] ), .B(n2297), 
        .C(n2880), .Q(n339) );
  XNR31 U320 ( .A(\u_decoder/fir_filter/dp_cluster_0/r177/A2[8] ), .B(n2368), 
        .C(n2794), .Q(n340) );
  INV3 U321 ( .A(\u_decoder/fir_filter/dp_cluster_0/r166/A1[8] ), .Q(n2247) );
  INV3 U322 ( .A(\u_decoder/fir_filter/dp_cluster_0/r179/A1[8] ), .Q(n2318) );
  INV3 U323 ( .A(\u_decoder/fir_filter/dp_cluster_0/r164/A1[8] ), .Q(n2297) );
  INV3 U324 ( .A(\u_decoder/fir_filter/dp_cluster_0/r177/A1[8] ), .Q(n2368) );
  INV3 U325 ( .A(\u_decoder/fir_filter/dp_cluster_0/r165/A1[8] ), .Q(n2240) );
  INV3 U326 ( .A(\u_decoder/fir_filter/dp_cluster_0/r178/A1[8] ), .Q(n2311) );
  NOR21 U327 ( .A(n627), .B(n628), .Q(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[7][0] ) );
  INV3 U328 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_308/SUMB[4][3] ), .Q(
        n627) );
  INV3 U329 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[6][0] ), 
        .Q(n628) );
  NOR21 U330 ( .A(\u_decoder/fir_filter/dp_cluster_0/r167/A2[10] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r167/A1[10] ), .Q(n2934) );
  NOR21 U331 ( .A(\u_decoder/fir_filter/dp_cluster_0/r180/A2[10] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r180/A1[10] ), .Q(n2848) );
  NAND22 U332 ( .A(\u_decoder/fir_filter/dp_cluster_0/r167/A2[9] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r167/A1[9] ), .Q(n2923) );
  NAND22 U333 ( .A(\u_decoder/fir_filter/dp_cluster_0/r180/A2[9] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r180/A1[9] ), .Q(n2837) );
  NAND22 U334 ( .A(\u_decoder/fir_filter/dp_cluster_0/r167/A2[10] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r167/A1[10] ), .Q(n2937) );
  NAND22 U335 ( .A(\u_decoder/fir_filter/dp_cluster_0/r180/A2[10] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r180/A1[10] ), .Q(n2851) );
  NOR21 U336 ( .A(n2888), .B(n2295), .Q(n2889) );
  NOR21 U337 ( .A(n2802), .B(n2366), .Q(n2803) );
  INV3 U338 ( .A(\u_decoder/fir_filter/dp_cluster_0/r164/A1[4] ), .Q(n2295) );
  INV3 U339 ( .A(\u_decoder/fir_filter/dp_cluster_0/r177/A1[4] ), .Q(n2366) );
  XNR31 U340 ( .A(\u_decoder/fir_filter/dp_cluster_0/r167/A1[7] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r167/A2[7] ), .C(n2929), .Q(n341)
         );
  XNR31 U341 ( .A(\u_decoder/fir_filter/dp_cluster_0/r180/A1[7] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r180/A2[7] ), .C(n2843), .Q(n342)
         );
  BUF2 U342 ( .A(\u_inFIFO/n224 ), .Q(n1203) );
  BUF2 U343 ( .A(\u_inFIFO/n224 ), .Q(n1204) );
  BUF2 U344 ( .A(\u_inFIFO/n224 ), .Q(n1205) );
  BUF2 U345 ( .A(\u_inFIFO/n224 ), .Q(n1206) );
  BUF2 U346 ( .A(\u_inFIFO/n224 ), .Q(n1207) );
  INV3 U347 ( .A(n1167), .Q(n1150) );
  INV3 U348 ( .A(n1191), .Q(n1184) );
  INV3 U349 ( .A(n1211), .Q(n1209) );
  INV3 U350 ( .A(\u_outFIFO/n1112 ), .Q(n1794) );
  XOR21 U351 ( .A(n2888), .B(\u_decoder/fir_filter/dp_cluster_0/r164/A1[4] ), 
        .Q(n343) );
  XOR21 U352 ( .A(n2802), .B(\u_decoder/fir_filter/dp_cluster_0/r177/A1[4] ), 
        .Q(n344) );
  INV3 U353 ( .A(\u_decoder/fir_filter/I_data_mult_3 [6]), .Q(n2284) );
  INV3 U354 ( .A(\u_decoder/fir_filter/I_data_mult_3 [5]), .Q(n2285) );
  INV3 U355 ( .A(\u_decoder/fir_filter/dp_cluster_0/r166/SUMB[5][1] ), .Q(
        n2252) );
  INV3 U356 ( .A(\u_decoder/fir_filter/Q_data_mult_3 [6]), .Q(n2355) );
  INV3 U357 ( .A(\u_decoder/fir_filter/Q_data_mult_3 [5]), .Q(n2356) );
  INV3 U358 ( .A(\u_decoder/fir_filter/dp_cluster_0/r179/SUMB[5][1] ), .Q(
        n2323) );
  BUF2 U359 ( .A(\u_inFIFO/n224 ), .Q(n1208) );
  INV3 U360 ( .A(n1145), .Q(n1144) );
  INV3 U361 ( .A(n1148), .Q(n1140) );
  INV3 U362 ( .A(n1146), .Q(n1139) );
  INV3 U363 ( .A(n1148), .Q(n1143) );
  INV3 U364 ( .A(n1146), .Q(n1142) );
  INV3 U365 ( .A(n1147), .Q(n1141) );
  INV3 U366 ( .A(n1149), .Q(n1138) );
  INV3 U367 ( .A(n1171), .Q(n1164) );
  INV3 U368 ( .A(n1171), .Q(n1165) );
  INV3 U369 ( .A(n1171), .Q(n1166) );
  INV3 U370 ( .A(n1170), .Q(n1162) );
  INV3 U371 ( .A(n1170), .Q(n1161) );
  INV3 U372 ( .A(n1171), .Q(n1163) );
  INV3 U373 ( .A(n1170), .Q(n1160) );
  INV3 U374 ( .A(n1168), .Q(n1156) );
  INV3 U375 ( .A(n1168), .Q(n1155) );
  INV3 U376 ( .A(n1168), .Q(n1154) );
  INV3 U377 ( .A(n1168), .Q(n1153) );
  INV3 U378 ( .A(n1167), .Q(n1152) );
  INV3 U379 ( .A(n1167), .Q(n1151) );
  INV3 U380 ( .A(n1169), .Q(n1159) );
  INV3 U381 ( .A(n1169), .Q(n1158) );
  INV3 U382 ( .A(n1169), .Q(n1157) );
  INV3 U383 ( .A(n1191), .Q(n1188) );
  INV3 U384 ( .A(n1191), .Q(n1185) );
  INV3 U385 ( .A(n1191), .Q(n1186) );
  INV3 U386 ( .A(n1191), .Q(n1187) );
  INV3 U387 ( .A(n1191), .Q(n1189) );
  INV3 U388 ( .A(n1191), .Q(n1190) );
  BUF2 U389 ( .A(n980), .Q(n1017) );
  BUF2 U390 ( .A(n979), .Q(n1016) );
  BUF2 U391 ( .A(n979), .Q(n1015) );
  BUF2 U392 ( .A(n978), .Q(n1014) );
  BUF2 U393 ( .A(n978), .Q(n1013) );
  BUF2 U394 ( .A(n977), .Q(n1012) );
  BUF2 U395 ( .A(n977), .Q(n1011) );
  BUF2 U396 ( .A(n976), .Q(n1010) );
  BUF2 U397 ( .A(n976), .Q(n1009) );
  BUF2 U398 ( .A(n975), .Q(n1008) );
  BUF2 U399 ( .A(n975), .Q(n1007) );
  BUF2 U400 ( .A(n974), .Q(n1006) );
  BUF2 U401 ( .A(n974), .Q(n1005) );
  BUF2 U402 ( .A(n973), .Q(n1004) );
  BUF2 U403 ( .A(n973), .Q(n1003) );
  BUF2 U404 ( .A(n972), .Q(n1002) );
  BUF2 U405 ( .A(n972), .Q(n1001) );
  BUF2 U406 ( .A(n971), .Q(n1000) );
  BUF2 U407 ( .A(n971), .Q(n999) );
  BUF2 U408 ( .A(n970), .Q(n998) );
  BUF2 U409 ( .A(n970), .Q(n997) );
  BUF2 U410 ( .A(n969), .Q(n996) );
  BUF2 U411 ( .A(n969), .Q(n995) );
  BUF2 U412 ( .A(n968), .Q(n994) );
  BUF2 U413 ( .A(n968), .Q(n993) );
  BUF2 U414 ( .A(n967), .Q(n992) );
  BUF2 U415 ( .A(n967), .Q(n991) );
  BUF2 U416 ( .A(n966), .Q(n990) );
  BUF2 U417 ( .A(n966), .Q(n989) );
  BUF2 U418 ( .A(n965), .Q(n988) );
  BUF2 U419 ( .A(n965), .Q(n987) );
  BUF2 U420 ( .A(n964), .Q(n986) );
  BUF2 U421 ( .A(n964), .Q(n985) );
  BUF2 U422 ( .A(n963), .Q(n984) );
  BUF2 U423 ( .A(n963), .Q(n983) );
  BUF2 U424 ( .A(n962), .Q(n982) );
  BUF2 U425 ( .A(n962), .Q(n981) );
  INV3 U426 ( .A(\u_decoder/fir_filter/I_data_mult_3 [4]), .Q(n2286) );
  INV3 U427 ( .A(\u_decoder/fir_filter/I_data_mult_3 [3]), .Q(n2287) );
  INV3 U428 ( .A(\u_decoder/fir_filter/dp_cluster_0/r166/SUMB[4][1] ), .Q(
        n2253) );
  INV3 U429 ( .A(\u_decoder/fir_filter/Q_data_mult_3 [4]), .Q(n2357) );
  INV3 U430 ( .A(\u_decoder/fir_filter/Q_data_mult_3 [3]), .Q(n2358) );
  INV3 U431 ( .A(\u_decoder/fir_filter/dp_cluster_0/r179/SUMB[4][1] ), .Q(
        n2324) );
  INV3 U432 ( .A(\u_decoder/fir_filter/I_data_mult_3 [2]), .Q(n2288) );
  INV3 U433 ( .A(\u_decoder/fir_filter/dp_cluster_0/r166/SUMB[3][1] ), .Q(
        n2254) );
  INV3 U434 ( .A(\u_decoder/fir_filter/I_data_mult_1[4] ), .Q(n2244) );
  INV3 U435 ( .A(\u_decoder/fir_filter/Q_data_mult_3 [2]), .Q(n2359) );
  INV3 U436 ( .A(\u_decoder/fir_filter/dp_cluster_0/r179/SUMB[3][1] ), .Q(
        n2325) );
  INV3 U437 ( .A(\u_decoder/fir_filter/Q_data_mult_1[4] ), .Q(n2315) );
  INV3 U438 ( .A(\u_decoder/fir_filter/I_data_mult_0 [3]), .Q(n2296) );
  INV3 U439 ( .A(\u_decoder/fir_filter/Q_data_mult_0 [3]), .Q(n2367) );
  BUF2 U440 ( .A(n980), .Q(n1018) );
  OAI2111 U441 ( .A(n1381), .B(n1363), .C(n1293), .D(n1337), .Q(
        \u_cdr/phd1/cnt_phd/N12 ) );
  NAND31 U442 ( .A(n1381), .B(n1380), .C(n1363), .Q(n1293) );
  AOI211 U443 ( .A(n1272), .B(n1275), .C(n1271), .Q(n1247) );
  OAI2111 U444 ( .A(n2663), .B(n2664), .C(n2665), .D(n2666), .Q(n3038) );
  NOR40 U445 ( .A(n2666), .B(n2665), .C(n2664), .D(n2663), .Q(
        \u_cordic/my_rotation/n57 ) );
  INV3 U446 ( .A(n767), .Q(n2674) );
  INV3 U447 ( .A(\u_cordic/my_rotation/n68 ), .Q(n2660) );
  AOI221 U448 ( .A(n768), .B(n2674), .C(\u_cordic/my_rotation/N40 ), .D(n767), 
        .Q(\u_cordic/my_rotation/n68 ) );
  XOR21 U449 ( .A(\u_cordic/my_rotation/add_38/carry [15]), .B(n767), .Q(
        \u_cordic/my_rotation/N40 ) );
  NOR21 U450 ( .A(n492), .B(n493), .Q(\u_cordic/my_rotation/add_38/carry [15])
         );
  AOI211 U451 ( .A(n3041), .B(n3040), .C(n2660), .Q(n3042) );
  NOR40 U452 ( .A(n2661), .B(n2662), .C(n2668), .D(n2667), .Q(n3040) );
  NOR40 U453 ( .A(n2673), .B(n2672), .C(n2671), .D(n3039), .Q(n3041) );
  AOI211 U454 ( .A(\u_cordic/my_rotation/n48 ), .B(n3038), .C(
        \u_cordic/my_rotation/n47 ), .Q(n3039) );
  INV3 U455 ( .A(\u_cordic/my_rotation/add_38/carry [14]), .Q(n492) );
  XOR21 U456 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_276/SUMB[7][3] ), 
        .B(\u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[7][2] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/A1[8] ) );
  XOR21 U457 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_308/SUMB[7][3] ), 
        .B(\u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[7][2] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/A1[8] ) );
  XOR21 U458 ( .A(\u_decoder/fir_filter/dp_cluster_0/r164/SUMB[7][1] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r164/CARRYB[7][0] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r164/A1[6] ) );
  XOR21 U459 ( .A(\u_decoder/fir_filter/dp_cluster_0/r177/SUMB[7][1] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r177/CARRYB[7][0] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r177/A1[6] ) );
  XOR21 U460 ( .A(\u_decoder/fir_filter/dp_cluster_0/r166/SUMB[7][1] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r166/CARRYB[7][0] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r166/A1[6] ) );
  XOR21 U461 ( .A(\u_decoder/fir_filter/dp_cluster_0/r179/SUMB[7][1] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r179/CARRYB[7][0] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r179/A1[6] ) );
  XOR21 U462 ( .A(\u_decoder/fir_filter/dp_cluster_0/r165/SUMB[7][1] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r165/CARRYB[7][0] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r165/A1[6] ) );
  XOR21 U463 ( .A(\u_decoder/fir_filter/dp_cluster_0/r178/SUMB[7][1] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r178/CARRYB[7][0] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r178/A1[6] ) );
  AOI311 U464 ( .A(n2894), .B(\u_decoder/fir_filter/dp_cluster_0/r164/A1[4] ), 
        .C(\u_decoder/fir_filter/dp_cluster_0/r164/A1[5] ), .D(n2895), .Q(
        n2880) );
  NOR21 U465 ( .A(n2896), .B(n2888), .Q(n2894) );
  MAJ31 U466 ( .A(\u_decoder/fir_filter/dp_cluster_0/r164/A2[7] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r164/A1[7] ), .C(n2292), .Q(n2895)
         );
  AOI311 U467 ( .A(n2808), .B(\u_decoder/fir_filter/dp_cluster_0/r177/A1[4] ), 
        .C(\u_decoder/fir_filter/dp_cluster_0/r177/A1[5] ), .D(n2809), .Q(
        n2794) );
  NOR21 U468 ( .A(n2810), .B(n2802), .Q(n2808) );
  MAJ31 U469 ( .A(\u_decoder/fir_filter/dp_cluster_0/r177/A2[7] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r177/A1[7] ), .C(n2363), .Q(n2809)
         );
  NOR40 U470 ( .A(n2933), .B(n2924), .C(n2934), .D(n2935), .Q(n2932) );
  NOR40 U471 ( .A(n2847), .B(n2838), .C(n2848), .D(n2849), .Q(n2846) );
  OAI311 U472 ( .A(n2243), .B(n2903), .C(n2902), .D(n2911), .Q(n2899) );
  NAND22 U473 ( .A(\u_decoder/fir_filter/dp_cluster_0/r165/A2[6] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r165/A1[6] ), .Q(n2911) );
  OAI311 U474 ( .A(n2314), .B(n2817), .C(n2816), .D(n2825), .Q(n2813) );
  NAND22 U475 ( .A(\u_decoder/fir_filter/dp_cluster_0/r178/A2[6] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r178/A1[6] ), .Q(n2825) );
  XOR21 U476 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_276/SUMB[7][4] ), 
        .B(\u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[7][3] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/A1[9] ) );
  XOR21 U477 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_308/SUMB[7][4] ), 
        .B(\u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[7][3] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/A1[9] ) );
  XOR21 U478 ( .A(\u_decoder/fir_filter/dp_cluster_0/r164/SUMB[7][2] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r164/CARRYB[7][1] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r164/A1[7] ) );
  XOR21 U479 ( .A(\u_decoder/fir_filter/dp_cluster_0/r177/SUMB[7][2] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r177/CARRYB[7][1] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r177/A1[7] ) );
  XOR21 U480 ( .A(\u_decoder/fir_filter/dp_cluster_0/r166/SUMB[7][2] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r166/CARRYB[7][1] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r166/A1[7] ) );
  XOR21 U481 ( .A(\u_decoder/fir_filter/dp_cluster_0/r165/SUMB[7][2] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r165/CARRYB[7][1] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r165/A1[7] ) );
  XOR21 U482 ( .A(\u_decoder/fir_filter/dp_cluster_0/r179/SUMB[7][2] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r179/CARRYB[7][1] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r179/A1[7] ) );
  XOR21 U483 ( .A(\u_decoder/fir_filter/dp_cluster_0/r178/SUMB[7][2] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r178/CARRYB[7][1] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r178/A1[7] ) );
  XNR31 U484 ( .A(\u_decoder/fir_filter/dp_cluster_0/r167/A2[11] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[7][5] ), .C(n2939), .Q(
        n345) );
  XNR31 U485 ( .A(\u_decoder/fir_filter/dp_cluster_0/r180/A2[11] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[7][5] ), .C(n2853), .Q(
        n346) );
  XOR21 U486 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_276/SUMB[7][2] ), 
        .B(\u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[7][1] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/A1[7] ) );
  XOR21 U487 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_308/SUMB[7][2] ), 
        .B(\u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[7][1] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/A1[7] ) );
  XOR21 U488 ( .A(n8), .B(\u_decoder/fir_filter/I_data_mult_0 [0]), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r167/SUMB[3][3] ) );
  XOR21 U489 ( .A(n7), .B(\u_decoder/fir_filter/Q_data_mult_0 [0]), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r180/SUMB[3][3] ) );
  XOR21 U490 ( .A(n4), .B(n84), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r165/SUMB[2][3] ) );
  XOR21 U491 ( .A(n3), .B(n88), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r178/SUMB[2][3] ) );
  XOR21 U492 ( .A(n4), .B(\u_decoder/fir_filter/I_data_mult_0 [0]), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r167/SUMB[2][1] ) );
  XOR21 U493 ( .A(n3), .B(\u_decoder/fir_filter/Q_data_mult_0 [0]), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r180/SUMB[2][1] ) );
  XOR21 U494 ( .A(n4), .B(n84), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r164/SUMB[2][2] ) );
  XOR21 U495 ( .A(n3), .B(n88), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r177/SUMB[2][2] ) );
  NOR21 U496 ( .A(n89), .B(\u_decoder/fir_filter/I_data_mult_0 [0]), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r165/CARRYB[2][3] ) );
  NOR21 U497 ( .A(n90), .B(\u_decoder/fir_filter/Q_data_mult_0 [0]), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r178/CARRYB[2][3] ) );
  NOR21 U498 ( .A(n89), .B(\u_decoder/fir_filter/I_data_mult_0 [0]), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r164/CARRYB[2][2] ) );
  NOR21 U499 ( .A(n90), .B(\u_decoder/fir_filter/Q_data_mult_0 [0]), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r177/CARRYB[2][2] ) );
  NOR21 U500 ( .A(n89), .B(n84), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r166/CARRYB[2][1] ) );
  XOR21 U501 ( .A(\u_decoder/fir_filter/I_data_mult_0 [0]), .B(n12), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r166/SUMB[1][3] ) );
  NOR21 U502 ( .A(n90), .B(n88), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r179/CARRYB[2][1] ) );
  XOR21 U503 ( .A(\u_decoder/fir_filter/Q_data_mult_0 [0]), .B(n11), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r179/SUMB[1][3] ) );
  NOR21 U504 ( .A(n89), .B(n84), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[2][1] ) );
  NOR21 U505 ( .A(n90), .B(n88), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[2][1] ) );
  NOR21 U506 ( .A(n89), .B(n84), .Q(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[2][3] ) );
  XOR21 U507 ( .A(\u_decoder/fir_filter/I_data_mult_0 [0]), .B(n12), .Q(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/SUMB[1][5] ) );
  NOR21 U508 ( .A(n90), .B(n88), .Q(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[2][3] ) );
  XOR21 U509 ( .A(\u_decoder/fir_filter/Q_data_mult_0 [0]), .B(n11), .Q(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/SUMB[1][5] ) );
  NOR21 U510 ( .A(n84), .B(n80), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r165/CARRYB[3][0] ) );
  NOR21 U511 ( .A(n88), .B(n81), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r178/CARRYB[3][0] ) );
  NOR21 U512 ( .A(n84), .B(n89), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r164/CARRYB[2][0] ) );
  NOR21 U513 ( .A(n88), .B(n90), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r177/CARRYB[2][0] ) );
  NOR21 U514 ( .A(n84), .B(n74), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r166/CARRYB[1][3] ) );
  NOR21 U515 ( .A(n88), .B(n75), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r179/CARRYB[1][3] ) );
  NOR21 U516 ( .A(n74), .B(n84), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[1][0] ) );
  NOR21 U517 ( .A(n75), .B(n88), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[1][0] ) );
  NOR21 U518 ( .A(n84), .B(n74), .Q(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[1][5] ) );
  NOR21 U519 ( .A(n88), .B(n75), .Q(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[1][5] ) );
  NAND22 U520 ( .A(\u_decoder/fir_filter/dp_cluster_0/r164/A2[6] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r164/A1[6] ), .Q(n2882) );
  NAND22 U521 ( .A(\u_decoder/fir_filter/dp_cluster_0/r177/A2[6] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r177/A1[6] ), .Q(n2796) );
  NOR21 U522 ( .A(n363), .B(n321), .Q(n2929) );
  NOR21 U523 ( .A(n364), .B(n322), .Q(n2843) );
  NOR21 U524 ( .A(n365), .B(n347), .Q(n2951) );
  NOR21 U525 ( .A(n366), .B(n348), .Q(n2865) );
  NOR21 U526 ( .A(\u_decoder/fir_filter/dp_cluster_0/r165/A2[6] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r165/A1[6] ), .Q(n2903) );
  NOR21 U527 ( .A(\u_decoder/fir_filter/dp_cluster_0/r178/A2[6] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r178/A1[6] ), .Q(n2817) );
  INV3 U528 ( .A(n2920), .Q(n2251) );
  NAND22 U529 ( .A(\u_decoder/fir_filter/dp_cluster_0/r166/A2[6] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r166/A1[6] ), .Q(n2920) );
  INV3 U530 ( .A(n2834), .Q(n2322) );
  NAND22 U531 ( .A(\u_decoder/fir_filter/dp_cluster_0/r179/A2[6] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r179/A1[6] ), .Q(n2834) );
  INV3 U532 ( .A(\u_decoder/fir_filter/dp_cluster_0/r165/A1[5] ), .Q(n2243) );
  INV3 U533 ( .A(\u_decoder/fir_filter/dp_cluster_0/r178/A1[5] ), .Q(n2314) );
  XNR21 U534 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_276/SUMB[7][1] ), 
        .B(\u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[7][0] ), .Q(n347) );
  XNR21 U535 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_308/SUMB[7][1] ), 
        .B(\u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[7][0] ), .Q(n348) );
  NOR21 U536 ( .A(n610), .B(n611), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r165/A2[7] ) );
  INV3 U537 ( .A(\u_decoder/fir_filter/dp_cluster_0/r165/CARRYB[7][0] ), .Q(
        n610) );
  INV3 U538 ( .A(\u_decoder/fir_filter/dp_cluster_0/r165/SUMB[7][1] ), .Q(n611) );
  NOR21 U539 ( .A(n671), .B(n672), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r178/A2[7] ) );
  INV3 U540 ( .A(\u_decoder/fir_filter/dp_cluster_0/r178/CARRYB[7][0] ), .Q(
        n671) );
  INV3 U541 ( .A(\u_decoder/fir_filter/dp_cluster_0/r178/SUMB[7][1] ), .Q(n672) );
  NOR21 U542 ( .A(n622), .B(n623), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r164/A2[7] ) );
  INV3 U543 ( .A(\u_decoder/fir_filter/dp_cluster_0/r164/CARRYB[7][0] ), .Q(
        n622) );
  INV3 U544 ( .A(\u_decoder/fir_filter/dp_cluster_0/r164/SUMB[7][1] ), .Q(n623) );
  NOR21 U545 ( .A(n683), .B(n684), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r177/A2[7] ) );
  INV3 U546 ( .A(\u_decoder/fir_filter/dp_cluster_0/r177/CARRYB[7][0] ), .Q(
        n683) );
  INV3 U547 ( .A(\u_decoder/fir_filter/dp_cluster_0/r177/SUMB[7][1] ), .Q(n684) );
  NAND22 U548 ( .A(\u_decoder/fir_filter/I_data_mult_0_15 ), .B(n1083), .Q(
        \u_decoder/fir_filter/n1019 ) );
  XOR21 U549 ( .A(n2891), .B(
        \u_decoder/fir_filter/dp_cluster_0/r164/CARRYB[7][3] ), .Q(
        \u_decoder/fir_filter/I_data_mult_0_15 ) );
  AOI211 U550 ( .A(n2879), .B(n2305), .C(n2289), .Q(n2891) );
  INV3 U551 ( .A(n2892), .Q(n2289) );
  NAND22 U552 ( .A(\u_decoder/fir_filter/Q_data_mult_0_15 ), .B(n1083), .Q(
        \u_decoder/fir_filter/n722 ) );
  XOR21 U553 ( .A(n2805), .B(
        \u_decoder/fir_filter/dp_cluster_0/r177/CARRYB[7][3] ), .Q(
        \u_decoder/fir_filter/Q_data_mult_0_15 ) );
  AOI211 U554 ( .A(n2793), .B(n2376), .C(n2360), .Q(n2805) );
  INV3 U555 ( .A(n2806), .Q(n2360) );
  NAND22 U556 ( .A(\u_decoder/fir_filter/I_data_mult_1_15 ), .B(n1083), .Q(
        \u_decoder/fir_filter/n1033 ) );
  XOR21 U557 ( .A(n2905), .B(
        \u_decoder/fir_filter/dp_cluster_0/r165/CARRYB[7][4] ), .Q(
        \u_decoder/fir_filter/I_data_mult_1_15 ) );
  AOI211 U558 ( .A(n2906), .B(n2305), .C(n2237), .Q(n2905) );
  INV3 U559 ( .A(n2907), .Q(n2237) );
  NAND22 U560 ( .A(\u_decoder/fir_filter/Q_data_mult_1_15 ), .B(n1083), .Q(
        \u_decoder/fir_filter/n736 ) );
  XOR21 U561 ( .A(n2819), .B(
        \u_decoder/fir_filter/dp_cluster_0/r178/CARRYB[7][4] ), .Q(
        \u_decoder/fir_filter/Q_data_mult_1_15 ) );
  AOI211 U562 ( .A(n2820), .B(n2376), .C(n2308), .Q(n2819) );
  INV3 U563 ( .A(n2821), .Q(n2308) );
  XOR21 U564 ( .A(\u_decoder/fir_filter/dp_cluster_0/r167/SUMB[7][3] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[7][2] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r167/A1[8] ) );
  XOR21 U565 ( .A(\u_decoder/fir_filter/dp_cluster_0/r180/SUMB[7][3] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[7][2] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r180/A1[8] ) );
  INV3 U566 ( .A(\u_decoder/iq_demod/dp_cluster_1/mult_150/CARRYB[3][3] ), .Q(
        n2389) );
  NOR21 U567 ( .A(n716), .B(n717), .Q(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/A2[5] ) );
  AOI211 U568 ( .A(n2773), .B(\u_decoder/iq_demod/dp_cluster_1/mult_150/A1[4] ), .C(n2380), .Q(n2772) );
  XOR21 U569 ( .A(\u_decoder/fir_filter/dp_cluster_0/r165/SUMB[7][4] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r165/CARRYB[7][3] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r165/A1[9] ) );
  XOR21 U570 ( .A(\u_decoder/fir_filter/dp_cluster_0/r178/SUMB[7][4] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r178/CARRYB[7][3] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r178/A1[9] ) );
  XOR21 U571 ( .A(\u_decoder/fir_filter/dp_cluster_0/r167/SUMB[7][4] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[7][3] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r167/A1[9] ) );
  XOR21 U572 ( .A(\u_decoder/fir_filter/dp_cluster_0/r180/SUMB[7][4] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[7][3] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r180/A1[9] ) );
  XOR21 U573 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_276/SUMB[7][5] ), 
        .B(\u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[7][4] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/A1[10] ) );
  XOR21 U574 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_308/SUMB[7][5] ), 
        .B(\u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[7][4] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/A1[10] ) );
  XOR21 U575 ( .A(n6), .B(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[6][5] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/SUMB[7][5] ) );
  XOR21 U576 ( .A(n6), .B(
        \u_decoder/fir_filter/dp_cluster_0/r166/CARRYB[6][3] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r166/SUMB[7][3] ) );
  XOR21 U577 ( .A(n5), .B(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[6][5] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/SUMB[7][5] ) );
  XOR21 U578 ( .A(n5), .B(
        \u_decoder/fir_filter/dp_cluster_0/r179/CARRYB[6][3] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r179/SUMB[7][3] ) );
  XOR21 U579 ( .A(\u_decoder/I_prefilter [4]), .B(
        \u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[6][3] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r167/SUMB[7][3] ) );
  XOR21 U580 ( .A(\u_decoder/Q_prefilter [4]), .B(
        \u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[6][3] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r180/SUMB[7][3] ) );
  XOR21 U581 ( .A(\u_decoder/fir_filter/dp_cluster_0/r166/SUMB[7][3] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r166/CARRYB[7][2] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r166/A1[8] ) );
  XOR21 U582 ( .A(\u_decoder/fir_filter/dp_cluster_0/r165/SUMB[7][3] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r165/CARRYB[7][2] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r165/A1[8] ) );
  XOR21 U583 ( .A(\u_decoder/fir_filter/dp_cluster_0/r179/SUMB[7][3] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r179/CARRYB[7][2] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r179/A1[8] ) );
  XOR21 U584 ( .A(\u_decoder/fir_filter/dp_cluster_0/r178/SUMB[7][3] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r178/CARRYB[7][2] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r178/A1[8] ) );
  XOR21 U585 ( .A(\u_decoder/fir_filter/dp_cluster_0/r164/SUMB[7][3] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r164/CARRYB[7][2] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r164/A1[8] ) );
  XOR21 U586 ( .A(\u_decoder/fir_filter/dp_cluster_0/r177/SUMB[7][3] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r177/CARRYB[7][2] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r177/A1[8] ) );
  NOR21 U587 ( .A(n588), .B(n589), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r167/A2[8] ) );
  INV3 U588 ( .A(\u_decoder/fir_filter/dp_cluster_0/r167/SUMB[7][2] ), .Q(n589) );
  INV3 U589 ( .A(\u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[7][1] ), .Q(
        n588) );
  NOR21 U590 ( .A(n649), .B(n650), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r180/A2[8] ) );
  INV3 U591 ( .A(\u_decoder/fir_filter/dp_cluster_0/r180/SUMB[7][2] ), .Q(n650) );
  INV3 U592 ( .A(\u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[7][1] ), .Q(
        n649) );
  NOR21 U593 ( .A(n573), .B(n574), .Q(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/A2[8] ) );
  INV3 U594 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[7][1] ), 
        .Q(n573) );
  INV3 U595 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_276/SUMB[7][2] ), .Q(
        n574) );
  NOR21 U596 ( .A(n634), .B(n635), .Q(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/A2[8] ) );
  INV3 U597 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[7][1] ), 
        .Q(n634) );
  INV3 U598 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_308/SUMB[7][2] ), .Q(
        n635) );
  NAND22 U599 ( .A(n2882), .B(n2883), .Q(n2881) );
  NAND22 U600 ( .A(n2796), .B(n2797), .Q(n2795) );
  AOI211 U601 ( .A(\u_decoder/iq_demod/dp_cluster_0/mult_151/A2[3] ), .B(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/A1[3] ), .C(n2789), .Q(n2792) );
  AOI211 U602 ( .A(\u_decoder/iq_demod/dp_cluster_1/mult_150/A2[3] ), .B(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/A1[3] ), .C(n2775), .Q(n2778) );
  AOI211 U603 ( .A(\u_decoder/iq_demod/dp_cluster_1/mult_149/A2[3] ), .B(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/A1[3] ), .C(n2768), .Q(n2771) );
  AOI211 U604 ( .A(\u_decoder/iq_demod/dp_cluster_0/mult_148/A2[3] ), .B(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/A1[3] ), .C(n2782), .Q(n2785) );
  AOI211 U605 ( .A(n2787), .B(\u_decoder/iq_demod/dp_cluster_0/mult_151/A1[4] ), .C(n2384), .Q(n2786) );
  INV3 U606 ( .A(n2788), .Q(n2384) );
  AOI211 U607 ( .A(n2766), .B(\u_decoder/iq_demod/dp_cluster_1/mult_149/A1[4] ), .C(n2390), .Q(n2765) );
  INV3 U608 ( .A(n2767), .Q(n2390) );
  XOR21 U609 ( .A(\u_decoder/fir_filter/dp_cluster_0/r167/SUMB[7][2] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[7][1] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r167/A1[7] ) );
  XOR21 U610 ( .A(\u_decoder/fir_filter/dp_cluster_0/r180/SUMB[7][2] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[7][1] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r180/A1[7] ) );
  XOR21 U611 ( .A(n4), .B(\u_decoder/fir_filter/I_data_mult_0 [0]), .Q(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/SUMB[2][3] ) );
  XOR21 U612 ( .A(n3), .B(\u_decoder/fir_filter/Q_data_mult_0 [0]), .Q(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/SUMB[2][3] ) );
  NOR21 U613 ( .A(n80), .B(n84), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[3][3] ) );
  NOR21 U614 ( .A(n81), .B(n88), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[3][3] ) );
  NOR21 U615 ( .A(n84), .B(n80), .Q(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[3][0] ) );
  NOR21 U616 ( .A(n88), .B(n81), .Q(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[3][0] ) );
  XNR21 U617 ( .A(\u_decoder/iq_demod/dp_cluster_1/mult_149/A1[2] ), .B(n2392), 
        .Q(\u_decoder/iq_demod/dp_cluster_1/mult_I_sin_out [4]) );
  XNR21 U618 ( .A(\u_decoder/iq_demod/dp_cluster_1/mult_150/A1[2] ), .B(n2382), 
        .Q(\u_decoder/iq_demod/dp_cluster_1/mult_Q_cos_out [4]) );
  NOR21 U619 ( .A(\u_decoder/fir_filter/dp_cluster_0/r164/A1[6] ), .B(n2293), 
        .Q(n2887) );
  INV3 U620 ( .A(\u_decoder/fir_filter/dp_cluster_0/r164/A2[6] ), .Q(n2293) );
  NOR21 U621 ( .A(\u_decoder/fir_filter/dp_cluster_0/r177/A1[6] ), .B(n2364), 
        .Q(n2801) );
  INV3 U622 ( .A(\u_decoder/fir_filter/dp_cluster_0/r177/A2[6] ), .Q(n2364) );
  XNR31 U623 ( .A(\u_decoder/iq_demod/dp_cluster_0/mult_151/A2[4] ), .B(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/A1[4] ), .C(n2787), .Q(n349)
         );
  XNR21 U624 ( .A(n2784), .B(n2785), .Q(
        \u_decoder/iq_demod/dp_cluster_0/mult_I_cos_out [5]) );
  XNR21 U625 ( .A(\u_decoder/iq_demod/dp_cluster_0/mult_148/A1[2] ), .B(n2395), 
        .Q(\u_decoder/iq_demod/dp_cluster_0/mult_I_cos_out [4]) );
  NOR21 U626 ( .A(\u_decoder/iq_demod/dp_cluster_0/mult_151/A2[3] ), .B(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/A1[3] ), .Q(n2789) );
  NOR21 U627 ( .A(\u_decoder/iq_demod/dp_cluster_1/mult_150/A2[3] ), .B(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/A1[3] ), .Q(n2775) );
  NOR21 U628 ( .A(\u_decoder/iq_demod/dp_cluster_1/mult_149/A2[3] ), .B(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/A1[3] ), .Q(n2768) );
  NOR21 U629 ( .A(\u_decoder/iq_demod/dp_cluster_0/mult_148/A2[3] ), .B(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/A1[3] ), .Q(n2782) );
  NOR21 U630 ( .A(n577), .B(n578), .Q(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/A2[10] ) );
  INV3 U631 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[7][3] ), 
        .Q(n577) );
  INV3 U632 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_276/SUMB[7][4] ), .Q(
        n578) );
  NOR21 U633 ( .A(n638), .B(n639), .Q(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/A2[10] ) );
  INV3 U634 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[7][3] ), 
        .Q(n638) );
  INV3 U635 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_308/SUMB[7][4] ), .Q(
        n639) );
  NOR21 U636 ( .A(n590), .B(n591), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r167/A2[9] ) );
  INV3 U637 ( .A(\u_decoder/fir_filter/dp_cluster_0/r167/SUMB[7][3] ), .Q(n591) );
  INV3 U638 ( .A(\u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[7][2] ), .Q(
        n590) );
  NOR21 U639 ( .A(n651), .B(n652), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r180/A2[9] ) );
  INV3 U640 ( .A(\u_decoder/fir_filter/dp_cluster_0/r180/SUMB[7][3] ), .Q(n652) );
  INV3 U641 ( .A(\u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[7][2] ), .Q(
        n651) );
  INV3 U642 ( .A(\u_decoder/fir_filter/I_data_mult_0 [8]), .Q(n2291) );
  IMUX21 U643 ( .A(n2887), .B(n2292), .S(n2884), .Q(n2886) );
  XNR21 U644 ( .A(\u_decoder/fir_filter/dp_cluster_0/r164/A1[6] ), .B(n2884), 
        .Q(n2885) );
  INV3 U645 ( .A(\u_decoder/fir_filter/Q_data_mult_0 [8]), .Q(n2362) );
  IMUX21 U646 ( .A(n2801), .B(n2363), .S(n2798), .Q(n2800) );
  XNR21 U647 ( .A(\u_decoder/fir_filter/dp_cluster_0/r177/A1[6] ), .B(n2798), 
        .Q(n2799) );
  NOR21 U648 ( .A(n579), .B(n580), .Q(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/A2[11] ) );
  INV3 U649 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[7][4] ), 
        .Q(n579) );
  INV3 U650 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_276/SUMB[7][5] ), .Q(
        n580) );
  NOR21 U651 ( .A(n640), .B(n641), .Q(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/A2[11] ) );
  INV3 U652 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[7][4] ), 
        .Q(n640) );
  INV3 U653 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_308/SUMB[7][5] ), .Q(
        n641) );
  NOR21 U654 ( .A(n571), .B(n572), .Q(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/A2[7] ) );
  INV3 U655 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[7][0] ), 
        .Q(n571) );
  INV3 U656 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_276/SUMB[7][1] ), .Q(
        n572) );
  NOR21 U657 ( .A(n632), .B(n633), .Q(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/A2[7] ) );
  INV3 U658 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[7][0] ), 
        .Q(n632) );
  INV3 U659 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_308/SUMB[7][1] ), .Q(
        n633) );
  INV3 U660 ( .A(\u_decoder/fir_filter/dp_cluster_0/r164/A1[5] ), .Q(n2294) );
  INV3 U661 ( .A(\u_decoder/fir_filter/dp_cluster_0/r177/A1[5] ), .Q(n2365) );
  NOR21 U662 ( .A(n600), .B(n601), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r166/A2[7] ) );
  INV3 U663 ( .A(\u_decoder/fir_filter/dp_cluster_0/r166/CARRYB[7][0] ), .Q(
        n600) );
  INV3 U664 ( .A(\u_decoder/fir_filter/dp_cluster_0/r166/SUMB[7][1] ), .Q(n601) );
  NOR21 U665 ( .A(n661), .B(n662), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r179/A2[7] ) );
  INV3 U666 ( .A(\u_decoder/fir_filter/dp_cluster_0/r179/CARRYB[7][0] ), .Q(
        n661) );
  INV3 U667 ( .A(\u_decoder/fir_filter/dp_cluster_0/r179/SUMB[7][1] ), .Q(n662) );
  NOR21 U668 ( .A(n604), .B(n605), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r166/A2[9] ) );
  INV3 U669 ( .A(\u_decoder/fir_filter/dp_cluster_0/r166/SUMB[7][3] ), .Q(n605) );
  INV3 U670 ( .A(\u_decoder/fir_filter/dp_cluster_0/r166/CARRYB[7][2] ), .Q(
        n604) );
  NOR21 U671 ( .A(n665), .B(n666), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r179/A2[9] ) );
  INV3 U672 ( .A(\u_decoder/fir_filter/dp_cluster_0/r179/SUMB[7][3] ), .Q(n666) );
  INV3 U673 ( .A(\u_decoder/fir_filter/dp_cluster_0/r179/CARRYB[7][2] ), .Q(
        n665) );
  OAI311 U674 ( .A(n2386), .B(n2789), .C(n2385), .D(n2790), .Q(n2787) );
  NAND22 U675 ( .A(\u_decoder/iq_demod/dp_cluster_0/mult_151/A2[3] ), .B(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/A1[3] ), .Q(n2790) );
  INV3 U676 ( .A(\u_decoder/iq_demod/dp_cluster_0/mult_151/A1[2] ), .Q(n2385)
         );
  OAI311 U677 ( .A(n2382), .B(n2775), .C(n2381), .D(n2776), .Q(n2773) );
  NAND22 U678 ( .A(\u_decoder/iq_demod/dp_cluster_1/mult_150/A2[3] ), .B(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/A1[3] ), .Q(n2776) );
  INV3 U679 ( .A(\u_decoder/iq_demod/dp_cluster_1/mult_150/A1[2] ), .Q(n2381)
         );
  OAI311 U680 ( .A(n2392), .B(n2768), .C(n2391), .D(n2769), .Q(n2766) );
  NAND22 U681 ( .A(\u_decoder/iq_demod/dp_cluster_1/mult_149/A2[3] ), .B(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/A1[3] ), .Q(n2769) );
  INV3 U682 ( .A(\u_decoder/iq_demod/dp_cluster_1/mult_149/A1[2] ), .Q(n2391)
         );
  OAI311 U683 ( .A(n2395), .B(n2782), .C(n2394), .D(n2783), .Q(n2780) );
  NAND22 U684 ( .A(\u_decoder/iq_demod/dp_cluster_0/mult_148/A2[3] ), .B(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/A1[3] ), .Q(n2783) );
  INV3 U685 ( .A(\u_decoder/iq_demod/dp_cluster_0/mult_148/A1[2] ), .Q(n2394)
         );
  XNR31 U686 ( .A(\u_decoder/iq_demod/dp_cluster_0/mult_151/A2[5] ), .B(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/CARRYB[3][3] ), .C(n2786), 
        .Q(n350) );
  NOR21 U687 ( .A(n602), .B(n603), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r166/A2[8] ) );
  INV3 U688 ( .A(\u_decoder/fir_filter/dp_cluster_0/r166/CARRYB[7][1] ), .Q(
        n602) );
  INV3 U689 ( .A(\u_decoder/fir_filter/dp_cluster_0/r166/SUMB[7][2] ), .Q(n603) );
  NOR21 U690 ( .A(n663), .B(n664), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r179/A2[8] ) );
  INV3 U691 ( .A(\u_decoder/fir_filter/dp_cluster_0/r179/CARRYB[7][1] ), .Q(
        n663) );
  INV3 U692 ( .A(\u_decoder/fir_filter/dp_cluster_0/r179/SUMB[7][2] ), .Q(n664) );
  NOR21 U693 ( .A(n612), .B(n613), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r165/A2[8] ) );
  INV3 U694 ( .A(\u_decoder/fir_filter/dp_cluster_0/r165/CARRYB[7][1] ), .Q(
        n612) );
  INV3 U695 ( .A(\u_decoder/fir_filter/dp_cluster_0/r165/SUMB[7][2] ), .Q(n613) );
  NOR21 U696 ( .A(n673), .B(n674), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r178/A2[8] ) );
  INV3 U697 ( .A(\u_decoder/fir_filter/dp_cluster_0/r178/CARRYB[7][1] ), .Q(
        n673) );
  INV3 U698 ( .A(\u_decoder/fir_filter/dp_cluster_0/r178/SUMB[7][2] ), .Q(n674) );
  NOR21 U699 ( .A(n575), .B(n576), .Q(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/A2[9] ) );
  INV3 U700 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[7][2] ), 
        .Q(n575) );
  INV3 U701 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_276/SUMB[7][3] ), .Q(
        n576) );
  NOR21 U702 ( .A(n636), .B(n637), .Q(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/A2[9] ) );
  INV3 U703 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[7][2] ), 
        .Q(n636) );
  INV3 U704 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_308/SUMB[7][3] ), .Q(
        n637) );
  NOR21 U705 ( .A(n614), .B(n615), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r165/A2[9] ) );
  INV3 U706 ( .A(\u_decoder/fir_filter/dp_cluster_0/r165/CARRYB[7][2] ), .Q(
        n614) );
  INV3 U707 ( .A(\u_decoder/fir_filter/dp_cluster_0/r165/SUMB[7][3] ), .Q(n615) );
  NOR21 U708 ( .A(n624), .B(n625), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r164/A2[8] ) );
  INV3 U709 ( .A(\u_decoder/fir_filter/dp_cluster_0/r164/CARRYB[7][1] ), .Q(
        n624) );
  INV3 U710 ( .A(\u_decoder/fir_filter/dp_cluster_0/r164/SUMB[7][2] ), .Q(n625) );
  NOR21 U711 ( .A(n675), .B(n676), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r178/A2[9] ) );
  INV3 U712 ( .A(\u_decoder/fir_filter/dp_cluster_0/r178/CARRYB[7][2] ), .Q(
        n675) );
  INV3 U713 ( .A(\u_decoder/fir_filter/dp_cluster_0/r178/SUMB[7][3] ), .Q(n676) );
  NOR21 U714 ( .A(n685), .B(n686), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r177/A2[8] ) );
  INV3 U715 ( .A(\u_decoder/fir_filter/dp_cluster_0/r177/CARRYB[7][1] ), .Q(
        n685) );
  INV3 U716 ( .A(\u_decoder/fir_filter/dp_cluster_0/r177/SUMB[7][2] ), .Q(n686) );
  NOR21 U717 ( .A(n164), .B(n585), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[7][3] ) );
  INV3 U718 ( .A(\u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[6][3] ), .Q(
        n585) );
  NOR21 U719 ( .A(n165), .B(n646), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[7][3] ) );
  INV3 U720 ( .A(\u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[6][3] ), .Q(
        n646) );
  NOR21 U721 ( .A(n18), .B(n570), .Q(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[7][5] ) );
  INV3 U722 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[6][5] ), 
        .Q(n570) );
  NOR21 U723 ( .A(n19), .B(n631), .Q(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[7][5] ) );
  INV3 U724 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[6][5] ), 
        .Q(n631) );
  INV3 U725 ( .A(\u_decoder/iq_demod/dp_cluster_1/mult_150/ab[0][2] ), .Q(n720) );
  INV3 U726 ( .A(\u_decoder/iq_demod/dp_cluster_1/mult_150/ab[0][1] ), .Q(n718) );
  INV3 U727 ( .A(\u_decoder/iq_demod/dp_cluster_0/mult_148/ab[0][2] ), .Q(n708) );
  INV3 U728 ( .A(\u_decoder/iq_demod/dp_cluster_0/mult_148/ab[0][1] ), .Q(n706) );
  INV3 U729 ( .A(\u_decoder/iq_demod/dp_cluster_0/mult_151/ab[0][2] ), .Q(n696) );
  INV3 U730 ( .A(\u_decoder/iq_demod/dp_cluster_0/mult_151/ab[0][1] ), .Q(n694) );
  INV3 U731 ( .A(\u_decoder/iq_demod/dp_cluster_1/mult_149/ab[0][2] ), .Q(n732) );
  INV3 U732 ( .A(\u_decoder/iq_demod/dp_cluster_1/mult_149/ab[0][1] ), .Q(n730) );
  INV3 U733 ( .A(\u_decoder/iq_demod/dp_cluster_0/mult_151/ab[1][0] ), .Q(n695) );
  INV3 U734 ( .A(\u_decoder/iq_demod/dp_cluster_1/mult_150/ab[1][1] ), .Q(n721) );
  INV3 U735 ( .A(\u_decoder/iq_demod/dp_cluster_1/mult_150/ab[1][0] ), .Q(n719) );
  INV3 U736 ( .A(\u_decoder/iq_demod/dp_cluster_1/mult_149/ab[1][0] ), .Q(n731) );
  INV3 U737 ( .A(\u_decoder/iq_demod/dp_cluster_0/mult_148/ab[1][1] ), .Q(n709) );
  INV3 U738 ( .A(\u_decoder/iq_demod/dp_cluster_0/mult_148/ab[1][0] ), .Q(n707) );
  INV3 U739 ( .A(\u_decoder/iq_demod/dp_cluster_1/mult_150/ab[1][2] ), .Q(n723) );
  INV3 U740 ( .A(\u_decoder/iq_demod/dp_cluster_0/mult_148/ab[1][2] ), .Q(n711) );
  INV3 U741 ( .A(\u_decoder/iq_demod/dp_cluster_0/mult_151/ab[1][1] ), .Q(n697) );
  INV3 U742 ( .A(\u_decoder/iq_demod/dp_cluster_1/mult_149/ab[1][1] ), .Q(n733) );
  INV3 U743 ( .A(\u_decoder/iq_demod/dp_cluster_0/mult_151/ab[1][2] ), .Q(n699) );
  INV3 U744 ( .A(\u_decoder/iq_demod/dp_cluster_1/mult_149/ab[1][2] ), .Q(n735) );
  INV3 U745 ( .A(n2774), .Q(n2380) );
  AOI211 U746 ( .A(n2780), .B(\u_decoder/iq_demod/dp_cluster_0/mult_148/A1[4] ), .C(n2393), .Q(n2779) );
  INV3 U747 ( .A(n2781), .Q(n2393) );
  INV3 U748 ( .A(n2936), .Q(n2277) );
  INV3 U749 ( .A(n2850), .Q(n2348) );
  NAND22 U750 ( .A(n1219), .B(\u_coder/n139 ), .Q(\u_coder/n255 ) );
  NAND22 U751 ( .A(n1218), .B(\u_coder/n182 ), .Q(\u_coder/n239 ) );
  INV3 U752 ( .A(\u_coder/n281 ), .Q(n1916) );
  AOI221 U753 ( .A(\u_coder/n120 ), .B(n2169), .C(n890), .D(\u_coder/j [0]), 
        .Q(\u_coder/n281 ) );
  INV3 U754 ( .A(\u_coder/n278 ), .Q(n1919) );
  AOI221 U755 ( .A(\u_coder/N1016 ), .B(n2169), .C(\u_coder/n263 ), .D(
        \u_coder/j [3]), .Q(\u_coder/n278 ) );
  NOR21 U756 ( .A(n2902), .B(n2243), .Q(n2901) );
  AOI211 U757 ( .A(\u_decoder/fir_filter/dp_cluster_0/r165/A1[6] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r165/A2[6] ), .C(n2903), .Q(n2900)
         );
  NOR21 U758 ( .A(n2816), .B(n2314), .Q(n2815) );
  AOI211 U759 ( .A(\u_decoder/fir_filter/dp_cluster_0/r178/A1[6] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r178/A2[6] ), .C(n2817), .Q(n2814)
         );
  NOR21 U760 ( .A(n736), .B(n737), .Q(
        \u_decoder/iq_demod/dp_cluster_1/add_154/carry [1]) );
  XOR21 U761 ( .A(\u_decoder/iq_demod/dp_cluster_1/mult_149/ab[0][1] ), .B(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/ab[1][0] ), .Q(
        \u_decoder/iq_demod/dp_cluster_1/mult_I_sin_out [1]) );
  XOR21 U762 ( .A(\u_decoder/iq_demod/dp_cluster_1/mult_150/ab[0][1] ), .B(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/ab[1][0] ), .Q(
        \u_decoder/iq_demod/dp_cluster_1/mult_Q_cos_out [1]) );
  INV3 U763 ( .A(n477), .Q(\u_decoder/iq_demod/dp_cluster_0/sub_153/carry [1])
         );
  XOR21 U764 ( .A(\u_decoder/iq_demod/dp_cluster_0/mult_148/ab[0][1] ), .B(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/ab[1][0] ), .Q(
        \u_decoder/iq_demod/dp_cluster_0/mult_I_cos_out [1]) );
  INV3 U765 ( .A(\u_decoder/iq_demod/dp_cluster_0/mult_Q_sin_out [2]), .Q(
        n2388) );
  NOR21 U766 ( .A(n592), .B(n593), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r167/A2[10] ) );
  INV3 U767 ( .A(\u_decoder/fir_filter/dp_cluster_0/r167/SUMB[7][4] ), .Q(n593) );
  INV3 U768 ( .A(\u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[7][3] ), .Q(
        n592) );
  NOR21 U769 ( .A(n653), .B(n654), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r180/A2[10] ) );
  INV3 U770 ( .A(\u_decoder/fir_filter/dp_cluster_0/r180/SUMB[7][4] ), .Q(n654) );
  INV3 U771 ( .A(\u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[7][3] ), .Q(
        n653) );
  INV3 U772 ( .A(\u_coder/n135 ), .Q(n1809) );
  INV3 U773 ( .A(\u_inFIFO/N375 ), .Q(n2143) );
  NOR21 U774 ( .A(n2383), .B(
        \u_decoder/iq_demod/dp_cluster_0/mult_I_cos_out [0]), .Q(n477) );
  NOR21 U775 ( .A(n616), .B(n617), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r165/A2[10] ) );
  INV3 U776 ( .A(\u_decoder/fir_filter/dp_cluster_0/r165/SUMB[7][4] ), .Q(n617) );
  INV3 U777 ( .A(\u_decoder/fir_filter/dp_cluster_0/r165/CARRYB[7][3] ), .Q(
        n616) );
  NOR21 U778 ( .A(n677), .B(n678), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r178/A2[10] ) );
  INV3 U779 ( .A(\u_decoder/fir_filter/dp_cluster_0/r178/SUMB[7][4] ), .Q(n678) );
  INV3 U780 ( .A(\u_decoder/fir_filter/dp_cluster_0/r178/CARRYB[7][3] ), .Q(
        n677) );
  NOR21 U781 ( .A(n626), .B(n617), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r164/A2[9] ) );
  INV3 U782 ( .A(\u_decoder/fir_filter/dp_cluster_0/r164/CARRYB[7][2] ), .Q(
        n626) );
  NOR21 U783 ( .A(n687), .B(n678), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r177/A2[9] ) );
  INV3 U784 ( .A(\u_decoder/fir_filter/dp_cluster_0/r177/CARRYB[7][2] ), .Q(
        n687) );
  INV3 U785 ( .A(\u_decoder/fir_filter/I_data_mult_2[8] ), .Q(n2250) );
  AOI211 U786 ( .A(\u_decoder/fir_filter/dp_cluster_0/r166/A1[6] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r166/A2[6] ), .C(n2914), .Q(
        \u_decoder/fir_filter/I_data_mult_2[8] ) );
  NOR21 U787 ( .A(\u_decoder/fir_filter/dp_cluster_0/r166/A2[6] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r166/A1[6] ), .Q(n2914) );
  INV3 U788 ( .A(\u_decoder/fir_filter/Q_data_mult_2[8] ), .Q(n2321) );
  AOI211 U789 ( .A(\u_decoder/fir_filter/dp_cluster_0/r179/A1[6] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r179/A2[6] ), .C(n2828), .Q(
        \u_decoder/fir_filter/Q_data_mult_2[8] ) );
  NOR21 U790 ( .A(\u_decoder/fir_filter/dp_cluster_0/r179/A2[6] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r179/A1[6] ), .Q(n2828) );
  INV3 U791 ( .A(\u_decoder/fir_filter/I_data_mult_3 [8]), .Q(n2283) );
  AOI211 U792 ( .A(n363), .B(n321), .C(n2929), .Q(
        \u_decoder/fir_filter/I_data_mult_3 [8]) );
  INV3 U793 ( .A(\u_decoder/fir_filter/Q_data_mult_3 [8]), .Q(n2354) );
  AOI211 U794 ( .A(n364), .B(n322), .C(n2843), .Q(
        \u_decoder/fir_filter/Q_data_mult_3 [8]) );
  INV3 U795 ( .A(\u_coder/n182 ), .Q(n2102) );
  NOR21 U796 ( .A(n18), .B(n598), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r166/CARRYB[7][3] ) );
  INV3 U797 ( .A(\u_decoder/fir_filter/dp_cluster_0/r166/CARRYB[6][3] ), .Q(
        n598) );
  NOR21 U798 ( .A(n19), .B(n659), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r179/CARRYB[7][3] ) );
  INV3 U799 ( .A(\u_decoder/fir_filter/dp_cluster_0/r179/CARRYB[6][3] ), .Q(
        n659) );
  INV3 U800 ( .A(\u_decoder/iq_demod/dp_cluster_1/mult_Q_cos_out [0]), .Q(n736) );
  INV3 U801 ( .A(\u_decoder/iq_demod/dp_cluster_1/mult_I_sin_out [0]), .Q(n737) );
  NAND22 U802 ( .A(n1219), .B(n1209), .Q(\u_inFIFO/n224 ) );
  NOR21 U803 ( .A(n1203), .B(n2146), .Q(\u_inFIFO/n513 ) );
  XOR21 U804 ( .A(\u_decoder/fir_filter/dp_cluster_0/r167/SUMB[7][5] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[7][4] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r167/A1[10] ) );
  XOR21 U805 ( .A(\u_decoder/fir_filter/dp_cluster_0/r180/SUMB[7][5] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[7][4] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r180/A1[10] ) );
  NAND22 U806 ( .A(n2168), .B(\u_coder/n251 ), .Q(\u_coder/n167 ) );
  NOR21 U807 ( .A(\u_coder/n212 ), .B(\u_coder/n218 ), .Q(\u_coder/n194 ) );
  NAND22 U808 ( .A(n1219), .B(n1191), .Q(\u_outFIFO/n1112 ) );
  INV3 U809 ( .A(\u_inFIFO/n231 ), .Q(n2091) );
  NOR21 U810 ( .A(n897), .B(\u_inFIFO/n233 ), .Q(\u_inFIFO/n232 ) );
  INV3 U811 ( .A(\u_inFIFO/n228 ), .Q(n2092) );
  NOR21 U812 ( .A(n897), .B(\u_inFIFO/n230 ), .Q(\u_inFIFO/n229 ) );
  BUF2 U813 ( .A(\u_decoder/fir_filter/n721 ), .Q(n1167) );
  BUF2 U814 ( .A(n1795), .Q(n952) );
  BUF2 U815 ( .A(n1795), .Q(n953) );
  BUF2 U816 ( .A(n1795), .Q(n954) );
  BUF2 U817 ( .A(n1795), .Q(n955) );
  BUF2 U818 ( .A(n1795), .Q(n956) );
  BUF2 U819 ( .A(n1795), .Q(n957) );
  BUF2 U820 ( .A(n1795), .Q(n958) );
  BUF2 U821 ( .A(n1795), .Q(n959) );
  BUF2 U822 ( .A(n1795), .Q(n960) );
  BUF2 U823 ( .A(n1795), .Q(n961) );
  INV3 U824 ( .A(\u_outFIFO/n660 ), .Q(n1191) );
  XOR21 U825 ( .A(n2902), .B(\u_decoder/fir_filter/dp_cluster_0/r165/A1[5] ), 
        .Q(n351) );
  XOR21 U826 ( .A(n2816), .B(\u_decoder/fir_filter/dp_cluster_0/r178/A1[5] ), 
        .Q(n352) );
  NAND22 U827 ( .A(n1219), .B(\u_coder/n167 ), .Q(\u_coder/n254 ) );
  NOR21 U828 ( .A(n594), .B(n595), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r167/A2[11] ) );
  INV3 U829 ( .A(\u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[7][4] ), .Q(
        n594) );
  INV3 U830 ( .A(\u_decoder/fir_filter/dp_cluster_0/r167/SUMB[7][5] ), .Q(n595) );
  NOR21 U831 ( .A(n655), .B(n656), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r180/A2[11] ) );
  INV3 U832 ( .A(\u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[7][4] ), .Q(
        n655) );
  INV3 U833 ( .A(\u_decoder/fir_filter/dp_cluster_0/r180/SUMB[7][5] ), .Q(n656) );
  INV3 U834 ( .A(\u_coder/n176 ), .Q(n2155) );
  NOR21 U835 ( .A(\u_coder/n169 ), .B(n2162), .Q(\u_coder/n176 ) );
  BUF2 U836 ( .A(\u_decoder/fir_filter/n554 ), .Q(n1145) );
  BUF2 U837 ( .A(\u_decoder/fir_filter/n554 ), .Q(n1148) );
  BUF2 U838 ( .A(\u_decoder/fir_filter/n554 ), .Q(n1146) );
  BUF2 U839 ( .A(\u_decoder/fir_filter/n554 ), .Q(n1147) );
  INV3 U840 ( .A(\u_coder/n309 ), .Q(n2161) );
  BUF2 U841 ( .A(\u_outFIFO/n545 ), .Q(n804) );
  BUF2 U842 ( .A(\u_outFIFO/n545 ), .Q(n805) );
  INV3 U843 ( .A(\u_coder/n251 ), .Q(n2162) );
  INV3 U844 ( .A(\u_inFIFO/n510 ), .Q(n1966) );
  NOR21 U845 ( .A(\u_inFIFO/n272 ), .B(n910), .Q(\u_inFIFO/n511 ) );
  INV3 U846 ( .A(\u_inFIFO/n508 ), .Q(n1967) );
  NOR21 U847 ( .A(\u_inFIFO/n269 ), .B(n910), .Q(\u_inFIFO/n509 ) );
  INV3 U848 ( .A(\u_inFIFO/n506 ), .Q(n1968) );
  NOR21 U849 ( .A(\u_inFIFO/n266 ), .B(n910), .Q(\u_inFIFO/n507 ) );
  INV3 U850 ( .A(\u_inFIFO/n503 ), .Q(n1969) );
  NOR21 U851 ( .A(\u_inFIFO/n263 ), .B(n910), .Q(\u_inFIFO/n504 ) );
  INV3 U852 ( .A(\u_inFIFO/n501 ), .Q(n1970) );
  NOR21 U853 ( .A(\u_inFIFO/n260 ), .B(n910), .Q(\u_inFIFO/n502 ) );
  INV3 U854 ( .A(\u_inFIFO/n499 ), .Q(n1971) );
  NOR21 U855 ( .A(\u_inFIFO/n257 ), .B(n910), .Q(\u_inFIFO/n500 ) );
  INV3 U856 ( .A(\u_inFIFO/n497 ), .Q(n1972) );
  NOR21 U857 ( .A(\u_inFIFO/n254 ), .B(n910), .Q(\u_inFIFO/n498 ) );
  INV3 U858 ( .A(\u_inFIFO/n494 ), .Q(n1973) );
  NOR21 U859 ( .A(\u_inFIFO/n251 ), .B(n910), .Q(\u_inFIFO/n495 ) );
  INV3 U860 ( .A(\u_inFIFO/n492 ), .Q(n1974) );
  NOR21 U861 ( .A(\u_inFIFO/n248 ), .B(n911), .Q(\u_inFIFO/n493 ) );
  INV3 U862 ( .A(\u_inFIFO/n490 ), .Q(n1975) );
  NOR21 U863 ( .A(\u_inFIFO/n245 ), .B(n911), .Q(\u_inFIFO/n491 ) );
  INV3 U864 ( .A(\u_inFIFO/n488 ), .Q(n1976) );
  NOR21 U865 ( .A(\u_inFIFO/n242 ), .B(n911), .Q(\u_inFIFO/n489 ) );
  INV3 U866 ( .A(\u_inFIFO/n485 ), .Q(n1977) );
  NOR21 U867 ( .A(\u_inFIFO/n239 ), .B(n911), .Q(\u_inFIFO/n486 ) );
  INV3 U868 ( .A(\u_inFIFO/n482 ), .Q(n1978) );
  NOR21 U869 ( .A(\u_inFIFO/n236 ), .B(n911), .Q(\u_inFIFO/n483 ) );
  INV3 U870 ( .A(\u_inFIFO/n479 ), .Q(n1979) );
  NOR21 U871 ( .A(\u_inFIFO/n233 ), .B(n911), .Q(\u_inFIFO/n480 ) );
  INV3 U872 ( .A(\u_inFIFO/n476 ), .Q(n1980) );
  NOR21 U873 ( .A(\u_inFIFO/n230 ), .B(n911), .Q(\u_inFIFO/n477 ) );
  INV3 U874 ( .A(\u_inFIFO/n471 ), .Q(n1981) );
  NOR21 U875 ( .A(\u_inFIFO/n226 ), .B(n911), .Q(\u_inFIFO/n472 ) );
  INV3 U876 ( .A(\u_inFIFO/n469 ), .Q(n1982) );
  NOR21 U877 ( .A(\u_inFIFO/n272 ), .B(n908), .Q(\u_inFIFO/n470 ) );
  INV3 U878 ( .A(\u_inFIFO/n467 ), .Q(n1983) );
  NOR21 U879 ( .A(\u_inFIFO/n269 ), .B(n908), .Q(\u_inFIFO/n468 ) );
  INV3 U880 ( .A(\u_inFIFO/n465 ), .Q(n1984) );
  NOR21 U881 ( .A(\u_inFIFO/n266 ), .B(n908), .Q(\u_inFIFO/n466 ) );
  INV3 U882 ( .A(\u_inFIFO/n463 ), .Q(n1985) );
  NOR21 U883 ( .A(\u_inFIFO/n263 ), .B(n908), .Q(\u_inFIFO/n464 ) );
  INV3 U884 ( .A(\u_inFIFO/n461 ), .Q(n1986) );
  NOR21 U885 ( .A(\u_inFIFO/n260 ), .B(n908), .Q(\u_inFIFO/n462 ) );
  INV3 U886 ( .A(\u_inFIFO/n459 ), .Q(n1987) );
  NOR21 U887 ( .A(\u_inFIFO/n257 ), .B(n908), .Q(\u_inFIFO/n460 ) );
  INV3 U888 ( .A(\u_inFIFO/n457 ), .Q(n1988) );
  NOR21 U889 ( .A(\u_inFIFO/n254 ), .B(n908), .Q(\u_inFIFO/n458 ) );
  INV3 U890 ( .A(\u_inFIFO/n455 ), .Q(n1989) );
  NOR21 U891 ( .A(\u_inFIFO/n251 ), .B(n908), .Q(\u_inFIFO/n456 ) );
  INV3 U892 ( .A(\u_inFIFO/n453 ), .Q(n1990) );
  NOR21 U893 ( .A(\u_inFIFO/n248 ), .B(n909), .Q(\u_inFIFO/n454 ) );
  INV3 U894 ( .A(\u_inFIFO/n451 ), .Q(n1991) );
  NOR21 U895 ( .A(\u_inFIFO/n245 ), .B(n909), .Q(\u_inFIFO/n452 ) );
  INV3 U896 ( .A(\u_inFIFO/n449 ), .Q(n1992) );
  NOR21 U897 ( .A(\u_inFIFO/n242 ), .B(n909), .Q(\u_inFIFO/n450 ) );
  INV3 U898 ( .A(\u_inFIFO/n447 ), .Q(n1993) );
  NOR21 U899 ( .A(\u_inFIFO/n239 ), .B(n909), .Q(\u_inFIFO/n448 ) );
  INV3 U900 ( .A(\u_inFIFO/n445 ), .Q(n1994) );
  NOR21 U901 ( .A(\u_inFIFO/n236 ), .B(n909), .Q(\u_inFIFO/n446 ) );
  INV3 U902 ( .A(\u_inFIFO/n443 ), .Q(n1995) );
  NOR21 U903 ( .A(\u_inFIFO/n233 ), .B(n909), .Q(\u_inFIFO/n444 ) );
  INV3 U904 ( .A(\u_inFIFO/n441 ), .Q(n1996) );
  NOR21 U905 ( .A(\u_inFIFO/n230 ), .B(n909), .Q(\u_inFIFO/n442 ) );
  INV3 U906 ( .A(\u_inFIFO/n438 ), .Q(n1997) );
  NOR21 U907 ( .A(\u_inFIFO/n226 ), .B(n909), .Q(\u_inFIFO/n439 ) );
  INV3 U908 ( .A(\u_inFIFO/n436 ), .Q(n1998) );
  NOR21 U909 ( .A(\u_inFIFO/n272 ), .B(n906), .Q(\u_inFIFO/n437 ) );
  INV3 U910 ( .A(\u_inFIFO/n434 ), .Q(n1999) );
  NOR21 U911 ( .A(\u_inFIFO/n269 ), .B(n906), .Q(\u_inFIFO/n435 ) );
  INV3 U912 ( .A(\u_inFIFO/n432 ), .Q(n2000) );
  NOR21 U913 ( .A(\u_inFIFO/n266 ), .B(n906), .Q(\u_inFIFO/n433 ) );
  INV3 U914 ( .A(\u_inFIFO/n430 ), .Q(n2001) );
  NOR21 U915 ( .A(\u_inFIFO/n263 ), .B(n906), .Q(\u_inFIFO/n431 ) );
  INV3 U916 ( .A(\u_inFIFO/n428 ), .Q(n2002) );
  NOR21 U917 ( .A(\u_inFIFO/n260 ), .B(n906), .Q(\u_inFIFO/n429 ) );
  INV3 U918 ( .A(\u_inFIFO/n426 ), .Q(n2003) );
  NOR21 U919 ( .A(\u_inFIFO/n257 ), .B(n906), .Q(\u_inFIFO/n427 ) );
  INV3 U920 ( .A(\u_inFIFO/n424 ), .Q(n2004) );
  NOR21 U921 ( .A(\u_inFIFO/n254 ), .B(n906), .Q(\u_inFIFO/n425 ) );
  INV3 U922 ( .A(\u_inFIFO/n422 ), .Q(n2005) );
  NOR21 U923 ( .A(\u_inFIFO/n251 ), .B(n906), .Q(\u_inFIFO/n423 ) );
  INV3 U924 ( .A(\u_inFIFO/n420 ), .Q(n2006) );
  NOR21 U925 ( .A(\u_inFIFO/n248 ), .B(n907), .Q(\u_inFIFO/n421 ) );
  INV3 U926 ( .A(\u_inFIFO/n418 ), .Q(n2007) );
  NOR21 U927 ( .A(\u_inFIFO/n245 ), .B(n907), .Q(\u_inFIFO/n419 ) );
  INV3 U928 ( .A(\u_inFIFO/n416 ), .Q(n2008) );
  NOR21 U929 ( .A(\u_inFIFO/n242 ), .B(n907), .Q(\u_inFIFO/n417 ) );
  INV3 U930 ( .A(\u_inFIFO/n414 ), .Q(n2009) );
  NOR21 U931 ( .A(\u_inFIFO/n239 ), .B(n907), .Q(\u_inFIFO/n415 ) );
  INV3 U932 ( .A(\u_inFIFO/n412 ), .Q(n2010) );
  NOR21 U933 ( .A(\u_inFIFO/n236 ), .B(n907), .Q(\u_inFIFO/n413 ) );
  INV3 U934 ( .A(\u_inFIFO/n410 ), .Q(n2011) );
  NOR21 U935 ( .A(\u_inFIFO/n233 ), .B(n907), .Q(\u_inFIFO/n411 ) );
  INV3 U936 ( .A(\u_inFIFO/n408 ), .Q(n2012) );
  NOR21 U937 ( .A(\u_inFIFO/n230 ), .B(n907), .Q(\u_inFIFO/n409 ) );
  INV3 U938 ( .A(\u_inFIFO/n405 ), .Q(n2013) );
  NOR21 U939 ( .A(\u_inFIFO/n226 ), .B(n907), .Q(\u_inFIFO/n406 ) );
  INV3 U940 ( .A(\u_inFIFO/n403 ), .Q(n2014) );
  NOR21 U941 ( .A(\u_inFIFO/n272 ), .B(n904), .Q(\u_inFIFO/n404 ) );
  INV3 U942 ( .A(\u_inFIFO/n401 ), .Q(n2015) );
  NOR21 U943 ( .A(\u_inFIFO/n269 ), .B(n904), .Q(\u_inFIFO/n402 ) );
  INV3 U944 ( .A(\u_inFIFO/n399 ), .Q(n2016) );
  NOR21 U945 ( .A(\u_inFIFO/n266 ), .B(n904), .Q(\u_inFIFO/n400 ) );
  INV3 U946 ( .A(\u_inFIFO/n397 ), .Q(n2017) );
  NOR21 U947 ( .A(\u_inFIFO/n263 ), .B(n904), .Q(\u_inFIFO/n398 ) );
  INV3 U948 ( .A(\u_inFIFO/n395 ), .Q(n2018) );
  NOR21 U949 ( .A(\u_inFIFO/n260 ), .B(n904), .Q(\u_inFIFO/n396 ) );
  INV3 U950 ( .A(\u_inFIFO/n393 ), .Q(n2019) );
  NOR21 U951 ( .A(\u_inFIFO/n257 ), .B(n904), .Q(\u_inFIFO/n394 ) );
  INV3 U952 ( .A(\u_inFIFO/n391 ), .Q(n2020) );
  NOR21 U953 ( .A(\u_inFIFO/n254 ), .B(n904), .Q(\u_inFIFO/n392 ) );
  INV3 U954 ( .A(\u_inFIFO/n389 ), .Q(n2021) );
  NOR21 U955 ( .A(\u_inFIFO/n251 ), .B(n904), .Q(\u_inFIFO/n390 ) );
  INV3 U956 ( .A(\u_inFIFO/n387 ), .Q(n2022) );
  NOR21 U957 ( .A(\u_inFIFO/n248 ), .B(n905), .Q(\u_inFIFO/n388 ) );
  INV3 U958 ( .A(\u_inFIFO/n385 ), .Q(n2023) );
  NOR21 U959 ( .A(\u_inFIFO/n245 ), .B(n905), .Q(\u_inFIFO/n386 ) );
  INV3 U960 ( .A(\u_inFIFO/n383 ), .Q(n2024) );
  NOR21 U961 ( .A(\u_inFIFO/n242 ), .B(n905), .Q(\u_inFIFO/n384 ) );
  INV3 U962 ( .A(\u_inFIFO/n381 ), .Q(n2025) );
  NOR21 U963 ( .A(\u_inFIFO/n239 ), .B(n905), .Q(\u_inFIFO/n382 ) );
  INV3 U964 ( .A(\u_inFIFO/n379 ), .Q(n2026) );
  NOR21 U965 ( .A(\u_inFIFO/n236 ), .B(n905), .Q(\u_inFIFO/n380 ) );
  INV3 U966 ( .A(\u_inFIFO/n377 ), .Q(n2027) );
  NOR21 U967 ( .A(\u_inFIFO/n233 ), .B(n905), .Q(\u_inFIFO/n378 ) );
  INV3 U968 ( .A(\u_inFIFO/n375 ), .Q(n2028) );
  NOR21 U969 ( .A(\u_inFIFO/n230 ), .B(n905), .Q(\u_inFIFO/n376 ) );
  INV3 U970 ( .A(\u_inFIFO/n372 ), .Q(n2029) );
  NOR21 U971 ( .A(\u_inFIFO/n226 ), .B(n905), .Q(\u_inFIFO/n373 ) );
  INV3 U972 ( .A(\u_inFIFO/n370 ), .Q(n2030) );
  NOR21 U973 ( .A(\u_inFIFO/n272 ), .B(n902), .Q(\u_inFIFO/n371 ) );
  INV3 U974 ( .A(\u_inFIFO/n368 ), .Q(n2031) );
  NOR21 U975 ( .A(\u_inFIFO/n269 ), .B(n902), .Q(\u_inFIFO/n369 ) );
  INV3 U976 ( .A(\u_inFIFO/n366 ), .Q(n2032) );
  NOR21 U977 ( .A(\u_inFIFO/n266 ), .B(n902), .Q(\u_inFIFO/n367 ) );
  INV3 U978 ( .A(\u_inFIFO/n364 ), .Q(n2033) );
  NOR21 U979 ( .A(\u_inFIFO/n263 ), .B(n902), .Q(\u_inFIFO/n365 ) );
  INV3 U980 ( .A(\u_inFIFO/n362 ), .Q(n2034) );
  NOR21 U981 ( .A(\u_inFIFO/n260 ), .B(n902), .Q(\u_inFIFO/n363 ) );
  INV3 U982 ( .A(\u_inFIFO/n360 ), .Q(n2035) );
  NOR21 U983 ( .A(\u_inFIFO/n257 ), .B(n902), .Q(\u_inFIFO/n361 ) );
  INV3 U984 ( .A(\u_inFIFO/n358 ), .Q(n2036) );
  NOR21 U985 ( .A(\u_inFIFO/n254 ), .B(n902), .Q(\u_inFIFO/n359 ) );
  INV3 U986 ( .A(\u_inFIFO/n356 ), .Q(n2037) );
  NOR21 U987 ( .A(\u_inFIFO/n251 ), .B(n902), .Q(\u_inFIFO/n357 ) );
  INV3 U988 ( .A(\u_inFIFO/n354 ), .Q(n2038) );
  NOR21 U989 ( .A(\u_inFIFO/n248 ), .B(n903), .Q(\u_inFIFO/n355 ) );
  INV3 U990 ( .A(\u_inFIFO/n352 ), .Q(n2039) );
  NOR21 U991 ( .A(\u_inFIFO/n245 ), .B(n903), .Q(\u_inFIFO/n353 ) );
  INV3 U992 ( .A(\u_inFIFO/n350 ), .Q(n2040) );
  NOR21 U993 ( .A(\u_inFIFO/n242 ), .B(n903), .Q(\u_inFIFO/n351 ) );
  INV3 U994 ( .A(\u_inFIFO/n348 ), .Q(n2041) );
  NOR21 U995 ( .A(\u_inFIFO/n239 ), .B(n903), .Q(\u_inFIFO/n349 ) );
  INV3 U996 ( .A(\u_inFIFO/n346 ), .Q(n2042) );
  NOR21 U997 ( .A(\u_inFIFO/n236 ), .B(n903), .Q(\u_inFIFO/n347 ) );
  INV3 U998 ( .A(\u_inFIFO/n344 ), .Q(n2043) );
  NOR21 U999 ( .A(\u_inFIFO/n233 ), .B(n903), .Q(\u_inFIFO/n345 ) );
  INV3 U1000 ( .A(\u_inFIFO/n342 ), .Q(n2044) );
  NOR21 U1001 ( .A(\u_inFIFO/n230 ), .B(n903), .Q(\u_inFIFO/n343 ) );
  INV3 U1002 ( .A(\u_inFIFO/n339 ), .Q(n2045) );
  NOR21 U1003 ( .A(\u_inFIFO/n226 ), .B(n903), .Q(\u_inFIFO/n340 ) );
  INV3 U1004 ( .A(\u_inFIFO/n337 ), .Q(n2046) );
  NOR21 U1005 ( .A(\u_inFIFO/n272 ), .B(n900), .Q(\u_inFIFO/n338 ) );
  INV3 U1006 ( .A(\u_inFIFO/n335 ), .Q(n2047) );
  NOR21 U1007 ( .A(\u_inFIFO/n269 ), .B(n900), .Q(\u_inFIFO/n336 ) );
  INV3 U1008 ( .A(\u_inFIFO/n333 ), .Q(n2048) );
  NOR21 U1009 ( .A(\u_inFIFO/n266 ), .B(n900), .Q(\u_inFIFO/n334 ) );
  INV3 U1010 ( .A(\u_inFIFO/n331 ), .Q(n2049) );
  NOR21 U1011 ( .A(\u_inFIFO/n263 ), .B(n900), .Q(\u_inFIFO/n332 ) );
  INV3 U1012 ( .A(\u_inFIFO/n329 ), .Q(n2050) );
  NOR21 U1013 ( .A(\u_inFIFO/n260 ), .B(n900), .Q(\u_inFIFO/n330 ) );
  INV3 U1014 ( .A(\u_inFIFO/n327 ), .Q(n2051) );
  NOR21 U1015 ( .A(\u_inFIFO/n257 ), .B(n900), .Q(\u_inFIFO/n328 ) );
  INV3 U1016 ( .A(\u_inFIFO/n325 ), .Q(n2052) );
  NOR21 U1017 ( .A(\u_inFIFO/n254 ), .B(n900), .Q(\u_inFIFO/n326 ) );
  INV3 U1018 ( .A(\u_inFIFO/n323 ), .Q(n2053) );
  NOR21 U1019 ( .A(\u_inFIFO/n251 ), .B(n900), .Q(\u_inFIFO/n324 ) );
  INV3 U1020 ( .A(\u_inFIFO/n321 ), .Q(n2054) );
  NOR21 U1021 ( .A(\u_inFIFO/n248 ), .B(n901), .Q(\u_inFIFO/n322 ) );
  INV3 U1022 ( .A(\u_inFIFO/n319 ), .Q(n2055) );
  NOR21 U1023 ( .A(\u_inFIFO/n245 ), .B(n901), .Q(\u_inFIFO/n320 ) );
  INV3 U1024 ( .A(\u_inFIFO/n317 ), .Q(n2056) );
  NOR21 U1025 ( .A(\u_inFIFO/n242 ), .B(n901), .Q(\u_inFIFO/n318 ) );
  INV3 U1026 ( .A(\u_inFIFO/n315 ), .Q(n2057) );
  NOR21 U1027 ( .A(\u_inFIFO/n239 ), .B(n901), .Q(\u_inFIFO/n316 ) );
  INV3 U1028 ( .A(\u_inFIFO/n313 ), .Q(n2058) );
  NOR21 U1029 ( .A(\u_inFIFO/n236 ), .B(n901), .Q(\u_inFIFO/n314 ) );
  INV3 U1030 ( .A(\u_inFIFO/n311 ), .Q(n2059) );
  NOR21 U1031 ( .A(\u_inFIFO/n233 ), .B(n901), .Q(\u_inFIFO/n312 ) );
  INV3 U1032 ( .A(\u_inFIFO/n309 ), .Q(n2060) );
  NOR21 U1033 ( .A(\u_inFIFO/n230 ), .B(n901), .Q(\u_inFIFO/n310 ) );
  INV3 U1034 ( .A(\u_inFIFO/n306 ), .Q(n2061) );
  NOR21 U1035 ( .A(\u_inFIFO/n226 ), .B(n901), .Q(\u_inFIFO/n307 ) );
  INV3 U1036 ( .A(\u_inFIFO/n304 ), .Q(n2062) );
  NOR21 U1037 ( .A(\u_inFIFO/n272 ), .B(n898), .Q(\u_inFIFO/n305 ) );
  INV3 U1038 ( .A(\u_inFIFO/n302 ), .Q(n2063) );
  NOR21 U1039 ( .A(\u_inFIFO/n269 ), .B(n898), .Q(\u_inFIFO/n303 ) );
  INV3 U1040 ( .A(\u_inFIFO/n300 ), .Q(n2064) );
  NOR21 U1041 ( .A(\u_inFIFO/n266 ), .B(n898), .Q(\u_inFIFO/n301 ) );
  INV3 U1042 ( .A(\u_inFIFO/n298 ), .Q(n2065) );
  NOR21 U1043 ( .A(\u_inFIFO/n263 ), .B(n898), .Q(\u_inFIFO/n299 ) );
  INV3 U1044 ( .A(\u_inFIFO/n296 ), .Q(n2066) );
  NOR21 U1045 ( .A(\u_inFIFO/n260 ), .B(n898), .Q(\u_inFIFO/n297 ) );
  INV3 U1046 ( .A(\u_inFIFO/n294 ), .Q(n2067) );
  NOR21 U1047 ( .A(\u_inFIFO/n257 ), .B(n898), .Q(\u_inFIFO/n295 ) );
  INV3 U1048 ( .A(\u_inFIFO/n292 ), .Q(n2068) );
  NOR21 U1049 ( .A(\u_inFIFO/n254 ), .B(n898), .Q(\u_inFIFO/n293 ) );
  INV3 U1050 ( .A(\u_inFIFO/n290 ), .Q(n2069) );
  NOR21 U1051 ( .A(\u_inFIFO/n251 ), .B(n898), .Q(\u_inFIFO/n291 ) );
  INV3 U1052 ( .A(\u_inFIFO/n288 ), .Q(n2070) );
  NOR21 U1053 ( .A(\u_inFIFO/n248 ), .B(n899), .Q(\u_inFIFO/n289 ) );
  INV3 U1054 ( .A(\u_inFIFO/n286 ), .Q(n2071) );
  NOR21 U1055 ( .A(\u_inFIFO/n245 ), .B(n899), .Q(\u_inFIFO/n287 ) );
  INV3 U1056 ( .A(\u_inFIFO/n284 ), .Q(n2072) );
  NOR21 U1057 ( .A(\u_inFIFO/n242 ), .B(n899), .Q(\u_inFIFO/n285 ) );
  INV3 U1058 ( .A(\u_inFIFO/n282 ), .Q(n2073) );
  NOR21 U1059 ( .A(\u_inFIFO/n239 ), .B(n899), .Q(\u_inFIFO/n283 ) );
  INV3 U1060 ( .A(\u_inFIFO/n280 ), .Q(n2074) );
  NOR21 U1061 ( .A(\u_inFIFO/n236 ), .B(n899), .Q(\u_inFIFO/n281 ) );
  INV3 U1062 ( .A(\u_inFIFO/n278 ), .Q(n2075) );
  NOR21 U1063 ( .A(\u_inFIFO/n233 ), .B(n899), .Q(\u_inFIFO/n279 ) );
  INV3 U1064 ( .A(\u_inFIFO/n276 ), .Q(n2076) );
  NOR21 U1065 ( .A(\u_inFIFO/n230 ), .B(n899), .Q(\u_inFIFO/n277 ) );
  INV3 U1066 ( .A(\u_inFIFO/n273 ), .Q(n2077) );
  NOR21 U1067 ( .A(\u_inFIFO/n226 ), .B(n899), .Q(\u_inFIFO/n274 ) );
  INV3 U1068 ( .A(\u_inFIFO/n270 ), .Q(n2078) );
  NOR21 U1069 ( .A(n896), .B(\u_inFIFO/n272 ), .Q(\u_inFIFO/n271 ) );
  INV3 U1070 ( .A(\u_inFIFO/n267 ), .Q(n2079) );
  NOR21 U1071 ( .A(n896), .B(\u_inFIFO/n269 ), .Q(\u_inFIFO/n268 ) );
  INV3 U1072 ( .A(\u_inFIFO/n264 ), .Q(n2080) );
  NOR21 U1073 ( .A(n896), .B(\u_inFIFO/n266 ), .Q(\u_inFIFO/n265 ) );
  INV3 U1074 ( .A(\u_inFIFO/n261 ), .Q(n2081) );
  NOR21 U1075 ( .A(n896), .B(\u_inFIFO/n263 ), .Q(\u_inFIFO/n262 ) );
  INV3 U1076 ( .A(\u_inFIFO/n258 ), .Q(n2082) );
  NOR21 U1077 ( .A(n896), .B(\u_inFIFO/n260 ), .Q(\u_inFIFO/n259 ) );
  INV3 U1078 ( .A(\u_inFIFO/n255 ), .Q(n2083) );
  NOR21 U1079 ( .A(n896), .B(\u_inFIFO/n257 ), .Q(\u_inFIFO/n256 ) );
  INV3 U1080 ( .A(\u_inFIFO/n252 ), .Q(n2084) );
  NOR21 U1081 ( .A(n896), .B(\u_inFIFO/n254 ), .Q(\u_inFIFO/n253 ) );
  INV3 U1082 ( .A(\u_inFIFO/n249 ), .Q(n2085) );
  NOR21 U1083 ( .A(n896), .B(\u_inFIFO/n251 ), .Q(\u_inFIFO/n250 ) );
  INV3 U1084 ( .A(\u_inFIFO/n246 ), .Q(n2086) );
  NOR21 U1085 ( .A(n897), .B(\u_inFIFO/n248 ), .Q(\u_inFIFO/n247 ) );
  INV3 U1086 ( .A(\u_inFIFO/n243 ), .Q(n2087) );
  NOR21 U1087 ( .A(n897), .B(\u_inFIFO/n245 ), .Q(\u_inFIFO/n244 ) );
  INV3 U1088 ( .A(\u_inFIFO/n240 ), .Q(n2088) );
  NOR21 U1089 ( .A(n897), .B(\u_inFIFO/n242 ), .Q(\u_inFIFO/n241 ) );
  INV3 U1090 ( .A(\u_inFIFO/n237 ), .Q(n2089) );
  NOR21 U1091 ( .A(n897), .B(\u_inFIFO/n239 ), .Q(\u_inFIFO/n238 ) );
  INV3 U1092 ( .A(\u_inFIFO/n234 ), .Q(n2090) );
  NOR21 U1093 ( .A(n897), .B(\u_inFIFO/n236 ), .Q(\u_inFIFO/n235 ) );
  INV3 U1094 ( .A(\u_inFIFO/n218 ), .Q(n2093) );
  NOR21 U1095 ( .A(\u_inFIFO/n226 ), .B(n897), .Q(\u_inFIFO/n223 ) );
  BUF2 U1096 ( .A(\u_decoder/fir_filter/n554 ), .Q(n1149) );
  BUF2 U1097 ( .A(\u_outFIFO/n549 ), .Q(n809) );
  BUF2 U1098 ( .A(\u_outFIFO/n547 ), .Q(n806) );
  BUF2 U1099 ( .A(\u_outFIFO/n480 ), .Q(n799) );
  BUF2 U1100 ( .A(\u_outFIFO/n478 ), .Q(n796) );
  BUF2 U1101 ( .A(\u_outFIFO/n476 ), .Q(n793) );
  BUF2 U1102 ( .A(\u_outFIFO/n411 ), .Q(n788) );
  BUF2 U1103 ( .A(\u_outFIFO/n409 ), .Q(n785) );
  BUF2 U1104 ( .A(\u_outFIFO/n407 ), .Q(n782) );
  BUF2 U1105 ( .A(\u_outFIFO/n549 ), .Q(n811) );
  BUF2 U1106 ( .A(\u_outFIFO/n547 ), .Q(n808) );
  BUF2 U1107 ( .A(\u_outFIFO/n549 ), .Q(n810) );
  BUF2 U1108 ( .A(\u_outFIFO/n547 ), .Q(n807) );
  BUF2 U1109 ( .A(\u_outFIFO/n480 ), .Q(n801) );
  BUF2 U1110 ( .A(\u_outFIFO/n478 ), .Q(n798) );
  BUF2 U1111 ( .A(\u_outFIFO/n476 ), .Q(n795) );
  BUF2 U1112 ( .A(\u_outFIFO/n480 ), .Q(n800) );
  BUF2 U1113 ( .A(\u_outFIFO/n478 ), .Q(n797) );
  BUF2 U1114 ( .A(\u_outFIFO/n476 ), .Q(n794) );
  BUF2 U1115 ( .A(\u_outFIFO/n411 ), .Q(n790) );
  BUF2 U1116 ( .A(\u_outFIFO/n409 ), .Q(n787) );
  BUF2 U1117 ( .A(\u_outFIFO/n407 ), .Q(n784) );
  BUF2 U1118 ( .A(\u_outFIFO/n411 ), .Q(n789) );
  BUF2 U1119 ( .A(\u_outFIFO/n409 ), .Q(n786) );
  BUF2 U1120 ( .A(\u_outFIFO/n407 ), .Q(n783) );
  INV3 U1121 ( .A(\u_decoder/iq_demod/dp_cluster_0/mult_151/SUMB[3][3] ), .Q(
        n693) );
  INV3 U1122 ( .A(\u_decoder/iq_demod/dp_cluster_1/mult_150/SUMB[3][3] ), .Q(
        n717) );
  INV3 U1123 ( .A(\u_decoder/iq_demod/dp_cluster_1/mult_149/CARRYB[3][3] ), 
        .Q(n2396) );
  INV3 U1124 ( .A(\u_decoder/iq_demod/dp_cluster_0/mult_148/CARRYB[3][3] ), 
        .Q(n2397) );
  NOR31 U1125 ( .A(\u_inFIFO/n551 ), .B(n2146), .C(\u_inFIFO/n549 ), .Q(
        \u_inFIFO/n533 ) );
  NAND22 U1126 ( .A(n1217), .B(\u_outFIFO/n1113 ), .Q(\u_outFIFO/n1114 ) );
  NOR21 U1127 ( .A(\u_outFIFO/n1127 ), .B(\u_outFIFO/n1120 ), .Q(
        \u_outFIFO/n1119 ) );
  INV3 U1128 ( .A(\u_inFIFO/n549 ), .Q(n1828) );
  NAND22 U1129 ( .A(n1219), .B(\u_cdr/n44 ), .Q(\u_cdr/n47 ) );
  NAND22 U1130 ( .A(n2217), .B(n1212), .Q(\u_outFIFO/n1127 ) );
  BUF2 U1131 ( .A(\u_decoder/fir_filter/n721 ), .Q(n1168) );
  BUF2 U1132 ( .A(\u_decoder/fir_filter/n721 ), .Q(n1170) );
  BUF2 U1133 ( .A(\u_decoder/fir_filter/n721 ), .Q(n1171) );
  BUF2 U1134 ( .A(\u_decoder/fir_filter/n721 ), .Q(n1169) );
  NAND22 U1135 ( .A(n1219), .B(n2098), .Q(\u_cdr/n24 ) );
  INV3 U1136 ( .A(\u_cdr/n39 ), .Q(n2098) );
  NOR31 U1137 ( .A(\u_coder/j [0]), .B(\u_coder/j [3]), .C(n2184), .Q(
        \u_coder/n206 ) );
  BUF2 U1138 ( .A(\u_decoder/fir_filter/n721 ), .Q(n1172) );
  NAND22 U1139 ( .A(\u_outFIFO/n1117 ), .B(n1216), .Q(\u_outFIFO/n1153 ) );
  NAND22 U1140 ( .A(n2176), .B(\u_coder/j [3]), .Q(\u_coder/n241 ) );
  BUF2 U1141 ( .A(\u_outFIFO/n326 ), .Q(n840) );
  BUF2 U1142 ( .A(\u_outFIFO/n326 ), .Q(n839) );
  BUF2 U1143 ( .A(\u_outFIFO/n376 ), .Q(n871) );
  BUF2 U1144 ( .A(\u_outFIFO/n376 ), .Q(n870) );
  BUF2 U1145 ( .A(\u_outFIFO/n356 ), .Q(n859) );
  BUF2 U1146 ( .A(\u_outFIFO/n356 ), .Q(n858) );
  BUF2 U1147 ( .A(\u_outFIFO/n361 ), .Q(n862) );
  BUF2 U1148 ( .A(\u_outFIFO/n361 ), .Q(n861) );
  BUF2 U1149 ( .A(\u_outFIFO/n341 ), .Q(n850) );
  BUF2 U1150 ( .A(\u_outFIFO/n341 ), .Q(n849) );
  BUF2 U1151 ( .A(\u_outFIFO/n371 ), .Q(n868) );
  BUF2 U1152 ( .A(\u_outFIFO/n371 ), .Q(n867) );
  BUF2 U1153 ( .A(\u_outFIFO/n366 ), .Q(n865) );
  BUF2 U1154 ( .A(\u_outFIFO/n366 ), .Q(n864) );
  BUF2 U1155 ( .A(\u_outFIFO/n351 ), .Q(n856) );
  BUF2 U1156 ( .A(\u_outFIFO/n351 ), .Q(n855) );
  BUF2 U1157 ( .A(\u_outFIFO/n346 ), .Q(n853) );
  BUF2 U1158 ( .A(\u_outFIFO/n346 ), .Q(n852) );
  BUF2 U1159 ( .A(\u_outFIFO/n326 ), .Q(n838) );
  BUF2 U1160 ( .A(\u_outFIFO/n376 ), .Q(n869) );
  BUF2 U1161 ( .A(\u_outFIFO/n356 ), .Q(n857) );
  BUF2 U1162 ( .A(\u_outFIFO/n361 ), .Q(n860) );
  BUF2 U1163 ( .A(\u_outFIFO/n341 ), .Q(n848) );
  BUF2 U1164 ( .A(\u_outFIFO/n371 ), .Q(n866) );
  BUF2 U1165 ( .A(\u_outFIFO/n366 ), .Q(n863) );
  BUF2 U1166 ( .A(\u_outFIFO/n351 ), .Q(n854) );
  BUF2 U1167 ( .A(\u_outFIFO/n346 ), .Q(n851) );
  NOR21 U1168 ( .A(\u_coder/n218 ), .B(n2097), .Q(\u_coder/n228 ) );
  NAND22 U1169 ( .A(n2175), .B(n2185), .Q(\u_coder/n224 ) );
  INV3 U1170 ( .A(\u_coder/n241 ), .Q(n2175) );
  BUF2 U1171 ( .A(\u_outFIFO/n612 ), .Q(n812) );
  BUF2 U1172 ( .A(\u_outFIFO/n612 ), .Q(n813) );
  BUF2 U1173 ( .A(\u_outFIFO/n975 ), .Q(n880) );
  BUF2 U1174 ( .A(\u_outFIFO/n975 ), .Q(n881) );
  BUF2 U1175 ( .A(\u_outFIFO/n474 ), .Q(n791) );
  BUF2 U1176 ( .A(\u_outFIFO/n474 ), .Q(n792) );
  BUF2 U1177 ( .A(\u_outFIFO/n405 ), .Q(n780) );
  BUF2 U1178 ( .A(\u_outFIFO/n405 ), .Q(n781) );
  BUF2 U1179 ( .A(\u_outFIFO/n972 ), .Q(n878) );
  BUF2 U1180 ( .A(\u_outFIFO/n972 ), .Q(n879) );
  BUF2 U1181 ( .A(\u_outFIFO/n839 ), .Q(n825) );
  BUF2 U1182 ( .A(\u_outFIFO/n839 ), .Q(n826) );
  BUF2 U1183 ( .A(\u_outFIFO/n706 ), .Q(n814) );
  BUF2 U1184 ( .A(\u_outFIFO/n706 ), .Q(n815) );
  BUF2 U1185 ( .A(\u_outFIFO/n543 ), .Q(n802) );
  BUF2 U1186 ( .A(\u_outFIFO/n543 ), .Q(n803) );
  BUF2 U1187 ( .A(n843), .Q(n844) );
  BUF2 U1188 ( .A(n843), .Q(n845) );
  BUF2 U1189 ( .A(\u_outFIFO/n336 ), .Q(n846) );
  BUF2 U1190 ( .A(\u_outFIFO/n336 ), .Q(n847) );
  INV3 U1191 ( .A(n888), .Q(n889) );
  INV3 U1192 ( .A(n876), .Q(n877) );
  INV3 U1193 ( .A(n874), .Q(n875) );
  INV3 U1194 ( .A(n841), .Q(n842) );
  INV3 U1195 ( .A(n872), .Q(n873) );
  INV3 U1196 ( .A(\u_decoder/fir_filter/dp_cluster_0/r164/CARRYB[7][3] ), .Q(
        n2305) );
  INV3 U1197 ( .A(\u_decoder/fir_filter/dp_cluster_0/r177/CARRYB[7][3] ), .Q(
        n2376) );
  INV3 U1198 ( .A(n836), .Q(n837) );
  INV3 U1199 ( .A(\u_coder/n235 ), .Q(n2173) );
  BUF2 U1200 ( .A(\u_outFIFO/n842 ), .Q(n827) );
  BUF2 U1201 ( .A(\u_outFIFO/n709 ), .Q(n816) );
  BUF2 U1202 ( .A(\u_outFIFO/n978 ), .Q(n882) );
  BUF2 U1203 ( .A(\u_outFIFO/n845 ), .Q(n830) );
  BUF2 U1204 ( .A(\u_outFIFO/n712 ), .Q(n819) );
  BUF2 U1205 ( .A(\u_outFIFO/n981 ), .Q(n885) );
  BUF2 U1206 ( .A(\u_outFIFO/n848 ), .Q(n833) );
  BUF2 U1207 ( .A(\u_outFIFO/n715 ), .Q(n822) );
  BUF2 U1208 ( .A(\u_outFIFO/n842 ), .Q(n829) );
  BUF2 U1209 ( .A(\u_outFIFO/n842 ), .Q(n828) );
  BUF2 U1210 ( .A(\u_outFIFO/n709 ), .Q(n818) );
  BUF2 U1211 ( .A(\u_outFIFO/n709 ), .Q(n817) );
  BUF2 U1212 ( .A(\u_outFIFO/n978 ), .Q(n884) );
  BUF2 U1213 ( .A(\u_outFIFO/n978 ), .Q(n883) );
  BUF2 U1214 ( .A(\u_outFIFO/n845 ), .Q(n832) );
  BUF2 U1215 ( .A(\u_outFIFO/n845 ), .Q(n831) );
  BUF2 U1216 ( .A(\u_outFIFO/n712 ), .Q(n821) );
  BUF2 U1217 ( .A(\u_outFIFO/n712 ), .Q(n820) );
  BUF2 U1218 ( .A(\u_outFIFO/n981 ), .Q(n887) );
  BUF2 U1219 ( .A(\u_outFIFO/n981 ), .Q(n886) );
  BUF2 U1220 ( .A(\u_outFIFO/n848 ), .Q(n835) );
  BUF2 U1221 ( .A(\u_outFIFO/n848 ), .Q(n834) );
  BUF2 U1222 ( .A(\u_outFIFO/n715 ), .Q(n824) );
  BUF2 U1223 ( .A(\u_outFIFO/n715 ), .Q(n823) );
  BUF2 U1224 ( .A(n1911), .Q(n980) );
  BUF2 U1225 ( .A(n1911), .Q(n979) );
  BUF2 U1226 ( .A(n1911), .Q(n978) );
  BUF2 U1227 ( .A(n1911), .Q(n977) );
  BUF2 U1228 ( .A(n1911), .Q(n976) );
  BUF2 U1229 ( .A(n1911), .Q(n975) );
  BUF2 U1230 ( .A(n1911), .Q(n974) );
  BUF2 U1231 ( .A(n1911), .Q(n973) );
  BUF2 U1232 ( .A(n1911), .Q(n972) );
  BUF2 U1233 ( .A(n1911), .Q(n971) );
  BUF2 U1234 ( .A(n1911), .Q(n970) );
  BUF2 U1235 ( .A(n1911), .Q(n969) );
  BUF2 U1236 ( .A(n1911), .Q(n968) );
  BUF2 U1237 ( .A(n1911), .Q(n967) );
  BUF2 U1238 ( .A(n1911), .Q(n966) );
  BUF2 U1239 ( .A(n1911), .Q(n965) );
  BUF2 U1240 ( .A(n1911), .Q(n964) );
  BUF2 U1241 ( .A(n1911), .Q(n963) );
  BUF2 U1242 ( .A(n1911), .Q(n962) );
  NAND22 U1243 ( .A(n1219), .B(n1796), .Q(\u_outFIFO/n1143 ) );
  INV3 U1244 ( .A(\u_cordic/mycordic/n548 ), .Q(n1907) );
  NAND22 U1245 ( .A(\u_cordic/mycordic/present_Q_table[4][7] ), .B(n1212), .Q(
        \u_cordic/mycordic/n548 ) );
  NAND22 U1246 ( .A(n1219), .B(\u_inFIFO/n531 ), .Q(\u_inFIFO/n217 ) );
  BUF2 U1247 ( .A(\u_cordic/mycordic/n363 ), .Q(n777) );
  XNR21 U1248 ( .A(n4), .B(\u_decoder/fir_filter/I_data_mult_0 [0]), .Q(n353)
         );
  XNR21 U1249 ( .A(n3), .B(\u_decoder/fir_filter/Q_data_mult_0 [0]), .Q(n354)
         );
  NAND22 U1250 ( .A(n1219), .B(\u_inFIFO/n217 ), .Q(\u_inFIFO/n216 ) );
  NAND22 U1251 ( .A(\u_decoder/iq_demod/cossin_dig/n41 ), .B(
        \u_decoder/iq_demod/cossin_dig/n40 ), .Q(
        \u_decoder/iq_demod/cossin_dig/n39 ) );
  NAND22 U1252 ( .A(n1218), .B(\u_decoder/iq_demod/cossin_dig/n42 ), .Q(
        \u_decoder/iq_demod/cossin_dig/n41 ) );
  BUF2 U1253 ( .A(\u_decoder/fir_filter/n721 ), .Q(n1174) );
  BUF2 U1254 ( .A(\u_decoder/fir_filter/n721 ), .Q(n1173) );
  BUF2 U1255 ( .A(\u_decoder/fir_filter/n721 ), .Q(n1175) );
  XNR21 U1256 ( .A(n8), .B(\u_decoder/fir_filter/I_data_mult_0 [0]), .Q(n355)
         );
  XNR21 U1257 ( .A(n7), .B(\u_decoder/fir_filter/Q_data_mult_0 [0]), .Q(n356)
         );
  XNR21 U1258 ( .A(\u_decoder/fir_filter/I_data_mult_0 [0]), .B(n12), .Q(n357)
         );
  XNR21 U1259 ( .A(\u_decoder/fir_filter/Q_data_mult_0 [0]), .B(n11), .Q(n358)
         );
  XNR21 U1260 ( .A(n4), .B(\u_decoder/fir_filter/I_data_mult_0 [0]), .Q(n359)
         );
  XNR21 U1261 ( .A(n3), .B(\u_decoder/fir_filter/Q_data_mult_0 [0]), .Q(n360)
         );
  INV3 U1262 ( .A(\u_decoder/iq_demod/n69 ), .Q(n1910) );
  NOR31 U1263 ( .A(n2208), .B(n1397), .C(n1237), .Q(\u_cdr/dec1/cnt_dec/n17 )
         );
  NOR31 U1264 ( .A(n1235), .B(n1397), .C(\u_cdr/dec1/cnt_dec/n24 ), .Q(
        \u_cdr/dec1/cnt_dec/n18 ) );
  NAND31 U1265 ( .A(n1219), .B(n2208), .C(n1392), .Q(n1393) );
  NOR31 U1266 ( .A(n1233), .B(n1396), .C(\u_cdr/div1/cnt_div/n41 ), .Q(
        \u_cdr/div1/cnt_div/n34 ) );
  NOR31 U1267 ( .A(n1234), .B(n1398), .C(n3064), .Q(n3057) );
  NOR31 U1268 ( .A(n2208), .B(n1396), .C(n1237), .Q(\u_cdr/div1/cnt_div/n35 )
         );
  INV3 U1269 ( .A(\u_cdr/div1/cnt_div/n41 ), .Q(n2208) );
  NOR31 U1270 ( .A(n2208), .B(n1398), .C(n1238), .Q(n3058) );
  NAND22 U1271 ( .A(n1283), .B(\u_cdr/div1/n7 ), .Q(n1388) );
  NAND31 U1272 ( .A(n1391), .B(n1392), .C(n1217), .Q(n1390) );
  INV3 U1273 ( .A(n3067), .Q(n1836) );
  NAND22 U1274 ( .A(\u_cdr/phd1/cnt_phd/N42 ), .B(n1217), .Q(n3067) );
  NOR40 U1275 ( .A(n3051), .B(n3050), .C(n2677), .D(\u_cdr/phd1/cnt_phd/N41 ), 
        .Q(\u_cdr/phd1/cnt_phd/N42 ) );
  NAND22 U1276 ( .A(n2679), .B(n3049), .Q(n3050) );
  OAI2111 U1277 ( .A(\u_cdr/div1/n9 ), .B(n59), .C(n1287), .D(n1313), .Q(n1349) );
  NOR21 U1278 ( .A(n1232), .B(n2675), .Q(\u_cdr/div1/cnt_div/N88 ) );
  AOI211 U1279 ( .A(n1265), .B(\u_cdr/w_sE ), .C(n1271), .Q(n1252) );
  NAND22 U1280 ( .A(n1218), .B(\u_cdr/phd1/n21 ), .Q(\u_cdr/phd1/n17 ) );
  INV3 U1281 ( .A(\u_cdr/phd1/n21 ), .Q(n1850) );
  AOI221 U1282 ( .A(\u_cordic/my_rotation/delta [7]), .B(n2674), .C(
        \u_cordic/my_rotation/N32 ), .D(n768), .Q(\u_cordic/my_rotation/n47 )
         );
  XOR21 U1283 ( .A(\u_cordic/my_rotation/delta [7]), .B(
        \u_cordic/my_rotation/add_38/carry [7]), .Q(\u_cordic/my_rotation/N32 ) );
  AOI221 U1284 ( .A(\u_cordic/my_rotation/delta [6]), .B(n2674), .C(
        \u_cordic/my_rotation/N31 ), .D(n768), .Q(\u_cordic/my_rotation/n48 )
         );
  XNR21 U1285 ( .A(\u_cordic/my_rotation/delta [6]), .B(
        \u_cordic/my_rotation/add_38/carry [6]), .Q(\u_cordic/my_rotation/N31 ) );
  NOR40 U1286 ( .A(n2669), .B(n2660), .C(n2668), .D(n2667), .Q(
        \u_cordic/my_rotation/n56 ) );
  INV3 U1287 ( .A(\u_cordic/my_rotation/n69 ), .Q(n2669) );
  AOI221 U1288 ( .A(\u_cordic/my_rotation/delta [1]), .B(n2674), .C(
        \u_cordic/my_rotation/delta [1]), .D(n767), .Q(
        \u_cordic/my_rotation/n69 ) );
  INV3 U1289 ( .A(\u_cordic/my_rotation/n64 ), .Q(n2665) );
  AOI221 U1290 ( .A(\u_cordic/my_rotation/delta [4]), .B(n2674), .C(
        \u_cordic/my_rotation/N29 ), .D(n768), .Q(\u_cordic/my_rotation/n64 )
         );
  XOR21 U1291 ( .A(\u_cordic/my_rotation/delta [4]), .B(
        \u_cordic/my_rotation/delta [3]), .Q(\u_cordic/my_rotation/N29 ) );
  INV3 U1292 ( .A(\u_cordic/my_rotation/n72 ), .Q(n2672) );
  AOI221 U1293 ( .A(\u_cordic/my_rotation/delta [11]), .B(n2674), .C(
        \u_cordic/my_rotation/N36 ), .D(n767), .Q(\u_cordic/my_rotation/n72 )
         );
  XOR21 U1294 ( .A(\u_cordic/my_rotation/delta [11]), .B(
        \u_cordic/my_rotation/add_38/carry [11]), .Q(
        \u_cordic/my_rotation/N36 ) );
  INV3 U1295 ( .A(\u_cordic/my_rotation/n71 ), .Q(n2671) );
  AOI221 U1296 ( .A(\u_cordic/my_rotation/delta [10]), .B(n2674), .C(
        \u_cordic/my_rotation/N35 ), .D(n767), .Q(\u_cordic/my_rotation/n71 )
         );
  XOR21 U1297 ( .A(\u_cordic/my_rotation/delta [10]), .B(
        \u_cordic/my_rotation/add_38/carry [10]), .Q(
        \u_cordic/my_rotation/N35 ) );
  INV3 U1298 ( .A(\u_cordic/my_rotation/n60 ), .Q(n2661) );
  AOI221 U1299 ( .A(\u_cordic/my_rotation/delta [9]), .B(n2674), .C(
        \u_cordic/my_rotation/N34 ), .D(n768), .Q(\u_cordic/my_rotation/n60 )
         );
  XOR21 U1300 ( .A(\u_cordic/my_rotation/delta [9]), .B(
        \u_cordic/my_rotation/add_38/carry [9]), .Q(\u_cordic/my_rotation/N34 ) );
  INV3 U1301 ( .A(\u_cordic/my_rotation/n61 ), .Q(n2662) );
  AOI221 U1302 ( .A(\u_cordic/my_rotation/delta [8]), .B(n2674), .C(
        \u_cordic/my_rotation/N33 ), .D(n768), .Q(\u_cordic/my_rotation/n61 )
         );
  XNR21 U1303 ( .A(\u_cordic/my_rotation/delta [8]), .B(
        \u_cordic/my_rotation/add_38/carry [8]), .Q(\u_cordic/my_rotation/N33 ) );
  INV3 U1304 ( .A(\u_cordic/my_rotation/n67 ), .Q(n2668) );
  AOI221 U1305 ( .A(\u_cordic/my_rotation/delta [14]), .B(n2674), .C(
        \u_cordic/my_rotation/N39 ), .D(n767), .Q(\u_cordic/my_rotation/n67 )
         );
  XOR21 U1306 ( .A(\u_cordic/my_rotation/delta [14]), .B(
        \u_cordic/my_rotation/add_38/carry [14]), .Q(
        \u_cordic/my_rotation/N39 ) );
  INV3 U1307 ( .A(\u_cordic/my_rotation/n66 ), .Q(n2667) );
  AOI221 U1308 ( .A(\u_cordic/my_rotation/delta [13]), .B(n2674), .C(
        \u_cordic/my_rotation/N38 ), .D(n768), .Q(\u_cordic/my_rotation/n66 )
         );
  XOR21 U1309 ( .A(\u_cordic/my_rotation/delta [13]), .B(
        \u_cordic/my_rotation/add_38/carry [13]), .Q(
        \u_cordic/my_rotation/N38 ) );
  BUF2 U1310 ( .A(\u_cordic/my_rotation/N23 ), .Q(n767) );
  BUF2 U1311 ( .A(\u_cordic/my_rotation/N23 ), .Q(n768) );
  INV3 U1312 ( .A(\u_cordic/my_rotation/n73 ), .Q(n2673) );
  AOI221 U1313 ( .A(\u_cordic/my_rotation/delta [12]), .B(n2674), .C(
        \u_cordic/my_rotation/N37 ), .D(n767), .Q(\u_cordic/my_rotation/n73 )
         );
  XOR21 U1314 ( .A(\u_cordic/my_rotation/delta [12]), .B(
        \u_cordic/my_rotation/add_38/carry [12]), .Q(
        \u_cordic/my_rotation/N37 ) );
  INV3 U1315 ( .A(\u_cordic/my_rotation/n63 ), .Q(n2664) );
  AOI221 U1316 ( .A(\u_cordic/my_rotation/delta [3]), .B(n2674), .C(n480), .D(
        n768), .Q(\u_cordic/my_rotation/n63 ) );
  INV3 U1317 ( .A(\u_cordic/my_rotation/n65 ), .Q(n2666) );
  AOI221 U1318 ( .A(\u_cordic/my_rotation/delta [5]), .B(n2674), .C(
        \u_cordic/my_rotation/N30 ), .D(n768), .Q(\u_cordic/my_rotation/n65 )
         );
  XNR21 U1319 ( .A(\u_cordic/my_rotation/delta [5]), .B(
        \u_cordic/my_rotation/add_38/carry [5]), .Q(\u_cordic/my_rotation/N30 ) );
  INV3 U1320 ( .A(\u_cordic/my_rotation/n62 ), .Q(n2663) );
  AOI221 U1321 ( .A(\u_cordic/my_rotation/delta [2]), .B(n2674), .C(
        \u_cordic/my_rotation/delta [2]), .D(n768), .Q(
        \u_cordic/my_rotation/n62 ) );
  INV3 U1322 ( .A(\u_cordic/my_rotation/delta [14]), .Q(n493) );
  INV3 U1323 ( .A(\u_cordic/my_rotation/n53 ), .Q(n1855) );
  NAND31 U1324 ( .A(n1219), .B(\u_cordic/my_rotation/n54 ), .C(n2659), .Q(
        \u_cordic/my_rotation/n53 ) );
  NAND41 U1325 ( .A(\u_cordic/my_rotation/n55 ), .B(\u_cordic/my_rotation/n56 ), .C(\u_cordic/my_rotation/n57 ), .D(\u_cordic/my_rotation/n58 ), .Q(
        \u_cordic/my_rotation/n54 ) );
  INV3 U1326 ( .A(n3042), .Q(n2659) );
  NOR21 U1327 ( .A(n396), .B(n482), .Q(\u_cordic/my_rotation/add_38/carry [8])
         );
  INV3 U1328 ( .A(\u_cordic/my_rotation/delta [7]), .Q(n482) );
  NOR21 U1329 ( .A(n484), .B(n485), .Q(\u_cordic/my_rotation/add_38/carry [11]) );
  INV3 U1330 ( .A(\u_cordic/my_rotation/add_38/carry [10]), .Q(n484) );
  INV3 U1331 ( .A(\u_cordic/my_rotation/delta [10]), .Q(n485) );
  NOR21 U1332 ( .A(n488), .B(n489), .Q(\u_cordic/my_rotation/add_38/carry [13]) );
  INV3 U1333 ( .A(\u_cordic/my_rotation/add_38/carry [12]), .Q(n488) );
  INV3 U1334 ( .A(\u_cordic/my_rotation/delta [12]), .Q(n489) );
  INV3 U1335 ( .A(n396), .Q(\u_cordic/my_rotation/add_38/carry [7]) );
  NOR21 U1336 ( .A(\u_cordic/my_rotation/add_38/carry [6]), .B(
        \u_cordic/my_rotation/delta [6]), .Q(n396) );
  INV3 U1337 ( .A(n397), .Q(\u_cordic/my_rotation/add_38/carry [9]) );
  NOR21 U1338 ( .A(\u_cordic/my_rotation/add_38/carry [8]), .B(
        \u_cordic/my_rotation/delta [8]), .Q(n397) );
  NOR21 U1339 ( .A(n397), .B(n483), .Q(\u_cordic/my_rotation/add_38/carry [10]) );
  INV3 U1340 ( .A(\u_cordic/my_rotation/delta [9]), .Q(n483) );
  NOR21 U1341 ( .A(n486), .B(n487), .Q(\u_cordic/my_rotation/add_38/carry [12]) );
  INV3 U1342 ( .A(\u_cordic/my_rotation/add_38/carry [11]), .Q(n486) );
  INV3 U1343 ( .A(\u_cordic/my_rotation/delta [11]), .Q(n487) );
  NOR21 U1344 ( .A(n490), .B(n491), .Q(\u_cordic/my_rotation/add_38/carry [14]) );
  INV3 U1345 ( .A(\u_cordic/my_rotation/add_38/carry [13]), .Q(n490) );
  INV3 U1346 ( .A(\u_cordic/my_rotation/delta [13]), .Q(n491) );
  NOR21 U1347 ( .A(\u_coder/n315 ), .B(n2188), .Q(\u_coder/N520 ) );
  INV3 U1348 ( .A(\u_coder/N475 ), .Q(n2188) );
  NOR21 U1349 ( .A(n895), .B(n2187), .Q(\u_coder/N521 ) );
  INV3 U1350 ( .A(\u_coder/N476 ), .Q(n2187) );
  XOR21 U1351 ( .A(n1192), .B(
        \u_decoder/fir_filter/dp_cluster_0/r166/SUMB[6][1] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r166/SUMB[7][0] ) );
  XOR21 U1352 ( .A(n1194), .B(
        \u_decoder/fir_filter/dp_cluster_0/r179/SUMB[6][1] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r179/SUMB[7][0] ) );
  XOR21 U1353 ( .A(n1193), .B(
        \u_decoder/fir_filter/dp_cluster_0/r165/SUMB[7][0] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r165/A1[5] ) );
  XOR21 U1354 ( .A(n1195), .B(
        \u_decoder/fir_filter/dp_cluster_0/r178/SUMB[7][0] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r178/A1[5] ) );
  XOR21 U1355 ( .A(n1192), .B(
        \u_decoder/fir_filter/dp_cluster_0/r166/SUMB[6][3] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r166/SUMB[7][2] ) );
  XOR21 U1356 ( .A(n1194), .B(
        \u_decoder/fir_filter/dp_cluster_0/r179/SUMB[6][3] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r179/SUMB[7][2] ) );
  XOR21 U1357 ( .A(n1192), .B(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/SUMB[6][5] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/SUMB[7][4] ) );
  XOR21 U1358 ( .A(n1194), .B(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/SUMB[6][5] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/SUMB[7][4] ) );
  XOR21 U1359 ( .A(n1192), .B(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/SUMB[5][3] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/SUMB[7][1] ) );
  XOR21 U1360 ( .A(n1194), .B(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/SUMB[5][3] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/SUMB[7][1] ) );
  XOR21 U1361 ( .A(n1192), .B(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/SUMB[6][3] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/SUMB[7][2] ) );
  XOR21 U1362 ( .A(n1194), .B(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/SUMB[6][3] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/SUMB[7][2] ) );
  XOR21 U1363 ( .A(n1193), .B(
        \u_decoder/fir_filter/dp_cluster_0/r165/SUMB[5][3] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r165/SUMB[7][1] ) );
  XOR21 U1364 ( .A(n1195), .B(
        \u_decoder/fir_filter/dp_cluster_0/r178/SUMB[5][3] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r178/SUMB[7][1] ) );
  XOR21 U1365 ( .A(n1193), .B(
        \u_decoder/fir_filter/dp_cluster_0/r165/SUMB[6][3] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r165/SUMB[7][2] ) );
  XOR21 U1366 ( .A(n1195), .B(
        \u_decoder/fir_filter/dp_cluster_0/r178/SUMB[6][3] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r178/SUMB[7][2] ) );
  XOR21 U1367 ( .A(n1193), .B(
        \u_decoder/fir_filter/dp_cluster_0/r164/SUMB[6][2] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r164/SUMB[7][1] ) );
  XOR21 U1368 ( .A(n1195), .B(
        \u_decoder/fir_filter/dp_cluster_0/r177/SUMB[6][2] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r177/SUMB[7][1] ) );
  NOR21 U1369 ( .A(n621), .B(n194), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r164/A2[6] ) );
  INV3 U1370 ( .A(\u_decoder/fir_filter/dp_cluster_0/r164/SUMB[7][0] ), .Q(
        n621) );
  NOR21 U1371 ( .A(n682), .B(n195), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r177/A2[6] ) );
  INV3 U1372 ( .A(\u_decoder/fir_filter/dp_cluster_0/r177/SUMB[7][0] ), .Q(
        n682) );
  NOR21 U1373 ( .A(n599), .B(n194), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r166/A2[6] ) );
  INV3 U1374 ( .A(\u_decoder/fir_filter/dp_cluster_0/r166/SUMB[7][0] ), .Q(
        n599) );
  NOR21 U1375 ( .A(n660), .B(n195), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r179/A2[6] ) );
  INV3 U1376 ( .A(\u_decoder/fir_filter/dp_cluster_0/r179/SUMB[7][0] ), .Q(
        n660) );
  NOR21 U1377 ( .A(n609), .B(n194), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r165/A2[6] ) );
  INV3 U1378 ( .A(\u_decoder/fir_filter/dp_cluster_0/r165/SUMB[7][0] ), .Q(
        n609) );
  NOR21 U1379 ( .A(n670), .B(n195), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r178/A2[6] ) );
  INV3 U1380 ( .A(\u_decoder/fir_filter/dp_cluster_0/r178/SUMB[7][0] ), .Q(
        n670) );
  INV3 U1381 ( .A(n2930), .Q(n2276) );
  AOI2111 U1382 ( .A(n2931), .B(
        \u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[7][5] ), .C(n2277), .D(
        n2932), .Q(n2930) );
  XNR21 U1383 ( .A(n1193), .B(n2916), .Q(n361) );
  INV3 U1384 ( .A(n2844), .Q(n2347) );
  AOI2111 U1385 ( .A(n2845), .B(
        \u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[7][5] ), .C(n2348), .D(
        n2846), .Q(n2844) );
  XNR21 U1386 ( .A(n1195), .B(n2830), .Q(n362) );
  NOR21 U1387 ( .A(n480), .B(n481), .Q(\u_cordic/my_rotation/add_38/carry [5])
         );
  INV3 U1388 ( .A(\u_cordic/my_rotation/delta [3]), .Q(n480) );
  INV3 U1389 ( .A(\u_cordic/my_rotation/delta [4]), .Q(n481) );
  NOR21 U1390 ( .A(n194), .B(n752), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r166/CARRYB[7][0] ) );
  INV3 U1391 ( .A(\u_decoder/fir_filter/dp_cluster_0/r166/SUMB[6][1] ), .Q(
        n752) );
  NOR21 U1392 ( .A(n195), .B(n743), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r179/CARRYB[7][0] ) );
  INV3 U1393 ( .A(\u_decoder/fir_filter/dp_cluster_0/r179/SUMB[6][1] ), .Q(
        n743) );
  NOR21 U1394 ( .A(n194), .B(n747), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r164/CARRYB[7][1] ) );
  INV3 U1395 ( .A(\u_decoder/fir_filter/dp_cluster_0/r164/SUMB[6][2] ), .Q(
        n747) );
  NOR21 U1396 ( .A(n195), .B(n738), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r177/CARRYB[7][1] ) );
  INV3 U1397 ( .A(\u_decoder/fir_filter/dp_cluster_0/r177/SUMB[6][2] ), .Q(
        n738) );
  NOR21 U1398 ( .A(n194), .B(n754), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r165/CARRYB[7][1] ) );
  INV3 U1399 ( .A(\u_decoder/fir_filter/dp_cluster_0/r165/SUMB[5][3] ), .Q(
        n754) );
  NOR21 U1400 ( .A(n195), .B(n745), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r178/CARRYB[7][1] ) );
  INV3 U1401 ( .A(\u_decoder/fir_filter/dp_cluster_0/r178/SUMB[5][3] ), .Q(
        n745) );
  NOR21 U1402 ( .A(n194), .B(n750), .Q(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[7][2] ) );
  INV3 U1403 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_276/SUMB[6][3] ), 
        .Q(n750) );
  NOR21 U1404 ( .A(n195), .B(n741), .Q(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[7][2] ) );
  INV3 U1405 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_308/SUMB[6][3] ), 
        .Q(n741) );
  NAND22 U1406 ( .A(\u_decoder/fir_filter/I_data_mult_2_15 ), .B(n1083), .Q(
        \u_decoder/fir_filter/n1050 ) );
  XNR21 U1407 ( .A(n1193), .B(n2915), .Q(
        \u_decoder/fir_filter/I_data_mult_2_15 ) );
  NAND22 U1408 ( .A(n2916), .B(n1193), .Q(n2915) );
  NAND22 U1409 ( .A(\u_decoder/fir_filter/Q_data_mult_2_15 ), .B(n1083), .Q(
        \u_decoder/fir_filter/n753 ) );
  XNR21 U1410 ( .A(n1195), .B(n2829), .Q(
        \u_decoder/fir_filter/Q_data_mult_2_15 ) );
  NAND22 U1411 ( .A(n2830), .B(n1195), .Q(n2829) );
  NOR21 U1412 ( .A(n895), .B(n2189), .Q(\u_coder/N519 ) );
  INV3 U1413 ( .A(\u_coder/N474 ), .Q(n2189) );
  INV3 U1414 ( .A(n395), .Q(\u_cordic/my_rotation/add_38/carry [6]) );
  NOR21 U1415 ( .A(\u_cordic/my_rotation/add_38/carry [5]), .B(
        \u_cordic/my_rotation/delta [5]), .Q(n395) );
  NAND22 U1416 ( .A(\u_decoder/fir_filter/dp_cluster_0/r167/SUMB[7][0] ), .B(
        n1192), .Q(n363) );
  NAND22 U1417 ( .A(\u_decoder/fir_filter/dp_cluster_0/r180/SUMB[7][0] ), .B(
        n1194), .Q(n364) );
  INV3 U1418 ( .A(n3002), .Q(n2528) );
  INV3 U1419 ( .A(n2983), .Q(n2408) );
  INV3 U1420 ( .A(n2993), .Q(n2536) );
  INV3 U1421 ( .A(n2974), .Q(n2416) );
  NOR21 U1422 ( .A(\u_coder/n315 ), .B(n2190), .Q(\u_coder/N518 ) );
  INV3 U1423 ( .A(\u_coder/N473 ), .Q(n2190) );
  NOR21 U1424 ( .A(n895), .B(n2191), .Q(\u_coder/N517 ) );
  INV3 U1425 ( .A(\u_coder/N472 ), .Q(n2191) );
  XOR21 U1426 ( .A(\u_decoder/iq_demod/dp_cluster_0/mult_151/SUMB[3][1] ), .B(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/CARRYB[3][0] ), .Q(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/A1[2] ) );
  XOR21 U1427 ( .A(\u_decoder/iq_demod/dp_cluster_1/mult_150/SUMB[3][1] ), .B(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/CARRYB[3][0] ), .Q(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/A1[2] ) );
  XOR21 U1428 ( .A(\u_decoder/iq_demod/dp_cluster_1/mult_149/SUMB[3][1] ), .B(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/CARRYB[3][0] ), .Q(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/A1[2] ) );
  XOR21 U1429 ( .A(\u_decoder/iq_demod/dp_cluster_0/mult_148/SUMB[3][1] ), .B(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/CARRYB[3][0] ), .Q(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/A1[2] ) );
  XOR21 U1430 ( .A(\u_decoder/iq_demod/dp_cluster_0/mult_151/SUMB[3][2] ), .B(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/CARRYB[3][1] ), .Q(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/A1[3] ) );
  XOR21 U1431 ( .A(\u_decoder/iq_demod/dp_cluster_1/mult_150/SUMB[3][2] ), .B(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/CARRYB[3][1] ), .Q(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/A1[3] ) );
  XOR21 U1432 ( .A(\u_decoder/iq_demod/dp_cluster_1/mult_149/SUMB[3][2] ), .B(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/CARRYB[3][1] ), .Q(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/A1[3] ) );
  XOR21 U1433 ( .A(\u_decoder/iq_demod/dp_cluster_0/mult_148/SUMB[3][2] ), .B(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/CARRYB[3][1] ), .Q(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/A1[3] ) );
  XOR21 U1434 ( .A(n1192), .B(
        \u_decoder/fir_filter/dp_cluster_0/r167/SUMB[6][3] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r167/SUMB[7][2] ) );
  XOR21 U1435 ( .A(n1194), .B(
        \u_decoder/fir_filter/dp_cluster_0/r180/SUMB[6][3] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r180/SUMB[7][2] ) );
  XOR21 U1436 ( .A(n1193), .B(
        \u_decoder/fir_filter/dp_cluster_0/r164/SUMB[7][0] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r164/A1[5] ) );
  XOR21 U1437 ( .A(n1195), .B(
        \u_decoder/fir_filter/dp_cluster_0/r177/SUMB[7][0] ), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r177/A1[5] ) );
  NOR21 U1438 ( .A(n124), .B(n41), .Q(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/ab[2][1] ) );
  NOR21 U1439 ( .A(n720), .B(n721), .Q(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/CARRYB[1][1] ) );
  XOR21 U1440 ( .A(\u_decoder/iq_demod/dp_cluster_1/mult_150/ab[0][3] ), .B(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/ab[1][2] ), .Q(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/SUMB[1][2] ) );
  NOR21 U1441 ( .A(n125), .B(n44), .Q(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/ab[2][1] ) );
  NOR21 U1442 ( .A(n732), .B(n733), .Q(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/CARRYB[1][1] ) );
  XOR21 U1443 ( .A(\u_decoder/iq_demod/dp_cluster_1/mult_149/ab[0][3] ), .B(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/ab[1][2] ), .Q(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/SUMB[1][2] ) );
  NOR21 U1444 ( .A(n125), .B(n41), .Q(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/ab[2][1] ) );
  NOR21 U1445 ( .A(n708), .B(n709), .Q(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/CARRYB[1][1] ) );
  XOR21 U1446 ( .A(\u_decoder/iq_demod/dp_cluster_0/mult_148/ab[0][3] ), .B(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/ab[1][2] ), .Q(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/SUMB[1][2] ) );
  NOR21 U1447 ( .A(n124), .B(n42), .Q(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/ab[2][0] ) );
  NOR21 U1448 ( .A(n694), .B(n695), .Q(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/CARRYB[1][0] ) );
  XOR21 U1449 ( .A(\u_decoder/iq_demod/dp_cluster_0/mult_151/ab[0][2] ), .B(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/ab[1][1] ), .Q(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/SUMB[1][1] ) );
  NOR21 U1450 ( .A(n124), .B(n40), .Q(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/ab[2][0] ) );
  NOR21 U1451 ( .A(n718), .B(n719), .Q(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/CARRYB[1][0] ) );
  XOR21 U1452 ( .A(\u_decoder/iq_demod/dp_cluster_1/mult_150/ab[0][2] ), .B(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/ab[1][1] ), .Q(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/SUMB[1][1] ) );
  NOR21 U1453 ( .A(n125), .B(n42), .Q(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/ab[2][0] ) );
  NOR21 U1454 ( .A(n730), .B(n731), .Q(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/CARRYB[1][0] ) );
  XOR21 U1455 ( .A(\u_decoder/iq_demod/dp_cluster_1/mult_149/ab[0][2] ), .B(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/ab[1][1] ), .Q(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/SUMB[1][1] ) );
  NOR21 U1456 ( .A(n125), .B(n40), .Q(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/ab[2][0] ) );
  NOR21 U1457 ( .A(n706), .B(n707), .Q(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/CARRYB[1][0] ) );
  XOR21 U1458 ( .A(\u_decoder/iq_demod/dp_cluster_0/mult_148/ab[0][2] ), .B(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/ab[1][1] ), .Q(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/SUMB[1][1] ) );
  NOR21 U1459 ( .A(n42), .B(n120), .Q(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/ab[1][0] ) );
  NOR21 U1460 ( .A(n45), .B(n120), .Q(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/ab[1][2] ) );
  NOR21 U1461 ( .A(n44), .B(n120), .Q(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/ab[1][1] ) );
  NOR21 U1462 ( .A(n43), .B(n120), .Q(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/ab[1][2] ) );
  NOR21 U1463 ( .A(n41), .B(n120), .Q(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/ab[1][1] ) );
  NOR21 U1464 ( .A(n45), .B(n121), .Q(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/ab[1][2] ) );
  NOR21 U1465 ( .A(n44), .B(n121), .Q(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/ab[1][1] ) );
  NOR21 U1466 ( .A(n43), .B(n121), .Q(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/ab[1][2] ) );
  NOR21 U1467 ( .A(n41), .B(n121), .Q(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/ab[1][1] ) );
  NOR21 U1468 ( .A(n40), .B(n120), .Q(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/ab[1][0] ) );
  NOR21 U1469 ( .A(n42), .B(n121), .Q(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/ab[1][0] ) );
  NOR21 U1470 ( .A(n40), .B(n121), .Q(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/ab[1][0] ) );
  NOR21 U1471 ( .A(n44), .B(n123), .Q(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/ab[0][1] ) );
  NOR21 U1472 ( .A(n45), .B(n123), .Q(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/ab[0][2] ) );
  NOR21 U1473 ( .A(n43), .B(n123), .Q(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/ab[0][2] ) );
  NOR21 U1474 ( .A(n45), .B(n122), .Q(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/ab[0][2] ) );
  NOR21 U1475 ( .A(n43), .B(n122), .Q(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/ab[0][2] ) );
  NOR21 U1476 ( .A(n41), .B(n123), .Q(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/ab[0][1] ) );
  NOR21 U1477 ( .A(n44), .B(n122), .Q(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/ab[0][1] ) );
  NOR21 U1478 ( .A(n41), .B(n122), .Q(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/ab[0][1] ) );
  XNR21 U1479 ( .A(n2770), .B(n2771), .Q(
        \u_decoder/iq_demod/dp_cluster_1/mult_I_sin_out [5]) );
  XNR21 U1480 ( .A(n2777), .B(n2778), .Q(
        \u_decoder/iq_demod/dp_cluster_1/mult_Q_cos_out [5]) );
  NAND22 U1481 ( .A(\u_decoder/iq_demod/dp_cluster_1/mult_149/A2[2] ), .B(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/A1[2] ), .Q(n2770) );
  INV3 U1482 ( .A(\u_decoder/iq_demod/dp_cluster_0/mult_Q_sin_out [3]), .Q(
        n2387) );
  NOR21 U1483 ( .A(n194), .B(n748), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[7][2] ) );
  INV3 U1484 ( .A(\u_decoder/fir_filter/dp_cluster_0/r167/SUMB[6][3] ), .Q(
        n748) );
  NOR21 U1485 ( .A(n195), .B(n739), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[7][2] ) );
  INV3 U1486 ( .A(\u_decoder/fir_filter/dp_cluster_0/r180/SUMB[6][3] ), .Q(
        n739) );
  NOR21 U1487 ( .A(n194), .B(n755), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r165/CARRYB[7][2] ) );
  INV3 U1488 ( .A(\u_decoder/fir_filter/dp_cluster_0/r165/SUMB[6][3] ), .Q(
        n755) );
  NOR21 U1489 ( .A(n195), .B(n746), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r178/CARRYB[7][2] ) );
  INV3 U1490 ( .A(\u_decoder/fir_filter/dp_cluster_0/r178/SUMB[6][3] ), .Q(
        n746) );
  NOR21 U1491 ( .A(n194), .B(n751), .Q(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[7][4] ) );
  INV3 U1492 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_276/SUMB[6][5] ), 
        .Q(n751) );
  NOR21 U1493 ( .A(n194), .B(n753), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r166/CARRYB[7][2] ) );
  INV3 U1494 ( .A(\u_decoder/fir_filter/dp_cluster_0/r166/SUMB[6][3] ), .Q(
        n753) );
  NOR21 U1495 ( .A(n195), .B(n742), .Q(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[7][4] ) );
  INV3 U1496 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_308/SUMB[6][5] ), 
        .Q(n742) );
  NOR21 U1497 ( .A(n195), .B(n744), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r179/CARRYB[7][2] ) );
  INV3 U1498 ( .A(\u_decoder/fir_filter/dp_cluster_0/r179/SUMB[6][3] ), .Q(
        n744) );
  NOR21 U1499 ( .A(n194), .B(n749), .Q(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[7][1] ) );
  INV3 U1500 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_276/SUMB[5][3] ), 
        .Q(n749) );
  NOR21 U1501 ( .A(n195), .B(n740), .Q(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[7][1] ) );
  INV3 U1502 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_308/SUMB[5][3] ), 
        .Q(n740) );
  NOR21 U1503 ( .A(n124), .B(n44), .Q(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/ab[2][1] ) );
  NOR21 U1504 ( .A(n696), .B(n697), .Q(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/CARRYB[1][1] ) );
  XOR21 U1505 ( .A(\u_decoder/iq_demod/dp_cluster_0/mult_151/ab[0][3] ), .B(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/ab[1][2] ), .Q(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/SUMB[1][2] ) );
  NAND22 U1506 ( .A(\u_decoder/iq_demod/dp_cluster_0/mult_151/A2[2] ), .B(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/A1[2] ), .Q(n2791) );
  NAND22 U1507 ( .A(\u_decoder/iq_demod/dp_cluster_1/mult_150/A2[2] ), .B(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/A1[2] ), .Q(n2777) );
  NAND22 U1508 ( .A(\u_decoder/iq_demod/dp_cluster_0/mult_148/A2[2] ), .B(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/A1[2] ), .Q(n2784) );
  NOR21 U1509 ( .A(\u_coder/n315 ), .B(n2192), .Q(\u_coder/N516 ) );
  INV3 U1510 ( .A(\u_coder/N471 ), .Q(n2192) );
  INV3 U1511 ( .A(\u_decoder/iq_demod/dp_cluster_0/mult_151/A2[2] ), .Q(n2386)
         );
  INV3 U1512 ( .A(\u_decoder/iq_demod/dp_cluster_1/mult_150/A2[2] ), .Q(n2382)
         );
  INV3 U1513 ( .A(\u_decoder/iq_demod/dp_cluster_1/mult_149/A2[2] ), .Q(n2392)
         );
  INV3 U1514 ( .A(\u_decoder/iq_demod/dp_cluster_0/mult_148/A2[2] ), .Q(n2395)
         );
  NAND22 U1515 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_276/SUMB[7][0] ), 
        .B(n1192), .Q(n365) );
  NAND22 U1516 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_308/SUMB[7][0] ), 
        .B(n1194), .Q(n366) );
  NOR21 U1517 ( .A(n688), .B(n689), .Q(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/A2[3] ) );
  INV3 U1518 ( .A(\u_decoder/iq_demod/dp_cluster_0/mult_151/CARRYB[3][0] ), 
        .Q(n688) );
  INV3 U1519 ( .A(\u_decoder/iq_demod/dp_cluster_0/mult_151/SUMB[3][1] ), .Q(
        n689) );
  NOR21 U1520 ( .A(n712), .B(n713), .Q(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/A2[3] ) );
  INV3 U1521 ( .A(\u_decoder/iq_demod/dp_cluster_1/mult_150/CARRYB[3][0] ), 
        .Q(n712) );
  INV3 U1522 ( .A(\u_decoder/iq_demod/dp_cluster_1/mult_150/SUMB[3][1] ), .Q(
        n713) );
  NOR21 U1523 ( .A(n724), .B(n725), .Q(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/A2[3] ) );
  INV3 U1524 ( .A(\u_decoder/iq_demod/dp_cluster_1/mult_149/CARRYB[3][0] ), 
        .Q(n724) );
  INV3 U1525 ( .A(\u_decoder/iq_demod/dp_cluster_1/mult_149/SUMB[3][1] ), .Q(
        n725) );
  NOR21 U1526 ( .A(n700), .B(n701), .Q(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/A2[3] ) );
  INV3 U1527 ( .A(\u_decoder/iq_demod/dp_cluster_0/mult_148/CARRYB[3][0] ), 
        .Q(n700) );
  INV3 U1528 ( .A(\u_decoder/iq_demod/dp_cluster_0/mult_148/SUMB[3][1] ), .Q(
        n701) );
  INV3 U1529 ( .A(\u_decoder/iq_demod/dp_cluster_0/mult_151/ab[0][3] ), .Q(
        n698) );
  INV3 U1530 ( .A(\u_decoder/iq_demod/dp_cluster_1/mult_150/ab[0][3] ), .Q(
        n722) );
  INV3 U1531 ( .A(\u_decoder/iq_demod/dp_cluster_1/mult_149/ab[0][3] ), .Q(
        n734) );
  INV3 U1532 ( .A(\u_decoder/iq_demod/dp_cluster_0/mult_148/ab[0][3] ), .Q(
        n710) );
  NOR21 U1533 ( .A(n895), .B(n2193), .Q(\u_coder/N515 ) );
  INV3 U1534 ( .A(\u_coder/N470 ), .Q(n2193) );
  INV3 U1535 ( .A(\u_decoder/iq_demod/n57 ), .Q(n2378) );
  AOI221 U1536 ( .A(\u_decoder/iq_demod/add_Q_out [7]), .B(n779), .C(n1195), 
        .D(\u_decoder/iq_demod/state [1]), .Q(\u_decoder/iq_demod/n57 ) );
  INV3 U1537 ( .A(\u_decoder/iq_demod/n56 ), .Q(n2377) );
  AOI221 U1538 ( .A(\u_decoder/iq_demod/add_Q_out [6]), .B(n779), .C(n5), .D(
        \u_decoder/iq_demod/state [1]), .Q(\u_decoder/iq_demod/n56 ) );
  INV3 U1539 ( .A(\u_decoder/iq_demod/n49 ), .Q(n2307) );
  AOI221 U1540 ( .A(\u_decoder/iq_demod/add_I_out [7]), .B(n779), .C(n1193), 
        .D(\u_decoder/iq_demod/state [1]), .Q(\u_decoder/iq_demod/n49 ) );
  INV3 U1541 ( .A(\u_decoder/iq_demod/n48 ), .Q(n2306) );
  AOI221 U1542 ( .A(\u_decoder/iq_demod/add_I_out [6]), .B(n779), .C(n6), .D(
        \u_decoder/iq_demod/state [1]), .Q(\u_decoder/iq_demod/n48 ) );
  AOI2111 U1543 ( .A(\u_coder/n170 ), .B(\u_coder/n91 ), .C(n2161), .D(
        \u_coder/n254 ), .Q(\u_coder/n245 ) );
  NAND22 U1544 ( .A(\u_coder/n91 ), .B(n2105), .Q(\u_coder/n139 ) );
  XOR21 U1545 ( .A(\u_decoder/iq_demod/dp_cluster_0/mult_151/SUMB[3][3] ), .B(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/CARRYB[3][2] ), .Q(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/A1[4] ) );
  XOR21 U1546 ( .A(\u_decoder/iq_demod/dp_cluster_1/mult_150/SUMB[3][3] ), .B(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/CARRYB[3][2] ), .Q(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/A1[4] ) );
  XOR21 U1547 ( .A(\u_decoder/iq_demod/dp_cluster_1/mult_149/SUMB[3][3] ), .B(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/CARRYB[3][2] ), .Q(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/A1[4] ) );
  XOR21 U1548 ( .A(\u_decoder/iq_demod/dp_cluster_0/mult_148/SUMB[3][3] ), .B(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/CARRYB[3][2] ), .Q(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/A1[4] ) );
  NOR40 U1549 ( .A(n2144), .B(n2692), .C(\u_inFIFO/N135 ), .D(\u_inFIFO/N134 ), 
        .Q(\u_inFIFO/N375 ) );
  NAND22 U1550 ( .A(\u_inFIFO/N140 ), .B(n2148), .Q(n2692) );
  INV3 U1551 ( .A(n2691), .Q(n2144) );
  INV3 U1552 ( .A(\u_inFIFO/N133 ), .Q(n2148) );
  NAND22 U1553 ( .A(\u_coder/n94 ), .B(\u_coder/n213 ), .Q(\u_coder/n182 ) );
  NOR40 U1554 ( .A(n2222), .B(n2745), .C(\u_outFIFO/N145 ), .D(
        \u_outFIFO/N144 ), .Q(\u_outFIFO/N1269 ) );
  NAND22 U1555 ( .A(\u_outFIFO/N150 ), .B(n2228), .Q(n2745) );
  INV3 U1556 ( .A(n2744), .Q(n2222) );
  INV3 U1557 ( .A(\u_outFIFO/N143 ), .Q(n2228) );
  NOR21 U1558 ( .A(n23), .B(\u_decoder/iq_demod/I_if_buff[3] ), .Q(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/ab[3][3] ) );
  NOR21 U1559 ( .A(n23), .B(\u_decoder/iq_demod/Q_if_buff[3] ), .Q(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/ab[3][3] ) );
  NOR21 U1560 ( .A(n22), .B(\u_decoder/iq_demod/I_if_buff[3] ), .Q(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/ab[3][3] ) );
  NOR21 U1561 ( .A(n22), .B(\u_decoder/iq_demod/Q_if_buff[3] ), .Q(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/ab[3][3] ) );
  NAND31 U1562 ( .A(\u_coder/n166 ), .B(\u_coder/n167 ), .C(\u_coder/n168 ), 
        .Q(\u_coder/n135 ) );
  AOI211 U1563 ( .A(n2168), .B(\u_coder/n169 ), .C(n1241), .Q(\u_coder/n168 )
         );
  OAI311 U1564 ( .A(\u_coder/n170 ), .B(\u_coder/n137 ), .C(\u_coder/n149 ), 
        .D(\u_coder/n91 ), .Q(\u_coder/n166 ) );
  NOR40 U1565 ( .A(\u_outFIFO/N149 ), .B(\u_outFIFO/N148 ), .C(
        \u_outFIFO/N147 ), .D(\u_outFIFO/N146 ), .Q(n2744) );
  NOR40 U1566 ( .A(\u_inFIFO/N139 ), .B(\u_inFIFO/N138 ), .C(\u_inFIFO/N137 ), 
        .D(\u_inFIFO/N136 ), .Q(n2691) );
  AOI211 U1567 ( .A(\u_outFIFO/n1149 ), .B(n2223), .C(\u_outFIFO/n1151 ), .Q(
        \u_outFIFO/n1150 ) );
  INV3 U1568 ( .A(\u_outFIFO/N1270 ), .Q(n2223) );
  INV3 U1569 ( .A(\u_coder/n280 ), .Q(n1917) );
  AOI221 U1570 ( .A(\u_coder/N1014 ), .B(n2169), .C(\u_coder/n263 ), .D(n762), 
        .Q(\u_coder/n280 ) );
  XNR21 U1571 ( .A(n1192), .B(
        \u_decoder/fir_filter/dp_cluster_0/r166/SUMB[7][0] ), .Q(n367) );
  XNR21 U1572 ( .A(n1194), .B(
        \u_decoder/fir_filter/dp_cluster_0/r179/SUMB[7][0] ), .Q(n368) );
  NOR21 U1573 ( .A(n40), .B(n122), .Q(
        \u_decoder/iq_demod/dp_cluster_0/mult_I_cos_out [0]) );
  NOR21 U1574 ( .A(n40), .B(n123), .Q(
        \u_decoder/iq_demod/dp_cluster_1/mult_Q_cos_out [0]) );
  NOR21 U1575 ( .A(n42), .B(n122), .Q(
        \u_decoder/iq_demod/dp_cluster_1/mult_I_sin_out [0]) );
  BUF2 U1576 ( .A(n891), .Q(n893) );
  AOI211 U1577 ( .A(n2168), .B(n2157), .C(\u_coder/n255 ), .Q(n891) );
  BUF2 U1578 ( .A(n892), .Q(n894) );
  AOI211 U1579 ( .A(n2168), .B(n2157), .C(\u_coder/n255 ), .Q(n892) );
  AOI311 U1580 ( .A(\u_inFIFO/n564 ), .B(\u_inFIFO/n531 ), .C(\u_inFIFO/n569 ), 
        .D(n1241), .Q(\u_inFIFO/N47 ) );
  AOI311 U1581 ( .A(n2142), .B(\u_inFIFO/n557 ), .C(\u_inFIFO/sig_fsm_start_R ), .D(\u_inFIFO/n570 ), .Q(\u_inFIFO/n569 ) );
  NOR21 U1582 ( .A(n2143), .B(\u_inFIFO/n563 ), .Q(\u_inFIFO/n570 ) );
  AOI221 U1583 ( .A(\u_inFIFO/n561 ), .B(n2143), .C(\u_inFIFO/n560 ), .D(n2711), .Q(\u_inFIFO/n562 ) );
  NOR21 U1584 ( .A(\u_coder/n315 ), .B(n2194), .Q(\u_coder/N514 ) );
  INV3 U1585 ( .A(\u_coder/N469 ), .Q(n2194) );
  INV3 U1586 ( .A(\u_coder/n170 ), .Q(n2105) );
  INV3 U1587 ( .A(\u_decoder/iq_demod/dp_cluster_0/mult_Q_sin_out [0]), .Q(
        n2383) );
  NOR21 U1588 ( .A(n42), .B(n123), .Q(
        \u_decoder/iq_demod/dp_cluster_0/mult_Q_sin_out [0]) );
  NOR21 U1589 ( .A(n714), .B(n715), .Q(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/A2[4] ) );
  INV3 U1590 ( .A(\u_decoder/iq_demod/dp_cluster_1/mult_150/CARRYB[3][1] ), 
        .Q(n714) );
  INV3 U1591 ( .A(\u_decoder/iq_demod/dp_cluster_1/mult_150/SUMB[3][2] ), .Q(
        n715) );
  NOR21 U1592 ( .A(n702), .B(n703), .Q(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/A2[4] ) );
  INV3 U1593 ( .A(\u_decoder/iq_demod/dp_cluster_0/mult_148/CARRYB[3][1] ), 
        .Q(n702) );
  INV3 U1594 ( .A(\u_decoder/iq_demod/dp_cluster_0/mult_148/SUMB[3][2] ), .Q(
        n703) );
  AOI211 U1595 ( .A(n2185), .B(n2170), .C(\u_coder/n239 ), .Q(n890) );
  AOI211 U1596 ( .A(n2185), .B(n2170), .C(\u_coder/n239 ), .Q(\u_coder/n263 )
         );
  XNR21 U1597 ( .A(n1192), .B(
        \u_decoder/fir_filter/dp_cluster_0/r167/SUMB[7][0] ), .Q(n369) );
  XNR21 U1598 ( .A(n1194), .B(
        \u_decoder/fir_filter/dp_cluster_0/r180/SUMB[7][0] ), .Q(n370) );
  INV3 U1599 ( .A(\u_decoder/iq_demod/dp_cluster_0/mult_151/CARRYB[3][2] ), 
        .Q(n692) );
  INV3 U1600 ( .A(\u_decoder/iq_demod/dp_cluster_1/mult_150/CARRYB[3][2] ), 
        .Q(n716) );
  NOR21 U1601 ( .A(n726), .B(n727), .Q(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/A2[4] ) );
  INV3 U1602 ( .A(\u_decoder/iq_demod/dp_cluster_1/mult_149/CARRYB[3][1] ), 
        .Q(n726) );
  INV3 U1603 ( .A(\u_decoder/iq_demod/dp_cluster_1/mult_149/SUMB[3][2] ), .Q(
        n727) );
  NOR21 U1604 ( .A(n690), .B(n691), .Q(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/A2[4] ) );
  INV3 U1605 ( .A(\u_decoder/iq_demod/dp_cluster_0/mult_151/CARRYB[3][1] ), 
        .Q(n690) );
  INV3 U1606 ( .A(\u_decoder/iq_demod/dp_cluster_0/mult_151/SUMB[3][2] ), .Q(
        n691) );
  NOR21 U1607 ( .A(n728), .B(n729), .Q(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/A2[5] ) );
  INV3 U1608 ( .A(\u_decoder/iq_demod/dp_cluster_1/mult_149/SUMB[3][3] ), .Q(
        n729) );
  INV3 U1609 ( .A(\u_decoder/iq_demod/dp_cluster_1/mult_149/CARRYB[3][2] ), 
        .Q(n728) );
  NOR21 U1610 ( .A(n704), .B(n705), .Q(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/A2[5] ) );
  INV3 U1611 ( .A(\u_decoder/iq_demod/dp_cluster_0/mult_148/SUMB[3][3] ), .Q(
        n705) );
  INV3 U1612 ( .A(\u_decoder/iq_demod/dp_cluster_0/mult_148/CARRYB[3][2] ), 
        .Q(n704) );
  INV3 U1613 ( .A(\u_cordic/mycordic/r173/carry [14]), .Q(n499) );
  INV3 U1614 ( .A(\u_cordic/mycordic/add_262/carry [14]), .Q(n561) );
  NOR21 U1615 ( .A(\u_coder/n315 ), .B(n2196), .Q(\u_coder/N512 ) );
  INV3 U1616 ( .A(\u_coder/N467 ), .Q(n2196) );
  NOR21 U1617 ( .A(n895), .B(n2195), .Q(\u_coder/N513 ) );
  INV3 U1618 ( .A(\u_coder/N468 ), .Q(n2195) );
  INV3 U1619 ( .A(\u_coder/n303 ), .Q(n1936) );
  AOI221 U1620 ( .A(n763), .B(n893), .C(n2156), .D(\u_coder/n105 ), .Q(
        \u_coder/n303 ) );
  INV3 U1621 ( .A(\u_decoder/iq_demod/n55 ), .Q(n2375) );
  AOI221 U1622 ( .A(\u_decoder/iq_demod/add_Q_out [5]), .B(n779), .C(n9), .D(
        \u_decoder/iq_demod/state [1]), .Q(\u_decoder/iq_demod/n55 ) );
  INV3 U1623 ( .A(\u_decoder/iq_demod/n54 ), .Q(n2374) );
  AOI221 U1624 ( .A(\u_decoder/iq_demod/add_Q_out [4]), .B(n779), .C(
        \u_decoder/Q_prefilter [4]), .D(\u_decoder/iq_demod/state [1]), .Q(
        \u_decoder/iq_demod/n54 ) );
  INV3 U1625 ( .A(\u_decoder/iq_demod/n53 ), .Q(n2373) );
  AOI221 U1626 ( .A(\u_decoder/iq_demod/add_Q_out [3]), .B(n779), .C(n7), .D(
        \u_decoder/iq_demod/state [1]), .Q(\u_decoder/iq_demod/n53 ) );
  INV3 U1627 ( .A(\u_decoder/iq_demod/n47 ), .Q(n2304) );
  AOI221 U1628 ( .A(\u_decoder/iq_demod/add_I_out [5]), .B(n779), .C(n10), .D(
        \u_decoder/iq_demod/state [1]), .Q(\u_decoder/iq_demod/n47 ) );
  INV3 U1629 ( .A(\u_decoder/iq_demod/n46 ), .Q(n2303) );
  AOI221 U1630 ( .A(\u_decoder/iq_demod/add_I_out [4]), .B(n779), .C(
        \u_decoder/I_prefilter [4]), .D(\u_decoder/iq_demod/state [1]), .Q(
        \u_decoder/iq_demod/n46 ) );
  INV3 U1631 ( .A(\u_decoder/iq_demod/n45 ), .Q(n2302) );
  AOI221 U1632 ( .A(\u_decoder/iq_demod/add_I_out [3]), .B(n779), .C(n8), .D(
        \u_decoder/iq_demod/state [1]), .Q(\u_decoder/iq_demod/n45 ) );
  NOR21 U1633 ( .A(n2231), .B(n1184), .Q(\u_outFIFO/n403 ) );
  INV3 U1634 ( .A(\u_outFIFO/n661 ), .Q(n2231) );
  NOR21 U1635 ( .A(n2230), .B(n1184), .Q(\u_outFIFO/n401 ) );
  INV3 U1636 ( .A(\u_outFIFO/n666 ), .Q(n2230) );
  NOR21 U1637 ( .A(n2229), .B(n1184), .Q(\u_outFIFO/n399 ) );
  INV3 U1638 ( .A(\u_outFIFO/n664 ), .Q(n2229) );
  NAND22 U1639 ( .A(n1219), .B(\u_inFIFO/n520 ), .Q(\u_inFIFO/n225 ) );
  NOR21 U1640 ( .A(n1150), .B(\u_decoder/fir_filter/n1149 ), .Q(
        \u_decoder/fir_filter/n554 ) );
  NAND22 U1641 ( .A(\u_outFIFO/n659 ), .B(\u_outFIFO/n401 ), .Q(
        \u_outFIFO/n616 ) );
  NAND22 U1642 ( .A(\u_outFIFO/n659 ), .B(\u_outFIFO/n399 ), .Q(
        \u_outFIFO/n614 ) );
  NAND22 U1643 ( .A(\u_outFIFO/n659 ), .B(\u_outFIFO/n403 ), .Q(
        \u_outFIFO/n618 ) );
  XOR21 U1644 ( .A(n1192), .B(n10), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r167/SUMB[7][4] ) );
  XOR21 U1645 ( .A(n1194), .B(n9), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r180/SUMB[7][4] ) );
  XOR21 U1646 ( .A(n1192), .B(n6), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r167/SUMB[7][5] ) );
  XOR21 U1647 ( .A(n1194), .B(n5), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r180/SUMB[7][5] ) );
  XOR21 U1648 ( .A(n1192), .B(n18), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r165/SUMB[7][4] ) );
  XOR21 U1649 ( .A(n1194), .B(n19), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r178/SUMB[7][4] ) );
  XOR21 U1650 ( .A(n1193), .B(n18), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r164/SUMB[7][3] ) );
  XOR21 U1651 ( .A(n1195), .B(n19), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r177/SUMB[7][3] ) );
  NAND22 U1652 ( .A(\u_coder/n206 ), .B(n2177), .Q(\u_coder/n218 ) );
  NOR21 U1653 ( .A(\u_coder/n183 ), .B(\u_coder/n218 ), .Q(\u_coder/n209 ) );
  NAND22 U1654 ( .A(n2639), .B(\u_decoder/fir_filter/n1153 ), .Q(
        \u_decoder/fir_filter/n721 ) );
  INV3 U1655 ( .A(\u_decoder/fir_filter/n1149 ), .Q(n2639) );
  INV3 U1656 ( .A(n198), .Q(n1198) );
  INV3 U1657 ( .A(n198), .Q(n1199) );
  INV3 U1658 ( .A(n198), .Q(n1197) );
  INV3 U1659 ( .A(n198), .Q(n1196) );
  AOI211 U1660 ( .A(\u_coder/n195 ), .B(\u_coder/n194 ), .C(n2151), .Q(
        \u_coder/n184 ) );
  INV3 U1661 ( .A(\u_coder/n192 ), .Q(n2151) );
  INV3 U1662 ( .A(\u_outFIFO/n1110 ), .Q(n1795) );
  NOR21 U1663 ( .A(\u_outFIFO/n315 ), .B(n1184), .Q(\u_outFIFO/n1110 ) );
  NOR21 U1664 ( .A(\u_coder/n194 ), .B(n2153), .Q(\u_coder/n216 ) );
  NOR21 U1665 ( .A(\u_coder/n159 ), .B(\u_coder/n256 ), .Q(\u_coder/n251 ) );
  INV3 U1666 ( .A(\u_cordic/mycordic/n377 ), .Q(n1474) );
  AOI221 U1667 ( .A(\u_cordic/mycordic/N321 ), .B(n772), .C(
        \u_cordic/mycordic/N353 ), .D(n1904), .Q(\u_cordic/mycordic/n377 ) );
  INV3 U1668 ( .A(\u_cordic/mycordic/n376 ), .Q(n1475) );
  AOI221 U1669 ( .A(\u_cordic/mycordic/N322 ), .B(n772), .C(
        \u_cordic/mycordic/N354 ), .D(n1904), .Q(\u_cordic/mycordic/n376 ) );
  INV3 U1670 ( .A(\u_cordic/mycordic/n337 ), .Q(n1483) );
  AOI221 U1671 ( .A(\u_cordic/mycordic/N330 ), .B(n772), .C(
        \u_cordic/mycordic/N362 ), .D(n1904), .Q(\u_cordic/mycordic/n337 ) );
  INV3 U1672 ( .A(\u_cordic/mycordic/n366 ), .Q(n1537) );
  AOI221 U1673 ( .A(\u_cordic/mycordic/N444 ), .B(n777), .C(
        \u_cordic/mycordic/N472 ), .D(n1907), .Q(\u_cordic/mycordic/n366 ) );
  INV3 U1674 ( .A(\u_cordic/mycordic/n541 ), .Q(n1519) );
  AOI221 U1675 ( .A(\u_cordic/mycordic/N454 ), .B(n777), .C(
        \u_cordic/mycordic/N482 ), .D(n1907), .Q(\u_cordic/mycordic/n541 ) );
  INV3 U1676 ( .A(\u_decoder/iq_demod/n44 ), .Q(n2301) );
  AOI221 U1677 ( .A(\u_decoder/iq_demod/add_I_out [2]), .B(n779), .C(n4), .D(
        \u_decoder/iq_demod/state [1]), .Q(\u_decoder/iq_demod/n44 ) );
  INV3 U1678 ( .A(\u_inFIFO/n525 ), .Q(n1818) );
  AOI221 U1679 ( .A(n912), .B(n765), .C(\u_inFIFO/n523 ), .D(\u_inFIFO/N129 ), 
        .Q(\u_inFIFO/n525 ) );
  BUF2 U1680 ( .A(n759), .Q(n1180) );
  AOI221 U1681 ( .A(\u_coder/n194 ), .B(\u_coder/n195 ), .C(n2153), .D(n2184), 
        .Q(\u_coder/n193 ) );
  AOI221 U1682 ( .A(\u_coder/n194 ), .B(\u_coder/n195 ), .C(n2153), .D(n2182), 
        .Q(\u_coder/n202 ) );
  INV3 U1683 ( .A(\u_coder/n201 ), .Q(n2182) );
  NOR21 U1684 ( .A(n1233), .B(\u_coder/n209 ), .Q(\u_coder/n236 ) );
  AOI211 U1685 ( .A(n2154), .B(\u_coder/n155 ), .C(\u_coder/n156 ), .Q(
        \u_coder/n154 ) );
  INV3 U1686 ( .A(\u_coder/n157 ), .Q(n2165) );
  AOI211 U1687 ( .A(n2154), .B(\u_coder/n145 ), .C(\u_coder/n146 ), .Q(
        \u_coder/n143 ) );
  NAND22 U1688 ( .A(\u_coder/n158 ), .B(\u_coder/n147 ), .Q(\u_coder/n169 ) );
  NAND22 U1689 ( .A(\u_coder/n192 ), .B(\u_coder/n217 ), .Q(\u_coder/n212 ) );
  NAND22 U1690 ( .A(\u_coder/n246 ), .B(n2168), .Q(\u_coder/n309 ) );
  NOR21 U1691 ( .A(n194), .B(n16), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[7][4] ) );
  NOR21 U1692 ( .A(n195), .B(n17), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[7][4] ) );
  NOR21 U1693 ( .A(\u_outFIFO/n308 ), .B(\u_outFIFO/n1159 ), .Q(
        \u_outFIFO/n1117 ) );
  AOI211 U1694 ( .A(\u_outFIFO/N1270 ), .B(\u_outFIFO/n1149 ), .C(
        \u_outFIFO/n1154 ), .Q(\u_outFIFO/n1152 ) );
  OAI311 U1695 ( .A(\u_outFIFO/n1155 ), .B(\u_outFIFO/n1156 ), .C(
        \u_outFIFO/n1144 ), .D(n2220), .Q(\u_outFIFO/n1154 ) );
  XNR21 U1696 ( .A(\u_outFIFO/sig_fsm_start_W ), .B(
        \u_outFIFO/sig_fsm_start_R ), .Q(\u_outFIFO/n1156 ) );
  NAND22 U1697 ( .A(\u_outFIFO/n538 ), .B(\u_outFIFO/n399 ), .Q(
        \u_outFIFO/n476 ) );
  NAND22 U1698 ( .A(\u_outFIFO/n469 ), .B(\u_outFIFO/n399 ), .Q(
        \u_outFIFO/n407 ) );
  NAND22 U1699 ( .A(\u_outFIFO/n607 ), .B(\u_outFIFO/n401 ), .Q(
        \u_outFIFO/n547 ) );
  NAND22 U1700 ( .A(\u_outFIFO/n538 ), .B(\u_outFIFO/n401 ), .Q(
        \u_outFIFO/n478 ) );
  NAND22 U1701 ( .A(\u_outFIFO/n469 ), .B(\u_outFIFO/n401 ), .Q(
        \u_outFIFO/n409 ) );
  NAND22 U1702 ( .A(\u_outFIFO/n607 ), .B(\u_outFIFO/n403 ), .Q(
        \u_outFIFO/n549 ) );
  NAND22 U1703 ( .A(\u_outFIFO/n538 ), .B(\u_outFIFO/n403 ), .Q(
        \u_outFIFO/n480 ) );
  NAND22 U1704 ( .A(\u_outFIFO/n469 ), .B(\u_outFIFO/n403 ), .Q(
        \u_outFIFO/n411 ) );
  NOR21 U1705 ( .A(n895), .B(n2197), .Q(\u_coder/N511 ) );
  INV3 U1706 ( .A(\u_coder/N466 ), .Q(n2197) );
  NAND22 U1707 ( .A(\u_outFIFO/n607 ), .B(\u_outFIFO/n399 ), .Q(
        \u_outFIFO/n545 ) );
  INV3 U1708 ( .A(n2707), .Q(n2149) );
  NAND22 U1709 ( .A(n126), .B(n2708), .Q(n2707) );
  NAND22 U1710 ( .A(\u_outFIFO/n403 ), .B(\u_outFIFO/n397 ), .Q(
        \u_outFIFO/n324 ) );
  NAND22 U1711 ( .A(\u_outFIFO/n401 ), .B(\u_outFIFO/n397 ), .Q(
        \u_outFIFO/n322 ) );
  NAND22 U1712 ( .A(\u_outFIFO/n399 ), .B(\u_outFIFO/n397 ), .Q(
        \u_outFIFO/n320 ) );
  INV3 U1713 ( .A(\u_coder/n173 ), .Q(n2096) );
  AOI221 U1714 ( .A(\u_coder/n138 ), .B(\u_coder/n174 ), .C(\u_coder/n174 ), 
        .D(\u_coder/n175 ), .Q(\u_coder/n173 ) );
  NAND22 U1715 ( .A(n2155), .B(\u_coder/n147 ), .Q(\u_coder/n175 ) );
  NOR21 U1716 ( .A(\u_coder/n315 ), .B(n2198), .Q(\u_coder/N510 ) );
  INV3 U1717 ( .A(\u_coder/N465 ), .Q(n2198) );
  NOR21 U1718 ( .A(n895), .B(n2199), .Q(\u_coder/N509 ) );
  INV3 U1719 ( .A(\u_coder/N464 ), .Q(n2199) );
  INV3 U1720 ( .A(\u_inFIFO/n524 ), .Q(n1819) );
  AOI221 U1721 ( .A(n912), .B(n49), .C(\u_inFIFO/n523 ), .D(\u_inFIFO/N130 ), 
        .Q(\u_inFIFO/n524 ) );
  INV3 U1722 ( .A(\u_decoder/iq_demod/n52 ), .Q(n2372) );
  AOI221 U1723 ( .A(\u_decoder/iq_demod/add_Q_out [2]), .B(n779), .C(n3), .D(
        \u_decoder/iq_demod/state [1]), .Q(\u_decoder/iq_demod/n52 ) );
  INV3 U1724 ( .A(\u_cordic/mycordic/n378 ), .Q(n1473) );
  AOI221 U1725 ( .A(\u_cordic/mycordic/N320 ), .B(n772), .C(
        \u_cordic/mycordic/N352 ), .D(n1904), .Q(\u_cordic/mycordic/n378 ) );
  INV3 U1726 ( .A(\u_cordic/mycordic/n339 ), .Q(n1481) );
  AOI221 U1727 ( .A(\u_cordic/mycordic/N328 ), .B(n772), .C(
        \u_cordic/mycordic/N360 ), .D(n1904), .Q(\u_cordic/mycordic/n339 ) );
  INV3 U1728 ( .A(\u_cordic/mycordic/n338 ), .Q(n1482) );
  AOI221 U1729 ( .A(\u_cordic/mycordic/N329 ), .B(n772), .C(
        \u_cordic/mycordic/N361 ), .D(n1904), .Q(\u_cordic/mycordic/n338 ) );
  INV3 U1730 ( .A(\u_cordic/mycordic/n368 ), .Q(n1568) );
  AOI221 U1731 ( .A(\u_cordic/mycordic/N386 ), .B(n778), .C(
        \u_cordic/mycordic/N418 ), .D(n1908), .Q(\u_cordic/mycordic/n368 ) );
  INV3 U1732 ( .A(\u_cordic/mycordic/n369 ), .Q(n1567) );
  AOI221 U1733 ( .A(\u_cordic/mycordic/N385 ), .B(n778), .C(
        \u_cordic/mycordic/N417 ), .D(n1908), .Q(\u_cordic/mycordic/n369 ) );
  INV3 U1734 ( .A(\u_cordic/mycordic/n370 ), .Q(n1566) );
  AOI221 U1735 ( .A(\u_cordic/mycordic/N384 ), .B(n778), .C(
        \u_cordic/mycordic/N416 ), .D(n1908), .Q(\u_cordic/mycordic/n370 ) );
  INV3 U1736 ( .A(\u_cordic/mycordic/n550 ), .Q(n1544) );
  AOI221 U1737 ( .A(\u_cordic/mycordic/N394 ), .B(\u_cordic/mycordic/n332 ), 
        .C(\u_cordic/mycordic/N426 ), .D(n1908), .Q(\u_cordic/mycordic/n550 )
         );
  INV3 U1738 ( .A(\u_cordic/mycordic/n551 ), .Q(n1543) );
  AOI221 U1739 ( .A(\u_cordic/mycordic/N393 ), .B(n778), .C(
        \u_cordic/mycordic/N425 ), .D(n1908), .Q(\u_cordic/mycordic/n551 ) );
  INV3 U1740 ( .A(\u_cordic/mycordic/n552 ), .Q(n1542) );
  AOI221 U1741 ( .A(\u_cordic/mycordic/N392 ), .B(\u_cordic/mycordic/n332 ), 
        .C(\u_cordic/mycordic/N424 ), .D(n1908), .Q(\u_cordic/mycordic/n552 )
         );
  INV3 U1742 ( .A(\u_cordic/mycordic/n365 ), .Q(n1538) );
  AOI221 U1743 ( .A(\u_cordic/mycordic/N445 ), .B(n777), .C(
        \u_cordic/mycordic/N473 ), .D(n1907), .Q(\u_cordic/mycordic/n365 ) );
  INV3 U1744 ( .A(\u_cordic/mycordic/n364 ), .Q(n1539) );
  AOI221 U1745 ( .A(\u_cordic/mycordic/N446 ), .B(n777), .C(
        \u_cordic/mycordic/N474 ), .D(n1907), .Q(\u_cordic/mycordic/n364 ) );
  INV3 U1746 ( .A(\u_cordic/mycordic/n543 ), .Q(n1517) );
  AOI221 U1747 ( .A(\u_cordic/mycordic/N452 ), .B(n777), .C(
        \u_cordic/mycordic/N480 ), .D(n1907), .Q(\u_cordic/mycordic/n543 ) );
  INV3 U1748 ( .A(\u_cordic/mycordic/n542 ), .Q(n1518) );
  AOI221 U1749 ( .A(\u_cordic/mycordic/N453 ), .B(n777), .C(
        \u_cordic/mycordic/N481 ), .D(n1907), .Q(\u_cordic/mycordic/n542 ) );
  NAND22 U1750 ( .A(\u_inFIFO/n474 ), .B(\u_inFIFO/n475 ), .Q(\u_inFIFO/n226 )
         );
  NAND22 U1751 ( .A(\u_inFIFO/n484 ), .B(\u_inFIFO/n475 ), .Q(\u_inFIFO/n236 )
         );
  NAND22 U1752 ( .A(\u_inFIFO/n481 ), .B(\u_inFIFO/n475 ), .Q(\u_inFIFO/n233 )
         );
  NAND22 U1753 ( .A(\u_inFIFO/n478 ), .B(\u_inFIFO/n475 ), .Q(\u_inFIFO/n230 )
         );
  NAND22 U1754 ( .A(\u_inFIFO/n505 ), .B(\u_inFIFO/n474 ), .Q(\u_inFIFO/n263 )
         );
  NAND22 U1755 ( .A(\u_inFIFO/n496 ), .B(\u_inFIFO/n474 ), .Q(\u_inFIFO/n251 )
         );
  NAND22 U1756 ( .A(\u_inFIFO/n487 ), .B(\u_inFIFO/n474 ), .Q(\u_inFIFO/n239 )
         );
  NAND22 U1757 ( .A(\u_inFIFO/n505 ), .B(\u_inFIFO/n481 ), .Q(\u_inFIFO/n269 )
         );
  NAND22 U1758 ( .A(\u_inFIFO/n496 ), .B(\u_inFIFO/n481 ), .Q(\u_inFIFO/n257 )
         );
  NAND22 U1759 ( .A(\u_inFIFO/n487 ), .B(\u_inFIFO/n481 ), .Q(\u_inFIFO/n245 )
         );
  NAND22 U1760 ( .A(\u_inFIFO/n505 ), .B(\u_inFIFO/n478 ), .Q(\u_inFIFO/n266 )
         );
  NAND22 U1761 ( .A(\u_inFIFO/n496 ), .B(\u_inFIFO/n478 ), .Q(\u_inFIFO/n254 )
         );
  NAND22 U1762 ( .A(\u_inFIFO/n487 ), .B(\u_inFIFO/n478 ), .Q(\u_inFIFO/n242 )
         );
  NAND22 U1763 ( .A(\u_inFIFO/n505 ), .B(\u_inFIFO/n484 ), .Q(\u_inFIFO/n272 )
         );
  NAND22 U1764 ( .A(\u_inFIFO/n496 ), .B(\u_inFIFO/n484 ), .Q(\u_inFIFO/n260 )
         );
  NAND22 U1765 ( .A(\u_inFIFO/n487 ), .B(\u_inFIFO/n484 ), .Q(\u_inFIFO/n248 )
         );
  NOR31 U1766 ( .A(\u_inFIFO/n549 ), .B(n1238), .C(\u_inFIFO/n550 ), .Q(
        \u_inFIFO/n534 ) );
  NAND22 U1767 ( .A(n1219), .B(\u_coder/n314 ), .Q(n895) );
  NAND22 U1768 ( .A(n1219), .B(\u_coder/n314 ), .Q(\u_coder/n315 ) );
  NAND22 U1769 ( .A(\u_outFIFO/n1128 ), .B(\u_outFIFO/n1129 ), .Q(
        \u_outFIFO/n1120 ) );
  NOR21 U1770 ( .A(\u_outFIFO/n1139 ), .B(n1796), .Q(\u_outFIFO/n1131 ) );
  NAND22 U1771 ( .A(n1219), .B(\u_outFIFO/n1115 ), .Q(\u_outFIFO/n1113 ) );
  NAND31 U1772 ( .A(n290), .B(n50), .C(n2099), .Q(\u_cdr/n30 ) );
  NAND22 U1773 ( .A(n1218), .B(n3114), .Q(\u_cdr/n44 ) );
  NAND22 U1774 ( .A(\u_outFIFO/n659 ), .B(\u_outFIFO/n661 ), .Q(
        \u_outFIFO/n669 ) );
  INV3 U1775 ( .A(\u_outFIFO/n1139 ), .Q(n1797) );
  NAND22 U1776 ( .A(\u_outFIFO/n659 ), .B(\u_outFIFO/n664 ), .Q(
        \u_outFIFO/n674 ) );
  NAND22 U1777 ( .A(\u_outFIFO/n659 ), .B(\u_outFIFO/n666 ), .Q(
        \u_outFIFO/n677 ) );
  NOR21 U1778 ( .A(\u_cdr/n38 ), .B(n1238), .Q(\u_cdr/n33 ) );
  AOI2111 U1779 ( .A(\u_coder/j [0]), .B(\u_coder/j [3]), .C(\u_coder/n206 ), 
        .D(n762), .Q(\u_coder/n200 ) );
  BUF2 U1780 ( .A(n759), .Q(n1176) );
  BUF2 U1781 ( .A(n759), .Q(n1177) );
  BUF2 U1782 ( .A(n759), .Q(n1178) );
  BUF2 U1783 ( .A(n759), .Q(n1179) );
  NOR21 U1784 ( .A(n1234), .B(\u_outFIFO/n311 ), .Q(\u_outFIFO/n310 ) );
  NAND22 U1785 ( .A(\u_inFIFO/n552 ), .B(\u_inFIFO/n553 ), .Q(\u_inFIFO/n549 )
         );
  NAND22 U1786 ( .A(n2141), .B(n1212), .Q(\u_inFIFO/n551 ) );
  INV3 U1787 ( .A(\u_inFIFO/n520 ), .Q(n2141) );
  INV3 U1788 ( .A(\u_coder/n283 ), .Q(n2169) );
  NAND22 U1789 ( .A(n2170), .B(n2185), .Q(\u_coder/n283 ) );
  INV3 U1790 ( .A(\u_outFIFO/n315 ), .Q(n1911) );
  NAND31 U1791 ( .A(\u_inFIFO/n550 ), .B(\u_inFIFO/n520 ), .C(n912), .Q(
        \u_inFIFO/n552 ) );
  INV3 U1792 ( .A(\u_cordic/mycordic/n380 ), .Q(n1471) );
  AOI221 U1793 ( .A(\u_cordic/mycordic/N318 ), .B(n772), .C(
        \u_cordic/mycordic/N350 ), .D(n1904), .Q(\u_cordic/mycordic/n380 ) );
  INV3 U1794 ( .A(\u_cordic/mycordic/n385 ), .Q(n1488) );
  AOI221 U1795 ( .A(n1905), .B(\u_cordic/mycordic/N289 ), .C(n773), .D(
        \u_cordic/mycordic/N257 ), .Q(\u_cordic/mycordic/n385 ) );
  INV3 U1796 ( .A(\u_cordic/mycordic/n384 ), .Q(n1489) );
  AOI221 U1797 ( .A(n1905), .B(\u_cordic/mycordic/N290 ), .C(n773), .D(
        \u_cordic/mycordic/N258 ), .Q(\u_cordic/mycordic/n384 ) );
  NOR21 U1798 ( .A(n194), .B(n18), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[7][5] ) );
  NOR21 U1799 ( .A(n195), .B(n19), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[7][5] ) );
  INV3 U1800 ( .A(\u_coder/n183 ), .Q(n2185) );
  INV3 U1801 ( .A(\u_inFIFO/n527 ), .Q(n1816) );
  AOI221 U1802 ( .A(n912), .B(n15), .C(\u_inFIFO/n523 ), .D(\u_inFIFO/N127 ), 
        .Q(\u_inFIFO/n527 ) );
  INV3 U1803 ( .A(\u_inFIFO/n526 ), .Q(n1817) );
  AOI221 U1804 ( .A(n912), .B(n1202), .C(\u_inFIFO/n523 ), .D(\u_inFIFO/N128 ), 
        .Q(\u_inFIFO/n526 ) );
  INV3 U1805 ( .A(\u_inFIFO/n528 ), .Q(n1815) );
  AOI221 U1806 ( .A(n912), .B(\u_inFIFO/N38 ), .C(\u_inFIFO/n523 ), .D(
        \u_inFIFO/N126 ), .Q(\u_inFIFO/n528 ) );
  NAND22 U1807 ( .A(n2174), .B(n2185), .Q(\u_coder/n235 ) );
  INV3 U1808 ( .A(\u_coder/n325 ), .Q(n2176) );
  NAND31 U1809 ( .A(n2177), .B(\u_coder/n190 ), .C(\u_coder/j [0]), .Q(
        \u_coder/n325 ) );
  INV3 U1810 ( .A(\u_coder/n144 ), .Q(n2168) );
  INV3 U1811 ( .A(\u_outFIFO/n391 ), .Q(n876) );
  NAND22 U1812 ( .A(\u_outFIFO/n1085 ), .B(\u_outFIFO/n1001 ), .Q(
        \u_outFIFO/n391 ) );
  INV3 U1813 ( .A(\u_outFIFO/n386 ), .Q(n874) );
  NAND22 U1814 ( .A(\u_outFIFO/n1085 ), .B(\u_outFIFO/n992 ), .Q(
        \u_outFIFO/n386 ) );
  XNR21 U1815 ( .A(n2209), .B(\u_cdr/n48 ), .Q(\u_cdr/n46 ) );
  INV3 U1816 ( .A(\u_cdr/dp_cluster_0/mult_add_59_aco/PROD_not[3] ), .Q(n2209)
         );
  NOR21 U1817 ( .A(\u_cdr/n49 ), .B(
        \u_cdr/dp_cluster_0/mult_add_59_aco/PROD_not[2] ), .Q(\u_cdr/n48 ) );
  NAND22 U1818 ( .A(n2211), .B(n2210), .Q(\u_cdr/n49 ) );
  XOR21 U1819 ( .A(n2211), .B(\u_cdr/dp_cluster_0/mult_add_59_aco/PROD_not[0] ), .Q(n371) );
  BUF2 U1820 ( .A(n764), .Q(n1200) );
  OAI311 U1821 ( .A(n289), .B(\u_cdr/n30 ), .C(n20), .D(n1220), .Q(\u_cdr/n45 ) );
  BUF2 U1822 ( .A(\u_inFIFO/n227 ), .Q(n896) );
  BUF2 U1823 ( .A(\u_inFIFO/n227 ), .Q(n897) );
  NAND22 U1824 ( .A(n2099), .B(\u_cdr/n43 ), .Q(\u_cdr/n39 ) );
  INV3 U1825 ( .A(\u_coder/n305 ), .Q(n2156) );
  NAND22 U1826 ( .A(n2157), .B(n2168), .Q(\u_coder/n305 ) );
  XNR21 U1827 ( .A(\u_cdr/dp_cluster_0/mult_add_59_aco/PROD_not[2] ), .B(
        \u_cdr/n49 ), .Q(n372) );
  BUF2 U1828 ( .A(\u_inFIFO/n473 ), .Q(n910) );
  BUF2 U1829 ( .A(\u_inFIFO/n473 ), .Q(n911) );
  BUF2 U1830 ( .A(\u_inFIFO/n440 ), .Q(n908) );
  BUF2 U1831 ( .A(\u_inFIFO/n440 ), .Q(n909) );
  BUF2 U1832 ( .A(\u_inFIFO/n407 ), .Q(n906) );
  BUF2 U1833 ( .A(\u_inFIFO/n407 ), .Q(n907) );
  BUF2 U1834 ( .A(\u_inFIFO/n374 ), .Q(n904) );
  BUF2 U1835 ( .A(\u_inFIFO/n374 ), .Q(n905) );
  BUF2 U1836 ( .A(\u_inFIFO/n341 ), .Q(n902) );
  BUF2 U1837 ( .A(\u_inFIFO/n341 ), .Q(n903) );
  BUF2 U1838 ( .A(\u_inFIFO/n308 ), .Q(n900) );
  BUF2 U1839 ( .A(\u_inFIFO/n308 ), .Q(n901) );
  BUF2 U1840 ( .A(\u_inFIFO/n275 ), .Q(n898) );
  BUF2 U1841 ( .A(\u_inFIFO/n275 ), .Q(n899) );
  BUF2 U1842 ( .A(n760), .Q(n1181) );
  NOR21 U1843 ( .A(n2162), .B(\u_coder/n148 ), .Q(\u_coder/n247 ) );
  INV3 U1844 ( .A(\u_outFIFO/n331 ), .Q(n841) );
  NAND22 U1845 ( .A(\u_outFIFO/n1001 ), .B(\u_outFIFO/n983 ), .Q(
        \u_outFIFO/n331 ) );
  NOR21 U1846 ( .A(\u_cordic/mycordic/present_Q_table[0][5] ), .B(n564), .Q(
        \u_cordic/mycordic/sub_add_151_b0/carry [6]) );
  INV3 U1847 ( .A(\u_cordic/mycordic/sub_add_151_b0/carry [5]), .Q(n564) );
  INV3 U1848 ( .A(\u_outFIFO/n381 ), .Q(n872) );
  NAND22 U1849 ( .A(\u_outFIFO/n1085 ), .B(\u_outFIFO/n982 ), .Q(
        \u_outFIFO/n381 ) );
  INV3 U1850 ( .A(\u_cordic/mycordic/n587 ), .Q(n766) );
  NAND22 U1851 ( .A(\u_outFIFO/n1010 ), .B(\u_outFIFO/n983 ), .Q(n843) );
  NAND22 U1852 ( .A(\u_outFIFO/n1010 ), .B(\u_outFIFO/n983 ), .Q(
        \u_outFIFO/n336 ) );
  INV3 U1853 ( .A(\u_inFIFO/n550 ), .Q(n2146) );
  NAND22 U1854 ( .A(\u_outFIFO/n992 ), .B(\u_outFIFO/n983 ), .Q(
        \u_outFIFO/n326 ) );
  NAND22 U1855 ( .A(\u_outFIFO/n963 ), .B(\u_outFIFO/n664 ), .Q(
        \u_outFIFO/n842 ) );
  NAND22 U1856 ( .A(\u_outFIFO/n830 ), .B(\u_outFIFO/n664 ), .Q(
        \u_outFIFO/n709 ) );
  NAND22 U1857 ( .A(\u_outFIFO/n1104 ), .B(\u_outFIFO/n666 ), .Q(
        \u_outFIFO/n978 ) );
  NAND22 U1858 ( .A(\u_outFIFO/n963 ), .B(\u_outFIFO/n666 ), .Q(
        \u_outFIFO/n845 ) );
  NAND22 U1859 ( .A(\u_outFIFO/n830 ), .B(\u_outFIFO/n666 ), .Q(
        \u_outFIFO/n712 ) );
  NAND22 U1860 ( .A(\u_outFIFO/n1052 ), .B(\u_outFIFO/n1010 ), .Q(
        \u_outFIFO/n376 ) );
  NAND22 U1861 ( .A(\u_outFIFO/n1019 ), .B(\u_outFIFO/n1010 ), .Q(
        \u_outFIFO/n356 ) );
  NAND22 U1862 ( .A(\u_outFIFO/n1104 ), .B(\u_outFIFO/n661 ), .Q(
        \u_outFIFO/n981 ) );
  NAND22 U1863 ( .A(\u_outFIFO/n963 ), .B(\u_outFIFO/n661 ), .Q(
        \u_outFIFO/n848 ) );
  NAND22 U1864 ( .A(\u_outFIFO/n830 ), .B(\u_outFIFO/n661 ), .Q(
        \u_outFIFO/n715 ) );
  NAND22 U1865 ( .A(\u_outFIFO/n1052 ), .B(\u_outFIFO/n982 ), .Q(
        \u_outFIFO/n361 ) );
  NAND22 U1866 ( .A(\u_outFIFO/n1019 ), .B(\u_outFIFO/n982 ), .Q(
        \u_outFIFO/n341 ) );
  NAND22 U1867 ( .A(\u_outFIFO/n1052 ), .B(\u_outFIFO/n1001 ), .Q(
        \u_outFIFO/n371 ) );
  NAND22 U1868 ( .A(\u_outFIFO/n1019 ), .B(\u_outFIFO/n1001 ), .Q(
        \u_outFIFO/n351 ) );
  NAND22 U1869 ( .A(\u_outFIFO/n1052 ), .B(\u_outFIFO/n992 ), .Q(
        \u_outFIFO/n366 ) );
  NAND22 U1870 ( .A(\u_outFIFO/n1019 ), .B(\u_outFIFO/n992 ), .Q(
        \u_outFIFO/n346 ) );
  INV3 U1871 ( .A(\u_outFIFO/n317 ), .Q(n836) );
  NAND22 U1872 ( .A(\u_outFIFO/n982 ), .B(\u_outFIFO/n983 ), .Q(
        \u_outFIFO/n317 ) );
  NAND22 U1873 ( .A(\u_outFIFO/n659 ), .B(\u_outFIFO/N198 ), .Q(
        \u_outFIFO/n612 ) );
  NOR21 U1874 ( .A(\u_coder/n315 ), .B(n2205), .Q(\u_coder/N504 ) );
  INV3 U1875 ( .A(\u_coder/N459 ), .Q(n2205) );
  NOR21 U1876 ( .A(n895), .B(n2204), .Q(\u_coder/N505 ) );
  INV3 U1877 ( .A(\u_coder/N460 ), .Q(n2204) );
  NOR21 U1878 ( .A(\u_coder/n315 ), .B(n2203), .Q(\u_coder/N506 ) );
  INV3 U1879 ( .A(\u_coder/N461 ), .Q(n2203) );
  NOR21 U1880 ( .A(\u_coder/n315 ), .B(n2200), .Q(\u_coder/N508 ) );
  INV3 U1881 ( .A(\u_coder/N463 ), .Q(n2200) );
  INV3 U1882 ( .A(n3114), .Q(n2099) );
  INV3 U1883 ( .A(\u_outFIFO/n396 ), .Q(n888) );
  NAND22 U1884 ( .A(\u_outFIFO/n1085 ), .B(\u_outFIFO/n1010 ), .Q(
        \u_outFIFO/n396 ) );
  NAND22 U1885 ( .A(\u_outFIFO/n1104 ), .B(\u_outFIFO/n664 ), .Q(
        \u_outFIFO/n975 ) );
  INV3 U1886 ( .A(\u_coder/n195 ), .Q(n2097) );
  INV3 U1887 ( .A(\u_coder/n217 ), .Q(n2153) );
  INV3 U1888 ( .A(\u_coder/n190 ), .Q(n2184) );
  NAND22 U1889 ( .A(\u_outFIFO/n469 ), .B(\u_outFIFO/N198 ), .Q(
        \u_outFIFO/n405 ) );
  NAND22 U1890 ( .A(\u_outFIFO/n538 ), .B(\u_outFIFO/N198 ), .Q(
        \u_outFIFO/n474 ) );
  NAND22 U1891 ( .A(\u_outFIFO/n830 ), .B(\u_outFIFO/N198 ), .Q(
        \u_outFIFO/n706 ) );
  NAND22 U1892 ( .A(\u_outFIFO/n607 ), .B(\u_outFIFO/N198 ), .Q(
        \u_outFIFO/n543 ) );
  NAND22 U1893 ( .A(\u_outFIFO/n1104 ), .B(\u_outFIFO/N198 ), .Q(
        \u_outFIFO/n972 ) );
  NAND22 U1894 ( .A(\u_outFIFO/n963 ), .B(\u_outFIFO/N198 ), .Q(
        \u_outFIFO/n839 ) );
  NOR21 U1895 ( .A(\u_cordic/mycordic/present_Q_table[0][6] ), .B(n565), .Q(
        \u_cordic/mycordic/sub_add_151_b0/carry [7]) );
  INV3 U1896 ( .A(\u_cordic/mycordic/sub_add_151_b0/carry [6]), .Q(n565) );
  INV3 U1897 ( .A(\u_cdr/dp_cluster_0/mult_add_59_aco/PROD_not[0] ), .Q(n2210)
         );
  NAND22 U1898 ( .A(\u_outFIFO/N198 ), .B(\u_outFIFO/n397 ), .Q(
        \u_outFIFO/n318 ) );
  INV3 U1899 ( .A(\u_coder/n150 ), .Q(n2167) );
  INV3 U1900 ( .A(n2764), .Q(n2224) );
  INV3 U1901 ( .A(\u_outFIFO/n1115 ), .Q(n2217) );
  INV3 U1902 ( .A(\u_outFIFO/n1159 ), .Q(n2218) );
  INV3 U1903 ( .A(\u_coder/n158 ), .Q(n2154) );
  NOR21 U1904 ( .A(n194), .B(n6), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r164/CARRYB[7][3] ) );
  NOR21 U1905 ( .A(n195), .B(n5), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r177/CARRYB[7][3] ) );
  NOR21 U1906 ( .A(n194), .B(n6), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r165/CARRYB[7][4] ) );
  NOR21 U1907 ( .A(n195), .B(n5), .Q(
        \u_decoder/fir_filter/dp_cluster_0/r178/CARRYB[7][4] ) );
  NOR21 U1908 ( .A(\u_cordic/mycordic/present_Q_table[0][4] ), .B(
        \u_cordic/mycordic/present_Q_table[0][3] ), .Q(
        \u_cordic/mycordic/sub_add_151_b0/carry [5]) );
  NOR21 U1909 ( .A(n895), .B(n2201), .Q(\u_coder/N507 ) );
  INV3 U1910 ( .A(\u_coder/N462 ), .Q(n2201) );
  NAND22 U1911 ( .A(n2159), .B(n2168), .Q(\u_coder/n223 ) );
  INV3 U1912 ( .A(\u_coder/n242 ), .Q(n2159) );
  BUF2 U1913 ( .A(n760), .Q(n1182) );
  INV3 U1914 ( .A(\u_cordic/mycordic/n348 ), .Q(n1492) );
  AOI221 U1915 ( .A(n1905), .B(\u_cordic/mycordic/N256 ), .C(n774), .D(
        \u_cordic/mycordic/N264 ), .Q(\u_cordic/mycordic/n348 ) );
  INV3 U1916 ( .A(\u_cordic/mycordic/n347 ), .Q(n1493) );
  AOI221 U1917 ( .A(n1905), .B(\u_cordic/mycordic/N257 ), .C(n774), .D(
        \u_cordic/mycordic/N265 ), .Q(\u_cordic/mycordic/n347 ) );
  INV3 U1918 ( .A(\u_cordic/mycordic/n346 ), .Q(n1494) );
  AOI221 U1919 ( .A(n1905), .B(\u_cordic/mycordic/N258 ), .C(n774), .D(
        \u_cordic/mycordic/N266 ), .Q(\u_cordic/mycordic/n346 ) );
  INV3 U1920 ( .A(\u_cordic/mycordic/n386 ), .Q(n1487) );
  AOI221 U1921 ( .A(n1905), .B(\u_cordic/mycordic/N288 ), .C(n773), .D(
        \u_cordic/mycordic/N256 ), .Q(\u_cordic/mycordic/n386 ) );
  BUF2 U1922 ( .A(n764), .Q(n1201) );
  INV3 U1923 ( .A(n2760), .Q(n2227) );
  NAND22 U1924 ( .A(n161), .B(n2761), .Q(n2760) );
  INV3 U1925 ( .A(\u_decoder/iq_demod/n51 ), .Q(n2370) );
  AOI221 U1926 ( .A(\u_decoder/iq_demod/add_Q_out [1]), .B(n779), .C(n11), .D(
        \u_decoder/iq_demod/state [1]), .Q(\u_decoder/iq_demod/n51 ) );
  INV3 U1927 ( .A(\u_decoder/iq_demod/n43 ), .Q(n2299) );
  AOI221 U1928 ( .A(\u_decoder/iq_demod/add_I_out [1]), .B(n779), .C(n12), .D(
        \u_decoder/iq_demod/state [1]), .Q(\u_decoder/iq_demod/n43 ) );
  INV3 U1929 ( .A(\u_cordic/mycordic/n342 ), .Q(n1478) );
  AOI221 U1930 ( .A(\u_cordic/mycordic/N325 ), .B(\u_cordic/mycordic/n336 ), 
        .C(\u_cordic/mycordic/N357 ), .D(n1904), .Q(\u_cordic/mycordic/n342 )
         );
  INV3 U1931 ( .A(\u_cordic/mycordic/n331 ), .Q(n1572) );
  AOI221 U1932 ( .A(\u_cordic/mycordic/N390 ), .B(\u_cordic/mycordic/n332 ), 
        .C(\u_cordic/mycordic/N422 ), .D(n1908), .Q(\u_cordic/mycordic/n331 )
         );
  INV3 U1933 ( .A(\u_cordic/mycordic/n372 ), .Q(n1564) );
  AOI221 U1934 ( .A(\u_cordic/mycordic/N382 ), .B(\u_cordic/mycordic/n332 ), 
        .C(\u_cordic/mycordic/N414 ), .D(n1908), .Q(\u_cordic/mycordic/n372 )
         );
  INV3 U1935 ( .A(\u_cordic/mycordic/n379 ), .Q(n1472) );
  AOI221 U1936 ( .A(\u_cordic/mycordic/N319 ), .B(\u_cordic/mycordic/n336 ), 
        .C(\u_cordic/mycordic/N351 ), .D(n1904), .Q(\u_cordic/mycordic/n379 )
         );
  INV3 U1937 ( .A(\u_cordic/mycordic/n341 ), .Q(n1479) );
  AOI221 U1938 ( .A(\u_cordic/mycordic/N326 ), .B(n772), .C(
        \u_cordic/mycordic/N358 ), .D(n1904), .Q(\u_cordic/mycordic/n341 ) );
  INV3 U1939 ( .A(\u_cordic/mycordic/n340 ), .Q(n1480) );
  AOI221 U1940 ( .A(\u_cordic/mycordic/N327 ), .B(\u_cordic/mycordic/n336 ), 
        .C(\u_cordic/mycordic/N359 ), .D(n1904), .Q(\u_cordic/mycordic/n340 )
         );
  INV3 U1941 ( .A(\u_cordic/mycordic/n371 ), .Q(n1565) );
  AOI221 U1942 ( .A(\u_cordic/mycordic/N383 ), .B(n778), .C(
        \u_cordic/mycordic/N415 ), .D(n1908), .Q(\u_cordic/mycordic/n371 ) );
  INV3 U1943 ( .A(\u_cordic/mycordic/n553 ), .Q(n1541) );
  AOI221 U1944 ( .A(\u_cordic/mycordic/N391 ), .B(n778), .C(
        \u_cordic/mycordic/N423 ), .D(n1908), .Q(\u_cordic/mycordic/n553 ) );
  INV3 U1945 ( .A(\u_cordic/mycordic/n544 ), .Q(n1516) );
  AOI221 U1946 ( .A(\u_cordic/mycordic/N451 ), .B(\u_cordic/mycordic/n363 ), 
        .C(\u_cordic/mycordic/N479 ), .D(n1907), .Q(\u_cordic/mycordic/n544 )
         );
  INV3 U1947 ( .A(\u_cordic/mycordic/n333 ), .Q(n1571) );
  AOI221 U1948 ( .A(\u_cordic/mycordic/N389 ), .B(n778), .C(
        \u_cordic/mycordic/N421 ), .D(n1908), .Q(\u_cordic/mycordic/n333 ) );
  INV3 U1949 ( .A(\u_cordic/mycordic/n546 ), .Q(n1514) );
  AOI221 U1950 ( .A(\u_cordic/mycordic/N449 ), .B(\u_cordic/mycordic/n363 ), 
        .C(\u_cordic/mycordic/N477 ), .D(n1907), .Q(\u_cordic/mycordic/n546 )
         );
  INV3 U1951 ( .A(\u_cordic/mycordic/n545 ), .Q(n1515) );
  AOI221 U1952 ( .A(\u_cordic/mycordic/N450 ), .B(n777), .C(
        \u_cordic/mycordic/N478 ), .D(n1907), .Q(\u_cordic/mycordic/n545 ) );
  NOR21 U1953 ( .A(\u_cordic/n19 ), .B(\u_cordic/n15 ), .Q(\u_cordic/n18 ) );
  NOR21 U1954 ( .A(n1234), .B(n912), .Q(\u_inFIFO/n523 ) );
  INV3 U1955 ( .A(\u_outFIFO/n1129 ), .Q(n1912) );
  NAND22 U1956 ( .A(\u_inFIFO/n215 ), .B(\u_inFIFO/n212 ), .Q(\u_inFIFO/n531 )
         );
  INV3 U1957 ( .A(\u_inFIFO/n553 ), .Q(n2094) );
  NAND22 U1958 ( .A(\u_decoder/iq_demod/cossin_dig/n37 ), .B(
        \u_decoder/iq_demod/cossin_dig/n26 ), .Q(
        \u_decoder/iq_demod/cossin_dig/n31 ) );
  BUF2 U1959 ( .A(\u_cordic/mycordic/n332 ), .Q(n778) );
  BUF2 U1960 ( .A(\u_cordic/mycordic/n336 ), .Q(n772) );
  INV3 U1961 ( .A(\u_cordic/mycordic/n387 ), .Q(n1486) );
  AOI221 U1962 ( .A(n1905), .B(\u_cordic/mycordic/N287 ), .C(n773), .D(
        \u_cordic/mycordic/N255 ), .Q(\u_cordic/mycordic/n387 ) );
  NAND22 U1963 ( .A(n1218), .B(\u_decoder/iq_demod/cossin_dig/n26 ), .Q(
        \u_decoder/iq_demod/cossin_dig/n42 ) );
  NAND22 U1964 ( .A(n2142), .B(\u_inFIFO/n212 ), .Q(\u_inFIFO/n564 ) );
  NOR21 U1965 ( .A(\u_outFIFO/n1155 ), .B(\u_outFIFO/n308 ), .Q(
        \u_outFIFO/n1149 ) );
  NOR21 U1966 ( .A(\u_cordic/mycordic/present_I_table[0][5] ), .B(n562), .Q(
        \u_cordic/mycordic/sub_add_150_b0/carry [6]) );
  INV3 U1967 ( .A(\u_cordic/mycordic/sub_add_150_b0/carry [5]), .Q(n562) );
  NOR21 U1968 ( .A(\u_cordic/mycordic/present_I_table[0][4] ), .B(
        \u_cordic/mycordic/present_I_table[0][3] ), .Q(
        \u_cordic/mycordic/sub_add_150_b0/carry [5]) );
  NOR21 U1969 ( .A(\u_coder/n190 ), .B(\u_coder/j [3]), .Q(\u_coder/n189 ) );
  NAND22 U1970 ( .A(\u_inFIFO/n563 ), .B(\u_inFIFO/n564 ), .Q(\u_inFIFO/n561 )
         );
  NOR21 U1971 ( .A(n1236), .B(\u_cordic/mycordic/present_Q_table[4][7] ), .Q(
        \u_cordic/mycordic/n363 ) );
  INV3 U1972 ( .A(\u_outFIFO/n1142 ), .Q(n1796) );
  AOI211 U1973 ( .A(\u_decoder/fir_filter/n1153 ), .B(
        \u_decoder/fir_filter/n1154 ), .C(n1240), .Q(
        \u_decoder/fir_filter/N11 ) );
  NAND22 U1974 ( .A(\u_decoder/fir_filter/n1151 ), .B(n294), .Q(
        \u_decoder/fir_filter/n1154 ) );
  INV3 U1975 ( .A(\u_cordic/mycordic/n391 ), .Q(n1901) );
  INV3 U1976 ( .A(\u_inFIFO/n568 ), .Q(n2142) );
  BUF2 U1977 ( .A(\u_cordic/mycordic/n345 ), .Q(n774) );
  BUF2 U1978 ( .A(\u_cordic/mycordic/n438 ), .Q(n770) );
  BUF2 U1979 ( .A(\u_cordic/mycordic/n438 ), .Q(n771) );
  BUF2 U1980 ( .A(\u_cordic/mycordic/n345 ), .Q(n773) );
  INV3 U1981 ( .A(n3074), .Q(n1842) );
  NAND22 U1982 ( .A(n1218), .B(n2101), .Q(n3074) );
  INV3 U1983 ( .A(n775), .Q(n776) );
  INV3 U1984 ( .A(\u_outFIFO/n1147 ), .Q(n2220) );
  INV3 U1985 ( .A(\u_coder/n314 ), .Q(n2186) );
  INV3 U1986 ( .A(\u_outFIFO/n1148 ), .Q(n2219) );
  NOR21 U1987 ( .A(\u_cordic/mycordic/present_I_table[0][6] ), .B(n563), .Q(
        \u_cordic/mycordic/sub_add_150_b0/carry [7]) );
  INV3 U1988 ( .A(\u_cordic/mycordic/sub_add_150_b0/carry [6]), .Q(n563) );
  NAND22 U1989 ( .A(n1847), .B(\u_decoder/iq_demod/cossin_dig/n37 ), .Q(
        \u_decoder/iq_demod/cossin_dig/n40 ) );
  INV3 U1990 ( .A(\u_decoder/iq_demod/cossin_dig/n42 ), .Q(n1847) );
  INV3 U1991 ( .A(\u_cdr/phd1/n15 ), .Q(n2689) );
  INV3 U1992 ( .A(\u_cordic/mycordic/n349 ), .Q(n1491) );
  AOI221 U1993 ( .A(n1905), .B(\u_cordic/mycordic/N255 ), .C(n774), .D(
        \u_cordic/mycordic/N263 ), .Q(\u_cordic/mycordic/n349 ) );
  INV3 U1994 ( .A(\u_decoder/iq_demod/n50 ), .Q(n2345) );
  AOI221 U1995 ( .A(\u_decoder/iq_demod/add_Q_out [0]), .B(n779), .C(
        \u_decoder/fir_filter/Q_data_mult_0 [0]), .D(
        \u_decoder/iq_demod/state [1]), .Q(\u_decoder/iq_demod/n50 ) );
  XOR21 U1996 ( .A(\u_decoder/iq_demod/dp_cluster_1/mult_I_sin_out [0]), .B(
        \u_decoder/iq_demod/dp_cluster_1/mult_Q_cos_out [0]), .Q(
        \u_decoder/iq_demod/add_Q_out [0]) );
  INV3 U1997 ( .A(\u_decoder/iq_demod/n41 ), .Q(n2274) );
  AOI221 U1998 ( .A(\u_decoder/iq_demod/add_I_out [0]), .B(n779), .C(
        \u_decoder/iq_demod/state [1]), .D(
        \u_decoder/fir_filter/I_data_mult_0 [0]), .Q(\u_decoder/iq_demod/n41 )
         );
  XNR21 U1999 ( .A(\u_decoder/iq_demod/dp_cluster_0/mult_I_cos_out [0]), .B(
        n2383), .Q(\u_decoder/iq_demod/add_I_out [0]) );
  INV3 U2000 ( .A(\u_inFIFO/n529 ), .Q(n1814) );
  AOI221 U2001 ( .A(n912), .B(n1199), .C(\u_inFIFO/n523 ), .D(n198), .Q(
        \u_inFIFO/n529 ) );
  INV3 U2002 ( .A(\u_cordic/mycordic/n381 ), .Q(n1470) );
  AOI221 U2003 ( .A(\u_cordic/mycordic/N317 ), .B(\u_cordic/mycordic/n336 ), 
        .C(\u_cordic/mycordic/N349 ), .D(n1904), .Q(\u_cordic/mycordic/n381 )
         );
  INV3 U2004 ( .A(\u_cordic/mycordic/n373 ), .Q(n1563) );
  AOI221 U2005 ( .A(\u_cordic/mycordic/N381 ), .B(n778), .C(
        \u_cordic/mycordic/N413 ), .D(n1908), .Q(\u_cordic/mycordic/n373 ) );
  INV3 U2006 ( .A(\u_cordic/mycordic/n536 ), .Q(n1485) );
  NOR21 U2007 ( .A(n773), .B(n1905), .Q(\u_cordic/mycordic/n536 ) );
  INV3 U2008 ( .A(\u_decoder/iq_demod/n70 ), .Q(n1909) );
  NAND22 U2009 ( .A(\u_decoder/iq_demod/n71 ), .B(n1212), .Q(
        \u_decoder/iq_demod/n70 ) );
  INV3 U2010 ( .A(n779), .Q(n2398) );
  NOR21 U2011 ( .A(n1237), .B(n1910), .Q(\u_decoder/iq_demod/n61 ) );
  INV3 U2012 ( .A(n1232), .Q(n1219) );
  INV3 U2013 ( .A(n1235), .Q(n1220) );
  INV3 U2014 ( .A(n1235), .Q(n1224) );
  INV3 U2015 ( .A(n1234), .Q(n1223) );
  INV3 U2016 ( .A(n1232), .Q(n1221) );
  INV3 U2017 ( .A(n1232), .Q(n1222) );
  INV3 U2018 ( .A(n1233), .Q(n1230) );
  INV3 U2019 ( .A(n1238), .Q(n1229) );
  INV3 U2020 ( .A(n1236), .Q(n1227) );
  INV3 U2021 ( .A(n1239), .Q(n1228) );
  INV3 U2022 ( .A(n1236), .Q(n1226) );
  INV3 U2023 ( .A(n1233), .Q(n1225) );
  INV3 U2024 ( .A(n1235), .Q(n1212) );
  INV3 U2025 ( .A(n1233), .Q(n1216) );
  INV3 U2026 ( .A(n1235), .Q(n1213) );
  INV3 U2027 ( .A(n1234), .Q(n1214) );
  INV3 U2028 ( .A(n1234), .Q(n1215) );
  INV3 U2029 ( .A(n1234), .Q(n1231) );
  INV3 U2030 ( .A(n1232), .Q(n1218) );
  INV3 U2031 ( .A(n1233), .Q(n1217) );
  NAND22 U2032 ( .A(n1219), .B(sig_DEMUX_outDEMUX1[0]), .Q(
        \u_decoder/iq_demod/n69 ) );
  NOR21 U2033 ( .A(n2118), .B(n2140), .Q(sig_DEMUX_outDEMUX18[7]) );
  NOR21 U2034 ( .A(n2120), .B(n2140), .Q(sig_DEMUX_outDEMUX18[6]) );
  NOR21 U2035 ( .A(n2122), .B(n2140), .Q(sig_DEMUX_outDEMUX18[5]) );
  NOR21 U2036 ( .A(n2124), .B(n2140), .Q(sig_DEMUX_outDEMUX18[4]) );
  NOR21 U2037 ( .A(n2110), .B(n2140), .Q(sig_DEMUX_outDEMUX17[7]) );
  NOR21 U2038 ( .A(n2112), .B(n2140), .Q(sig_DEMUX_outDEMUX17[6]) );
  NOR21 U2039 ( .A(n2114), .B(n2140), .Q(sig_DEMUX_outDEMUX17[5]) );
  NOR21 U2040 ( .A(n2116), .B(n2140), .Q(sig_DEMUX_outDEMUX17[4]) );
  BUF2 U2041 ( .A(n1958), .Q(n1082) );
  BUF2 U2042 ( .A(n1957), .Q(n1066) );
  BUF2 U2043 ( .A(n1956), .Q(n1050) );
  BUF2 U2044 ( .A(n1955), .Q(n1034) );
  BUF2 U2045 ( .A(n1958), .Q(n1081) );
  BUF2 U2046 ( .A(n1957), .Q(n1065) );
  BUF2 U2047 ( .A(n1956), .Q(n1049) );
  BUF2 U2048 ( .A(n1955), .Q(n1033) );
  BUF2 U2049 ( .A(n1958), .Q(n1080) );
  BUF2 U2050 ( .A(n1957), .Q(n1064) );
  BUF2 U2051 ( .A(n1956), .Q(n1048) );
  BUF2 U2052 ( .A(n1955), .Q(n1032) );
  BUF2 U2053 ( .A(n1958), .Q(n1079) );
  BUF2 U2054 ( .A(n1957), .Q(n1063) );
  BUF2 U2055 ( .A(n1956), .Q(n1047) );
  BUF2 U2056 ( .A(n1955), .Q(n1031) );
  BUF2 U2057 ( .A(n1958), .Q(n1078) );
  BUF2 U2058 ( .A(n1957), .Q(n1062) );
  BUF2 U2059 ( .A(n1956), .Q(n1046) );
  BUF2 U2060 ( .A(n1955), .Q(n1030) );
  BUF2 U2061 ( .A(n1958), .Q(n1077) );
  BUF2 U2062 ( .A(n1957), .Q(n1061) );
  BUF2 U2063 ( .A(n1956), .Q(n1045) );
  BUF2 U2064 ( .A(n1955), .Q(n1029) );
  BUF2 U2065 ( .A(n1958), .Q(n1076) );
  BUF2 U2066 ( .A(n1957), .Q(n1060) );
  BUF2 U2067 ( .A(n1956), .Q(n1044) );
  BUF2 U2068 ( .A(n1955), .Q(n1028) );
  BUF2 U2069 ( .A(n1958), .Q(n1075) );
  BUF2 U2070 ( .A(n1957), .Q(n1059) );
  BUF2 U2071 ( .A(n1956), .Q(n1043) );
  BUF2 U2072 ( .A(n1955), .Q(n1027) );
  BUF2 U2073 ( .A(n1958), .Q(n1074) );
  BUF2 U2074 ( .A(n1957), .Q(n1058) );
  BUF2 U2075 ( .A(n1956), .Q(n1042) );
  BUF2 U2076 ( .A(n1955), .Q(n1026) );
  BUF2 U2077 ( .A(n1958), .Q(n1073) );
  BUF2 U2078 ( .A(n1957), .Q(n1057) );
  BUF2 U2079 ( .A(n1956), .Q(n1041) );
  BUF2 U2080 ( .A(n1955), .Q(n1025) );
  BUF2 U2081 ( .A(n1958), .Q(n1072) );
  BUF2 U2082 ( .A(n1957), .Q(n1056) );
  BUF2 U2083 ( .A(n1956), .Q(n1040) );
  BUF2 U2084 ( .A(n1955), .Q(n1024) );
  BUF2 U2085 ( .A(n1958), .Q(n1071) );
  BUF2 U2086 ( .A(n1957), .Q(n1055) );
  BUF2 U2087 ( .A(n1956), .Q(n1039) );
  BUF2 U2088 ( .A(n1955), .Q(n1023) );
  BUF2 U2089 ( .A(n1958), .Q(n1070) );
  BUF2 U2090 ( .A(n1957), .Q(n1054) );
  BUF2 U2091 ( .A(n1956), .Q(n1038) );
  BUF2 U2092 ( .A(n1955), .Q(n1022) );
  BUF2 U2093 ( .A(n1958), .Q(n1069) );
  BUF2 U2094 ( .A(n1957), .Q(n1053) );
  BUF2 U2095 ( .A(n1956), .Q(n1037) );
  BUF2 U2096 ( .A(n1955), .Q(n1021) );
  BUF2 U2097 ( .A(n1958), .Q(n1068) );
  BUF2 U2098 ( .A(n1957), .Q(n1052) );
  BUF2 U2099 ( .A(n1956), .Q(n1036) );
  BUF2 U2100 ( .A(n1955), .Q(n1020) );
  BUF2 U2101 ( .A(n1958), .Q(n1067) );
  BUF2 U2102 ( .A(n1957), .Q(n1051) );
  BUF2 U2103 ( .A(n1956), .Q(n1035) );
  BUF2 U2104 ( .A(n1955), .Q(n1019) );
  NAND41 U2105 ( .A(n1389), .B(n1388), .C(n1387), .D(n1386), .Q(n1392) );
  NOR40 U2106 ( .A(n1385), .B(n1384), .C(n1383), .D(n1382), .Q(n1386) );
  NAND41 U2107 ( .A(n1376), .B(n1388), .C(n1375), .D(n1374), .Q(n2675) );
  NOR40 U2108 ( .A(n1373), .B(n1372), .C(n1371), .D(n1370), .Q(n1374) );
  NOR40 U2109 ( .A(n1358), .B(n1357), .C(n1356), .D(n1355), .Q(n1359) );
  NAND41 U2110 ( .A(n3046), .B(n3045), .C(n3044), .D(n3043), .Q(n3051) );
  XNR21 U2111 ( .A(\u_cdr/phd1/cnt_phd/N12 ), .B(\u_cdr/phd1/cnt_phd/cnt [2]), 
        .Q(n3044) );
  XNR21 U2112 ( .A(\u_cdr/phd1/cnt_phd/N13 ), .B(\u_cdr/phd1/cnt_phd/cnt [3]), 
        .Q(n3045) );
  XNR21 U2113 ( .A(n2678), .B(\u_cdr/phd1/cnt_phd/cnt [5]), .Q(n3043) );
  NAND41 U2114 ( .A(n1361), .B(n1388), .C(n1360), .D(n1359), .Q(n1362) );
  NAND41 U2115 ( .A(n61), .B(n1388), .C(n1320), .D(n1300), .Q(n1301) );
  NOR40 U2116 ( .A(n1299), .B(n1298), .C(n1297), .D(n1296), .Q(n1300) );
  XNR21 U2117 ( .A(\u_cdr/phd1/cnt_phd/N14 ), .B(\u_cdr/phd1/cnt_phd/cnt [4]), 
        .Q(n3046) );
  AOI221 U2118 ( .A(\u_cdr/dec1/cnt_r [0]), .B(n1395), .C(n248), .D(n1394), 
        .Q(\u_cdr/dec1/n33 ) );
  AOI221 U2119 ( .A(\u_cdr/dec1/cnt_r [5]), .B(n1395), .C(\u_cdr/dec1/N65 ), 
        .D(n1394), .Q(\u_cdr/dec1/n32 ) );
  XOR21 U2120 ( .A(\u_cdr/dec1/add_40/carry [5]), .B(\u_cdr/dec1/cnt_r [5]), 
        .Q(\u_cdr/dec1/N65 ) );
  AOI221 U2121 ( .A(\u_cdr/dec1/cnt_r [4]), .B(n1395), .C(\u_cdr/dec1/N64 ), 
        .D(n1394), .Q(\u_cdr/dec1/n26 ) );
  AOI221 U2122 ( .A(\u_cdr/dec1/cnt_r [3]), .B(n1395), .C(\u_cdr/dec1/N63 ), 
        .D(n1394), .Q(\u_cdr/dec1/n29 ) );
  AOI221 U2123 ( .A(\u_cdr/dec1/cnt_r [2]), .B(n1395), .C(\u_cdr/dec1/N62 ), 
        .D(n1394), .Q(\u_cdr/dec1/n30 ) );
  AOI221 U2124 ( .A(\u_cdr/dec1/cnt_r [1]), .B(n1395), .C(\u_cdr/dec1/N61 ), 
        .D(n1394), .Q(\u_cdr/dec1/n31 ) );
  INV3 U2125 ( .A(\u_cdr/div1/cnt_div/n40 ), .Q(n1414) );
  AOI221 U2126 ( .A(\u_cdr/div1/cnt_div/n34 ), .B(n262), .C(
        \u_cdr/div1/cnt_div/n35 ), .D(\u_cdr/div1/cnt_div/cnt [0]), .Q(
        \u_cdr/div1/cnt_div/n40 ) );
  INV3 U2127 ( .A(\u_cdr/div1/cnt_div/n39 ), .Q(n1415) );
  AOI221 U2128 ( .A(\u_cdr/div1/cnt_div/n34 ), .B(\u_cdr/div1/cnt_div/N76 ), 
        .C(\u_cdr/div1/cnt_div/n35 ), .D(\u_cdr/div1/cnt_div/cnt [5]), .Q(
        \u_cdr/div1/cnt_div/n39 ) );
  XOR21 U2129 ( .A(\u_cdr/div1/cnt_div/add_58/carry [5]), .B(
        \u_cdr/div1/cnt_div/cnt [5]), .Q(\u_cdr/div1/cnt_div/N76 ) );
  INV3 U2130 ( .A(\u_cdr/div1/cnt_div/n33 ), .Q(n1419) );
  AOI221 U2131 ( .A(\u_cdr/div1/cnt_div/n34 ), .B(\u_cdr/div1/cnt_div/N75 ), 
        .C(\u_cdr/div1/cnt_div/n35 ), .D(\u_cdr/div1/cnt_div/cnt [4]), .Q(
        \u_cdr/div1/cnt_div/n33 ) );
  INV3 U2132 ( .A(\u_cdr/div1/cnt_div/n36 ), .Q(n1418) );
  AOI221 U2133 ( .A(\u_cdr/div1/cnt_div/n34 ), .B(\u_cdr/div1/cnt_div/N74 ), 
        .C(\u_cdr/div1/cnt_div/n35 ), .D(\u_cdr/div1/cnt_div/cnt [3]), .Q(
        \u_cdr/div1/cnt_div/n36 ) );
  INV3 U2134 ( .A(\u_cdr/div1/cnt_div/n37 ), .Q(n1417) );
  AOI221 U2135 ( .A(\u_cdr/div1/cnt_div/n34 ), .B(\u_cdr/div1/cnt_div/N73 ), 
        .C(\u_cdr/div1/cnt_div/n35 ), .D(\u_cdr/div1/cnt_div/cnt [2]), .Q(
        \u_cdr/div1/cnt_div/n37 ) );
  INV3 U2136 ( .A(\u_cdr/div1/cnt_div/n38 ), .Q(n1416) );
  AOI221 U2137 ( .A(\u_cdr/div1/cnt_div/n34 ), .B(\u_cdr/div1/cnt_div/N72 ), 
        .C(\u_cdr/div1/cnt_div/n35 ), .D(\u_cdr/div1/cnt_div/cnt [1]), .Q(
        \u_cdr/div1/cnt_div/n38 ) );
  INV3 U2138 ( .A(n3063), .Q(n1402) );
  AOI221 U2139 ( .A(n3057), .B(n3055), .C(n3058), .D(
        \u_cdr/phd1/cnt_phd/cnt [0]), .Q(n3063) );
  INV3 U2140 ( .A(n3062), .Q(n1403) );
  AOI221 U2141 ( .A(n3057), .B(\u_cdr/phd1/cnt_phd/N76 ), .C(n3058), .D(
        \u_cdr/phd1/cnt_phd/cnt [5]), .Q(n3062) );
  XOR21 U2142 ( .A(\u_cdr/phd1/cnt_phd/add_58/carry [5]), .B(
        \u_cdr/phd1/cnt_phd/cnt [5]), .Q(\u_cdr/phd1/cnt_phd/N76 ) );
  INV3 U2143 ( .A(n3056), .Q(n1407) );
  AOI221 U2144 ( .A(n3057), .B(\u_cdr/phd1/cnt_phd/N75 ), .C(n3058), .D(
        \u_cdr/phd1/cnt_phd/cnt [4]), .Q(n3056) );
  INV3 U2145 ( .A(n3059), .Q(n1406) );
  AOI221 U2146 ( .A(n3057), .B(\u_cdr/phd1/cnt_phd/N74 ), .C(n3058), .D(
        \u_cdr/phd1/cnt_phd/cnt [3]), .Q(n3059) );
  INV3 U2147 ( .A(n3060), .Q(n1405) );
  AOI221 U2148 ( .A(n3057), .B(\u_cdr/phd1/cnt_phd/N73 ), .C(n3058), .D(
        \u_cdr/phd1/cnt_phd/cnt [2]), .Q(n3060) );
  INV3 U2149 ( .A(n3061), .Q(n1404) );
  AOI221 U2150 ( .A(n3057), .B(\u_cdr/phd1/cnt_phd/N72 ), .C(n3058), .D(
        \u_cdr/phd1/cnt_phd/cnt [1]), .Q(n3061) );
  INV3 U2151 ( .A(\u_cdr/dec1/cnt_dec/n23 ), .Q(n1408) );
  AOI221 U2152 ( .A(\u_cdr/dec1/cnt_dec/cnt_dec [0]), .B(
        \u_cdr/dec1/cnt_dec/n17 ), .C(n263), .D(\u_cdr/dec1/cnt_dec/n18 ), .Q(
        \u_cdr/dec1/cnt_dec/n23 ) );
  INV3 U2153 ( .A(\u_cdr/dec1/cnt_dec/n22 ), .Q(n1409) );
  AOI221 U2154 ( .A(\u_cdr/dec1/cnt_dec/cnt_dec [1]), .B(
        \u_cdr/dec1/cnt_dec/n17 ), .C(\u_cdr/dec1/cnt_dec/N5 ), .D(
        \u_cdr/dec1/cnt_dec/n18 ), .Q(\u_cdr/dec1/cnt_dec/n22 ) );
  INV3 U2155 ( .A(\u_cdr/dec1/cnt_dec/n21 ), .Q(n1410) );
  AOI221 U2156 ( .A(\u_cdr/dec1/cnt_dec/cnt_dec [2]), .B(
        \u_cdr/dec1/cnt_dec/n17 ), .C(\u_cdr/dec1/cnt_dec/N6 ), .D(
        \u_cdr/dec1/cnt_dec/n18 ), .Q(\u_cdr/dec1/cnt_dec/n21 ) );
  INV3 U2157 ( .A(\u_cdr/dec1/cnt_dec/n20 ), .Q(n1411) );
  AOI221 U2158 ( .A(\u_cdr/dec1/cnt_dec/cnt_dec [3]), .B(
        \u_cdr/dec1/cnt_dec/n17 ), .C(\u_cdr/dec1/cnt_dec/N7 ), .D(
        \u_cdr/dec1/cnt_dec/n18 ), .Q(\u_cdr/dec1/cnt_dec/n20 ) );
  INV3 U2159 ( .A(\u_cdr/dec1/cnt_dec/n19 ), .Q(n1412) );
  AOI221 U2160 ( .A(\u_cdr/dec1/cnt_dec/cnt_dec [4]), .B(
        \u_cdr/dec1/cnt_dec/n17 ), .C(\u_cdr/dec1/cnt_dec/N8 ), .D(
        \u_cdr/dec1/cnt_dec/n18 ), .Q(\u_cdr/dec1/cnt_dec/n19 ) );
  INV3 U2161 ( .A(\u_cdr/dec1/cnt_dec/n16 ), .Q(n1413) );
  AOI221 U2162 ( .A(\u_cdr/dec1/cnt_dec/cnt_dec [5]), .B(
        \u_cdr/dec1/cnt_dec/n17 ), .C(\u_cdr/dec1/cnt_dec/N9 ), .D(
        \u_cdr/dec1/cnt_dec/n18 ), .Q(\u_cdr/dec1/cnt_dec/n16 ) );
  XOR21 U2163 ( .A(\u_cdr/dec1/cnt_dec/add_20/carry [5]), .B(
        \u_cdr/dec1/cnt_dec/cnt_dec [5]), .Q(\u_cdr/dec1/cnt_dec/N9 ) );
  NOR40 U2164 ( .A(n1367), .B(n1366), .C(n1365), .D(n1364), .Q(n1368) );
  NAND41 U2165 ( .A(n1343), .B(n1342), .C(n1388), .D(n1341), .Q(n1353) );
  NOR31 U2166 ( .A(n1391), .B(n1240), .C(n316), .Q(n1341) );
  NOR40 U2167 ( .A(n1353), .B(n1352), .C(n1351), .D(n1350), .Q(
        \u_cdr/dec1/N73 ) );
  NOR21 U2168 ( .A(n2676), .B(n1237), .Q(\u_cdr/dec1/cnt_dec/N33 ) );
  NAND41 U2169 ( .A(n1369), .B(n1388), .C(n315), .D(n1368), .Q(n2676) );
  INV3 U2170 ( .A(n3048), .Q(n2679) );
  AOI221 U2171 ( .A(n293), .B(n3047), .C(n3047), .D(n1400), .Q(n3048) );
  INV3 U2172 ( .A(n3065), .Q(n1834) );
  NAND22 U2173 ( .A(\u_cdr/phd1/cnt_phd/N58 ), .B(n1217), .Q(n3065) );
  NOR40 U2174 ( .A(n61), .B(n1319), .C(n1318), .D(n1317), .Q(
        \u_cdr/phd1/cnt_phd/N58 ) );
  AOI311 U2175 ( .A(\u_cdr/div1/w_en_freq_synch ), .B(\u_cdr/w_sT ), .C(
        \u_cdr/div1/n32 ), .D(n1239), .Q(n1244) );
  NAND31 U2176 ( .A(n1251), .B(n1274), .C(n1250), .Q(\u_cdr/div1/n36 ) );
  IMUX21 U2177 ( .A(n1249), .B(n1248), .S(\u_cdr/w_nb_P [3]), .Q(n1250) );
  NOR31 U2178 ( .A(n1271), .B(n221), .C(n1313), .Q(n1249) );
  OAI311 U2179 ( .A(n1272), .B(n1271), .C(\u_cdr/w_sE ), .D(\u_cdr/div1/N35 ), 
        .Q(n1273) );
  IMUX21 U2180 ( .A(n1255), .B(n1254), .S(\u_cdr/w_nb_P [4]), .Q(n1256) );
  OAI311 U2181 ( .A(n1271), .B(n221), .C(n1265), .D(n1251), .Q(n1255) );
  INV3 U2182 ( .A(n3066), .Q(n1835) );
  NAND22 U2183 ( .A(\u_cdr/phd1/cnt_phd/N50 ), .B(n1217), .Q(n3066) );
  NOR40 U2184 ( .A(n1335), .B(n1334), .C(n1333), .D(n1332), .Q(
        \u_cdr/phd1/cnt_phd/N50 ) );
  NAND41 U2185 ( .A(n1212), .B(\u_cdr/div1/w_en_freq_synch ), .C(\u_cdr/w_sT ), 
        .D(\u_cdr/div1/n32 ), .Q(\u_cdr/div1/n31 ) );
  NAND31 U2186 ( .A(\u_cdr/div1/w_en_freq_synch ), .B(\u_cdr/w_sT ), .C(n1217), 
        .Q(\u_cdr/div1/n27 ) );
  NAND22 U2187 ( .A(n1218), .B(n62), .Q(\u_cdr/phd1/n21 ) );
  AOI221 U2188 ( .A(n1279), .B(n1269), .C(n1278), .D(n1268), .Q(n1270) );
  IMUX21 U2189 ( .A(n1279), .B(n1278), .S(n1277), .Q(n1280) );
  NOR21 U2190 ( .A(n1284), .B(n1276), .Q(n1277) );
  NAND22 U2191 ( .A(\u_cdr/w_sE ), .B(n1850), .Q(\u_cdr/phd1/n20 ) );
  XNR21 U2192 ( .A(\u_cdr/phd1/w_s4 ), .B(\u_cdr/phd1/w_s2 ), .Q(
        \u_cdr/phd1/n19 ) );
  NAND22 U2193 ( .A(\u_cdr/w_sT ), .B(n1850), .Q(\u_cdr/phd1/n18 ) );
  XNR21 U2194 ( .A(\u_cdr/phd1/w_s2 ), .B(\u_cdr/phd1/w_s1 ), .Q(
        \u_cdr/phd1/n16 ) );
  NOR40 U2195 ( .A(n2673), .B(n2672), .C(n2671), .D(n2670), .Q(
        \u_cordic/my_rotation/n55 ) );
  INV3 U2196 ( .A(\u_cordic/my_rotation/n70 ), .Q(n2670) );
  AOI221 U2197 ( .A(\u_cordic/my_rotation/N25 ), .B(n2674), .C(
        \u_cordic/my_rotation/N25 ), .D(n767), .Q(\u_cordic/my_rotation/n70 )
         );
  XNR21 U2198 ( .A(\u_cordic/my_rotation/present_angle[0][0] ), .B(n65), .Q(
        \u_cordic/my_rotation/N25 ) );
  NOR40 U2199 ( .A(\u_cordic/my_rotation/n59 ), .B(n2662), .C(\u_cordic/dir ), 
        .D(n2661), .Q(\u_cordic/my_rotation/n58 ) );
  NAND22 U2200 ( .A(\u_cordic/my_rotation/n48 ), .B(\u_cordic/my_rotation/n47 ), .Q(\u_cordic/my_rotation/n59 ) );
  BUF2 U2201 ( .A(\u_coder/j [1]), .Q(n762) );
  BUF2 U2202 ( .A(\u_coder/i [0]), .Q(n763) );
  INV3 U2203 ( .A(n394), .Q(\u_cordic/my_rotation/sub_35/carry [1]) );
  NOR21 U2204 ( .A(n65), .B(\u_cordic/my_rotation/present_angle[0][0] ), .Q(
        n394) );
  INV3 U2205 ( .A(\u_coder/n282 ), .Q(n1915) );
  AOI221 U2206 ( .A(n890), .B(\u_coder/j [19]), .C(n2169), .D(\u_coder/N1032 ), 
        .Q(\u_coder/n282 ) );
  XOR21 U2207 ( .A(\u_coder/add_282/carry [19]), .B(\u_coder/j [19]), .Q(
        \u_coder/N1032 ) );
  INV3 U2208 ( .A(\u_coder/n304 ), .Q(n1935) );
  AOI221 U2209 ( .A(n894), .B(\u_coder/i [19]), .C(n2156), .D(\u_coder/N726 ), 
        .Q(\u_coder/n304 ) );
  XOR21 U2210 ( .A(\u_coder/add_206/carry [19]), .B(\u_coder/i [19]), .Q(
        \u_coder/N726 ) );
  XNR21 U2211 ( .A(\u_coder/add_93/carry [19]), .B(\u_coder/c [19]), .Q(n373)
         );
  INV3 U2212 ( .A(\u_coder/n262 ), .Q(n1934) );
  AOI221 U2213 ( .A(\u_coder/n263 ), .B(\u_coder/j [18]), .C(n2169), .D(
        \u_coder/N1031 ), .Q(\u_coder/n262 ) );
  INV3 U2214 ( .A(\u_coder/n284 ), .Q(n1954) );
  AOI221 U2215 ( .A(n894), .B(\u_coder/i [18]), .C(n2156), .D(\u_coder/N725 ), 
        .Q(\u_coder/n284 ) );
  INV3 U2216 ( .A(\u_coder/n264 ), .Q(n1933) );
  AOI221 U2217 ( .A(n890), .B(\u_coder/j [17]), .C(n2169), .D(\u_coder/N1030 ), 
        .Q(\u_coder/n264 ) );
  INV3 U2218 ( .A(\u_coder/n286 ), .Q(n1953) );
  AOI221 U2219 ( .A(n894), .B(\u_coder/i [17]), .C(n2156), .D(\u_coder/N724 ), 
        .Q(\u_coder/n286 ) );
  INV3 U2220 ( .A(\u_coder/n265 ), .Q(n1932) );
  AOI221 U2221 ( .A(\u_coder/n263 ), .B(\u_coder/j [16]), .C(n2169), .D(
        \u_coder/N1029 ), .Q(\u_coder/n265 ) );
  INV3 U2222 ( .A(\u_coder/n287 ), .Q(n1952) );
  AOI221 U2223 ( .A(n893), .B(\u_coder/i [16]), .C(n2156), .D(\u_coder/N723 ), 
        .Q(\u_coder/n287 ) );
  INV3 U2224 ( .A(n2985), .Q(n2544) );
  INV3 U2225 ( .A(n2966), .Q(n2424) );
  INV3 U2226 ( .A(n2987), .Q(n2542) );
  INV3 U2227 ( .A(n2968), .Q(n2422) );
  INV3 U2228 ( .A(n2989), .Q(n2540) );
  INV3 U2229 ( .A(n2970), .Q(n2420) );
  INV3 U2230 ( .A(n2991), .Q(n2538) );
  INV3 U2231 ( .A(n2972), .Q(n2418) );
  OAI2111 U2232 ( .A(\u_decoder/fir_filter/I_data_mult_0_buff [1]), .B(
        \u_decoder/fir_filter/I_data_add_1_buff [1]), .C(
        \u_decoder/fir_filter/I_data_mult_0_buff [0]), .D(
        \u_decoder/fir_filter/I_data_add_1_buff [0]), .Q(n2984) );
  OAI2111 U2233 ( .A(\u_decoder/fir_filter/Q_data_mult_0_buff [1]), .B(
        \u_decoder/fir_filter/Q_data_add_1_buff [1]), .C(
        \u_decoder/fir_filter/Q_data_mult_0_buff [0]), .D(
        \u_decoder/fir_filter/Q_data_add_1_buff [0]), .Q(n2965) );
  AOI211 U2234 ( .A(n3000), .B(\u_decoder/fir_filter/I_data_mult_0_buff [9]), 
        .C(n2529), .Q(n3002) );
  INV3 U2235 ( .A(n2999), .Q(n2529) );
  AOI211 U2236 ( .A(n2981), .B(\u_decoder/fir_filter/Q_data_mult_0_buff [9]), 
        .C(n2409), .Q(n2983) );
  INV3 U2237 ( .A(n2980), .Q(n2409) );
  AOI211 U2238 ( .A(n2996), .B(\u_decoder/fir_filter/I_data_mult_0_buff [7]), 
        .C(n2533), .Q(n2998) );
  INV3 U2239 ( .A(n2995), .Q(n2533) );
  AOI211 U2240 ( .A(n2977), .B(\u_decoder/fir_filter/Q_data_mult_0_buff [7]), 
        .C(n2413), .Q(n2979) );
  INV3 U2241 ( .A(n2976), .Q(n2413) );
  INV3 U2242 ( .A(\u_coder/n267 ), .Q(n1930) );
  AOI221 U2243 ( .A(n890), .B(\u_coder/j [14]), .C(n2169), .D(\u_coder/N1027 ), 
        .Q(\u_coder/n267 ) );
  INV3 U2244 ( .A(\u_coder/n289 ), .Q(n1950) );
  AOI221 U2245 ( .A(n893), .B(\u_coder/i [14]), .C(n2156), .D(\u_coder/N721 ), 
        .Q(\u_coder/n289 ) );
  INV3 U2246 ( .A(\u_coder/n266 ), .Q(n1931) );
  AOI221 U2247 ( .A(\u_coder/n263 ), .B(\u_coder/j [15]), .C(n2169), .D(
        \u_coder/N1028 ), .Q(\u_coder/n266 ) );
  INV3 U2248 ( .A(\u_coder/n288 ), .Q(n1951) );
  AOI221 U2249 ( .A(n893), .B(\u_coder/i [15]), .C(n2156), .D(\u_coder/N722 ), 
        .Q(\u_coder/n288 ) );
  INV3 U2250 ( .A(\u_decoder/fir_filter/n622 ), .Q(n2458) );
  AOI221 U2251 ( .A(\u_decoder/fir_filter/Q_data_add_4 [13]), .B(n1087), .C(
        \u_decoder/fir_filter/Q_data_add_4_buff [13]), .D(n1162), .Q(
        \u_decoder/fir_filter/n622 ) );
  INV3 U2252 ( .A(\u_decoder/fir_filter/n920 ), .Q(n2578) );
  AOI221 U2253 ( .A(\u_decoder/fir_filter/I_data_add_4 [13]), .B(n1095), .C(
        \u_decoder/fir_filter/I_data_add_4_buff [13]), .D(n1153), .Q(
        \u_decoder/fir_filter/n920 ) );
  INV3 U2254 ( .A(\u_decoder/fir_filter/n1083 ), .Q(n2258) );
  AOI221 U2255 ( .A(\u_decoder/fir_filter/I_data_mult_4 [13]), .B(n1094), .C(
        \u_decoder/fir_filter/I_data_mult_4_buff [13]), .D(n1162), .Q(
        \u_decoder/fir_filter/n1083 ) );
  INV3 U2256 ( .A(\u_decoder/fir_filter/n786 ), .Q(n2329) );
  AOI221 U2257 ( .A(\u_decoder/fir_filter/Q_data_mult_4 [13]), .B(n1083), .C(
        \u_decoder/fir_filter/Q_data_mult_4_buff [13]), .D(n1163), .Q(
        \u_decoder/fir_filter/n786 ) );
  INV3 U2258 ( .A(n2998), .Q(n2532) );
  INV3 U2259 ( .A(n2979), .Q(n2412) );
  NAND22 U2260 ( .A(\u_decoder/fir_filter/I_data_mult_1_buff [12]), .B(n1160), 
        .Q(\u_decoder/fir_filter/n1130 ) );
  NAND22 U2261 ( .A(\u_decoder/fir_filter/I_data_mult_2_buff [11]), .B(n1159), 
        .Q(\u_decoder/fir_filter/n1113 ) );
  NAND22 U2262 ( .A(\u_decoder/fir_filter/I_data_mult_3_buff [13]), .B(n1158), 
        .Q(\u_decoder/fir_filter/n1099 ) );
  NAND22 U2263 ( .A(\u_decoder/fir_filter/I_data_mult_5_buff [13]), .B(n1158), 
        .Q(\u_decoder/fir_filter/n1067 ) );
  NAND22 U2264 ( .A(\u_decoder/fir_filter/I_data_mult_6_buff [11]), .B(n1157), 
        .Q(\u_decoder/fir_filter/n1048 ) );
  NAND22 U2265 ( .A(\u_decoder/fir_filter/I_data_mult_7_buff [12]), .B(n1156), 
        .Q(\u_decoder/fir_filter/n1032 ) );
  NAND22 U2266 ( .A(\u_decoder/fir_filter/Q_data_mult_1_buff [12]), .B(n1152), 
        .Q(\u_decoder/fir_filter/n833 ) );
  NAND22 U2267 ( .A(\u_decoder/fir_filter/Q_data_mult_2_buff [11]), .B(n1159), 
        .Q(\u_decoder/fir_filter/n816 ) );
  NAND22 U2268 ( .A(\u_decoder/fir_filter/Q_data_mult_3_buff [13]), .B(n1153), 
        .Q(\u_decoder/fir_filter/n802 ) );
  NAND22 U2269 ( .A(\u_decoder/fir_filter/Q_data_mult_5_buff [13]), .B(n1154), 
        .Q(\u_decoder/fir_filter/n770 ) );
  NAND22 U2270 ( .A(\u_decoder/fir_filter/Q_data_mult_6_buff [11]), .B(n1155), 
        .Q(\u_decoder/fir_filter/n751 ) );
  NAND22 U2271 ( .A(\u_decoder/fir_filter/Q_data_mult_7_buff [12]), .B(n1154), 
        .Q(\u_decoder/fir_filter/n735 ) );
  NAND22 U2272 ( .A(\u_decoder/fir_filter/I_data_mult_0_buff [11]), .B(n1160), 
        .Q(\u_decoder/fir_filter/n1145 ) );
  NAND22 U2273 ( .A(\u_decoder/fir_filter/Q_data_mult_0_buff [11]), .B(n1151), 
        .Q(\u_decoder/fir_filter/n848 ) );
  NAND22 U2274 ( .A(\u_decoder/fir_filter/I_data_mult_3_buff [10]), .B(n1158), 
        .Q(\u_decoder/fir_filter/n1096 ) );
  NAND22 U2275 ( .A(\u_decoder/fir_filter/I_data_mult_5_buff [10]), .B(n1156), 
        .Q(\u_decoder/fir_filter/n1064 ) );
  NAND22 U2276 ( .A(\u_decoder/fir_filter/Q_data_mult_3_buff [10]), .B(n1156), 
        .Q(\u_decoder/fir_filter/n799 ) );
  NAND22 U2277 ( .A(\u_decoder/fir_filter/Q_data_mult_5_buff [10]), .B(n1154), 
        .Q(\u_decoder/fir_filter/n767 ) );
  NAND22 U2278 ( .A(\u_decoder/fir_filter/I_data_mult_2_buff [12]), .B(n1159), 
        .Q(\u_decoder/fir_filter/n1114 ) );
  NAND22 U2279 ( .A(\u_decoder/fir_filter/I_data_mult_3_buff [14]), .B(n1158), 
        .Q(\u_decoder/fir_filter/n1100 ) );
  NAND22 U2280 ( .A(\u_decoder/fir_filter/I_data_mult_3_buff [12]), .B(n1158), 
        .Q(\u_decoder/fir_filter/n1098 ) );
  NAND22 U2281 ( .A(\u_decoder/fir_filter/I_data_mult_5_buff [14]), .B(n1151), 
        .Q(\u_decoder/fir_filter/n1068 ) );
  NAND22 U2282 ( .A(\u_decoder/fir_filter/I_data_mult_5_buff [12]), .B(n1157), 
        .Q(\u_decoder/fir_filter/n1066 ) );
  NAND22 U2283 ( .A(\u_decoder/fir_filter/I_data_mult_6_buff [12]), .B(n1157), 
        .Q(\u_decoder/fir_filter/n1049 ) );
  NAND22 U2284 ( .A(\u_decoder/fir_filter/Q_data_mult_2_buff [12]), .B(n1160), 
        .Q(\u_decoder/fir_filter/n817 ) );
  NAND22 U2285 ( .A(\u_decoder/fir_filter/Q_data_mult_3_buff [14]), .B(n1155), 
        .Q(\u_decoder/fir_filter/n803 ) );
  NAND22 U2286 ( .A(\u_decoder/fir_filter/Q_data_mult_3_buff [12]), .B(n1154), 
        .Q(\u_decoder/fir_filter/n801 ) );
  NAND22 U2287 ( .A(\u_decoder/fir_filter/Q_data_mult_5_buff [14]), .B(n1154), 
        .Q(\u_decoder/fir_filter/n771 ) );
  NAND22 U2288 ( .A(\u_decoder/fir_filter/Q_data_mult_5_buff [12]), .B(n1154), 
        .Q(\u_decoder/fir_filter/n769 ) );
  NAND22 U2289 ( .A(\u_decoder/fir_filter/Q_data_mult_6_buff [12]), .B(n1155), 
        .Q(\u_decoder/fir_filter/n752 ) );
  NAND22 U2290 ( .A(\u_decoder/fir_filter/I_data_mult_3_buff [11]), .B(n1158), 
        .Q(\u_decoder/fir_filter/n1097 ) );
  NAND22 U2291 ( .A(\u_decoder/fir_filter/I_data_mult_5_buff [11]), .B(n1155), 
        .Q(\u_decoder/fir_filter/n1065 ) );
  NAND22 U2292 ( .A(\u_decoder/fir_filter/Q_data_mult_3_buff [11]), .B(n1153), 
        .Q(\u_decoder/fir_filter/n800 ) );
  NAND22 U2293 ( .A(\u_decoder/fir_filter/Q_data_mult_5_buff [11]), .B(n1154), 
        .Q(\u_decoder/fir_filter/n768 ) );
  INV3 U2294 ( .A(\u_decoder/fir_filter/n919 ), .Q(n2577) );
  AOI221 U2295 ( .A(\u_decoder/fir_filter/I_data_add_4 [14]), .B(n1095), .C(
        \u_decoder/fir_filter/I_data_add_4_buff [14]), .D(n1161), .Q(
        \u_decoder/fir_filter/n919 ) );
  INV3 U2296 ( .A(\u_decoder/fir_filter/n621 ), .Q(n2457) );
  AOI221 U2297 ( .A(\u_decoder/fir_filter/Q_data_add_4 [14]), .B(n1087), .C(
        \u_decoder/fir_filter/Q_data_add_4_buff [14]), .D(n1162), .Q(
        \u_decoder/fir_filter/n621 ) );
  NOR21 U2298 ( .A(n106), .B(n26), .Q(\u_decoder/fir_filter/add_301/carry [1])
         );
  NOR21 U2299 ( .A(n108), .B(n27), .Q(\u_decoder/fir_filter/add_300/carry [1])
         );
  NOR21 U2300 ( .A(n109), .B(n28), .Q(\u_decoder/fir_filter/add_299/carry [1])
         );
  NOR21 U2301 ( .A(n110), .B(n29), .Q(\u_decoder/fir_filter/add_297/carry [1])
         );
  NOR21 U2302 ( .A(n111), .B(n30), .Q(\u_decoder/fir_filter/add_296/carry [1])
         );
  NOR21 U2303 ( .A(n112), .B(n31), .Q(\u_decoder/fir_filter/add_295/carry [1])
         );
  NOR21 U2304 ( .A(n107), .B(n32), .Q(\u_decoder/fir_filter/add_333/carry [1])
         );
  NOR21 U2305 ( .A(n113), .B(n33), .Q(\u_decoder/fir_filter/add_332/carry [1])
         );
  NOR21 U2306 ( .A(n114), .B(n34), .Q(\u_decoder/fir_filter/add_331/carry [1])
         );
  NOR21 U2307 ( .A(n115), .B(n35), .Q(\u_decoder/fir_filter/add_329/carry [1])
         );
  NOR21 U2308 ( .A(n116), .B(n36), .Q(\u_decoder/fir_filter/add_328/carry [1])
         );
  NOR21 U2309 ( .A(n117), .B(n37), .Q(\u_decoder/fir_filter/add_327/carry [1])
         );
  NOR21 U2310 ( .A(n118), .B(n38), .Q(\u_decoder/fir_filter/add_298/carry [1])
         );
  NOR21 U2311 ( .A(n119), .B(n39), .Q(\u_decoder/fir_filter/add_330/carry [1])
         );
  NAND22 U2312 ( .A(\u_decoder/fir_filter/n1019 ), .B(
        \u_decoder/fir_filter/n1148 ), .Q(\u_decoder/fir_filter/n1450 ) );
  NAND22 U2313 ( .A(\u_decoder/fir_filter/I_data_mult_0_buff [14]), .B(n1150), 
        .Q(\u_decoder/fir_filter/n1148 ) );
  NAND22 U2314 ( .A(\u_decoder/fir_filter/n1019 ), .B(
        \u_decoder/fir_filter/n1147 ), .Q(\u_decoder/fir_filter/n1449 ) );
  NAND22 U2315 ( .A(\u_decoder/fir_filter/I_data_mult_0_buff [13]), .B(n1156), 
        .Q(\u_decoder/fir_filter/n1147 ) );
  NAND22 U2316 ( .A(\u_decoder/fir_filter/n1019 ), .B(
        \u_decoder/fir_filter/n1146 ), .Q(\u_decoder/fir_filter/n1448 ) );
  NAND22 U2317 ( .A(\u_decoder/fir_filter/I_data_mult_0_buff [12]), .B(n1160), 
        .Q(\u_decoder/fir_filter/n1146 ) );
  NAND22 U2318 ( .A(\u_decoder/fir_filter/n1033 ), .B(
        \u_decoder/fir_filter/n1132 ), .Q(\u_decoder/fir_filter/n1434 ) );
  NAND22 U2319 ( .A(\u_decoder/fir_filter/I_data_mult_1_buff [14]), .B(n1160), 
        .Q(\u_decoder/fir_filter/n1132 ) );
  NAND22 U2320 ( .A(\u_decoder/fir_filter/n1033 ), .B(
        \u_decoder/fir_filter/n1131 ), .Q(\u_decoder/fir_filter/n1433 ) );
  NAND22 U2321 ( .A(\u_decoder/fir_filter/I_data_mult_1_buff [13]), .B(n1160), 
        .Q(\u_decoder/fir_filter/n1131 ) );
  NAND22 U2322 ( .A(\u_decoder/fir_filter/n1033 ), .B(
        \u_decoder/fir_filter/n1035 ), .Q(\u_decoder/fir_filter/n1354 ) );
  NAND22 U2323 ( .A(\u_decoder/fir_filter/I_data_mult_7_buff [14]), .B(n1156), 
        .Q(\u_decoder/fir_filter/n1035 ) );
  NAND22 U2324 ( .A(\u_decoder/fir_filter/n1033 ), .B(
        \u_decoder/fir_filter/n1034 ), .Q(\u_decoder/fir_filter/n1353 ) );
  NAND22 U2325 ( .A(\u_decoder/fir_filter/I_data_mult_7_buff [13]), .B(n1156), 
        .Q(\u_decoder/fir_filter/n1034 ) );
  NAND22 U2326 ( .A(\u_decoder/fir_filter/n1050 ), .B(
        \u_decoder/fir_filter/n1116 ), .Q(\u_decoder/fir_filter/n1418 ) );
  NAND22 U2327 ( .A(\u_decoder/fir_filter/I_data_mult_2_buff [14]), .B(n1159), 
        .Q(\u_decoder/fir_filter/n1116 ) );
  NAND22 U2328 ( .A(\u_decoder/fir_filter/n1050 ), .B(
        \u_decoder/fir_filter/n1115 ), .Q(\u_decoder/fir_filter/n1417 ) );
  NAND22 U2329 ( .A(\u_decoder/fir_filter/I_data_mult_2_buff [13]), .B(n1159), 
        .Q(\u_decoder/fir_filter/n1115 ) );
  NAND22 U2330 ( .A(\u_decoder/fir_filter/n1050 ), .B(
        \u_decoder/fir_filter/n1052 ), .Q(\u_decoder/fir_filter/n1370 ) );
  NAND22 U2331 ( .A(\u_decoder/fir_filter/I_data_mult_6_buff [14]), .B(n1157), 
        .Q(\u_decoder/fir_filter/n1052 ) );
  NAND22 U2332 ( .A(\u_decoder/fir_filter/n1050 ), .B(
        \u_decoder/fir_filter/n1051 ), .Q(\u_decoder/fir_filter/n1369 ) );
  NAND22 U2333 ( .A(\u_decoder/fir_filter/I_data_mult_6_buff [13]), .B(n1157), 
        .Q(\u_decoder/fir_filter/n1051 ) );
  NAND22 U2334 ( .A(\u_decoder/fir_filter/n722 ), .B(
        \u_decoder/fir_filter/n851 ), .Q(\u_decoder/fir_filter/n1302 ) );
  NAND22 U2335 ( .A(\u_decoder/fir_filter/Q_data_mult_0_buff [14]), .B(n1151), 
        .Q(\u_decoder/fir_filter/n851 ) );
  NAND22 U2336 ( .A(\u_decoder/fir_filter/n722 ), .B(
        \u_decoder/fir_filter/n850 ), .Q(\u_decoder/fir_filter/n1301 ) );
  NAND22 U2337 ( .A(\u_decoder/fir_filter/Q_data_mult_0_buff [13]), .B(n1151), 
        .Q(\u_decoder/fir_filter/n850 ) );
  NAND22 U2338 ( .A(\u_decoder/fir_filter/n722 ), .B(
        \u_decoder/fir_filter/n849 ), .Q(\u_decoder/fir_filter/n1300 ) );
  NAND22 U2339 ( .A(\u_decoder/fir_filter/Q_data_mult_0_buff [12]), .B(n1151), 
        .Q(\u_decoder/fir_filter/n849 ) );
  NAND22 U2340 ( .A(\u_decoder/fir_filter/n736 ), .B(
        \u_decoder/fir_filter/n835 ), .Q(\u_decoder/fir_filter/n1286 ) );
  NAND22 U2341 ( .A(\u_decoder/fir_filter/Q_data_mult_1_buff [14]), .B(n1152), 
        .Q(\u_decoder/fir_filter/n835 ) );
  NAND22 U2342 ( .A(\u_decoder/fir_filter/n736 ), .B(
        \u_decoder/fir_filter/n834 ), .Q(\u_decoder/fir_filter/n1285 ) );
  NAND22 U2343 ( .A(\u_decoder/fir_filter/Q_data_mult_1_buff [13]), .B(n1152), 
        .Q(\u_decoder/fir_filter/n834 ) );
  NAND22 U2344 ( .A(\u_decoder/fir_filter/n753 ), .B(
        \u_decoder/fir_filter/n819 ), .Q(\u_decoder/fir_filter/n1270 ) );
  NAND22 U2345 ( .A(\u_decoder/fir_filter/Q_data_mult_2_buff [14]), .B(n1151), 
        .Q(\u_decoder/fir_filter/n819 ) );
  NAND22 U2346 ( .A(\u_decoder/fir_filter/n753 ), .B(
        \u_decoder/fir_filter/n818 ), .Q(\u_decoder/fir_filter/n1269 ) );
  NAND22 U2347 ( .A(\u_decoder/fir_filter/Q_data_mult_2_buff [13]), .B(n1152), 
        .Q(\u_decoder/fir_filter/n818 ) );
  NAND22 U2348 ( .A(\u_decoder/fir_filter/n753 ), .B(
        \u_decoder/fir_filter/n755 ), .Q(\u_decoder/fir_filter/n1222 ) );
  NAND22 U2349 ( .A(\u_decoder/fir_filter/Q_data_mult_6_buff [14]), .B(n1155), 
        .Q(\u_decoder/fir_filter/n755 ) );
  NAND22 U2350 ( .A(\u_decoder/fir_filter/n753 ), .B(
        \u_decoder/fir_filter/n754 ), .Q(\u_decoder/fir_filter/n1221 ) );
  NAND22 U2351 ( .A(\u_decoder/fir_filter/Q_data_mult_6_buff [13]), .B(n1155), 
        .Q(\u_decoder/fir_filter/n754 ) );
  NAND22 U2352 ( .A(\u_decoder/fir_filter/n736 ), .B(
        \u_decoder/fir_filter/n738 ), .Q(\u_decoder/fir_filter/n1206 ) );
  NAND22 U2353 ( .A(\u_decoder/fir_filter/Q_data_mult_7_buff [14]), .B(n1154), 
        .Q(\u_decoder/fir_filter/n738 ) );
  NAND22 U2354 ( .A(\u_decoder/fir_filter/n736 ), .B(
        \u_decoder/fir_filter/n737 ), .Q(\u_decoder/fir_filter/n1205 ) );
  NAND22 U2355 ( .A(\u_decoder/fir_filter/Q_data_mult_7_buff [13]), .B(n1154), 
        .Q(\u_decoder/fir_filter/n737 ) );
  INV3 U2356 ( .A(\u_decoder/fir_filter/n1080 ), .Q(n2265) );
  AOI221 U2357 ( .A(\u_decoder/fir_filter/I_data_mult_4 [10]), .B(n1090), .C(
        \u_decoder/fir_filter/I_data_mult_4_buff [10]), .D(n1163), .Q(
        \u_decoder/fir_filter/n1080 ) );
  IMUX21 U2358 ( .A(n2949), .B(n2950), .S(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/A2[8] ), .Q(n2948) );
  INV3 U2359 ( .A(\u_decoder/fir_filter/n783 ), .Q(n2336) );
  AOI221 U2360 ( .A(\u_decoder/fir_filter/Q_data_mult_4 [10]), .B(n1084), .C(
        \u_decoder/fir_filter/Q_data_mult_4_buff [10]), .D(n1166), .Q(
        \u_decoder/fir_filter/n783 ) );
  IMUX21 U2361 ( .A(n2863), .B(n2864), .S(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/A2[8] ), .Q(n2862) );
  XNR21 U2362 ( .A(n1193), .B(n2952), .Q(
        \u_decoder/fir_filter/I_data_mult_4 [14]) );
  INV3 U2363 ( .A(\u_decoder/fir_filter/n1082 ), .Q(n2256) );
  AOI221 U2364 ( .A(\u_decoder/fir_filter/I_data_mult_4 [12]), .B(n1090), .C(
        \u_decoder/fir_filter/I_data_mult_4_buff [12]), .D(n1163), .Q(
        \u_decoder/fir_filter/n1082 ) );
  XOR21 U2365 ( .A(n2962), .B(n2963), .Q(
        \u_decoder/fir_filter/I_data_mult_4 [12]) );
  NAND22 U2366 ( .A(n2257), .B(n2959), .Q(n2963) );
  XNR21 U2367 ( .A(n1195), .B(n2866), .Q(
        \u_decoder/fir_filter/Q_data_mult_4 [14]) );
  INV3 U2368 ( .A(\u_decoder/fir_filter/n785 ), .Q(n2327) );
  AOI221 U2369 ( .A(\u_decoder/fir_filter/Q_data_mult_4 [12]), .B(n1083), .C(
        \u_decoder/fir_filter/Q_data_mult_4_buff [12]), .D(n1158), .Q(
        \u_decoder/fir_filter/n785 ) );
  XOR21 U2370 ( .A(n2876), .B(n2877), .Q(
        \u_decoder/fir_filter/Q_data_mult_4 [12]) );
  NAND22 U2371 ( .A(n2328), .B(n2873), .Q(n2877) );
  INV3 U2372 ( .A(\u_decoder/fir_filter/n983 ), .Q(n2623) );
  AOI221 U2373 ( .A(\u_decoder/fir_filter/I_data_add_7 [13]), .B(n1092), .C(
        \u_decoder/fir_filter/I_data_add_7_buff [13]), .D(n1165), .Q(
        \u_decoder/fir_filter/n983 ) );
  INV3 U2374 ( .A(\u_decoder/fir_filter/n982 ), .Q(n2622) );
  AOI221 U2375 ( .A(\u_decoder/fir_filter/I_data_add_7 [14]), .B(n1092), .C(
        \u_decoder/fir_filter/I_data_add_7_buff [14]), .D(n1165), .Q(
        \u_decoder/fir_filter/n982 ) );
  INV3 U2376 ( .A(\u_decoder/fir_filter/n962 ), .Q(n2608) );
  AOI221 U2377 ( .A(\u_decoder/fir_filter/I_data_add_6 [13]), .B(n1093), .C(
        \u_decoder/fir_filter/I_data_add_6_buff [13]), .D(n1165), .Q(
        \u_decoder/fir_filter/n962 ) );
  INV3 U2378 ( .A(\u_decoder/fir_filter/n961 ), .Q(n2607) );
  AOI221 U2379 ( .A(\u_decoder/fir_filter/I_data_add_6 [14]), .B(n1093), .C(
        \u_decoder/fir_filter/I_data_add_6_buff [14]), .D(n1166), .Q(
        \u_decoder/fir_filter/n961 ) );
  INV3 U2380 ( .A(\u_decoder/fir_filter/n941 ), .Q(n2593) );
  AOI221 U2381 ( .A(\u_decoder/fir_filter/I_data_add_5 [13]), .B(n1094), .C(
        \u_decoder/fir_filter/I_data_add_5_buff [13]), .D(n1166), .Q(
        \u_decoder/fir_filter/n941 ) );
  INV3 U2382 ( .A(\u_decoder/fir_filter/n940 ), .Q(n2592) );
  AOI221 U2383 ( .A(\u_decoder/fir_filter/I_data_add_5 [14]), .B(n1094), .C(
        \u_decoder/fir_filter/I_data_add_5_buff [14]), .D(n1166), .Q(
        \u_decoder/fir_filter/n940 ) );
  INV3 U2384 ( .A(\u_decoder/fir_filter/n899 ), .Q(n2563) );
  AOI221 U2385 ( .A(\u_decoder/fir_filter/I_data_add_3 [13]), .B(n1095), .C(
        \u_decoder/fir_filter/I_data_add_3_buff [13]), .D(n1156), .Q(
        \u_decoder/fir_filter/n899 ) );
  INV3 U2386 ( .A(\u_decoder/fir_filter/n898 ), .Q(n2562) );
  AOI221 U2387 ( .A(\u_decoder/fir_filter/I_data_add_3 [14]), .B(n1096), .C(
        \u_decoder/fir_filter/I_data_add_3_buff [14]), .D(n1151), .Q(
        \u_decoder/fir_filter/n898 ) );
  INV3 U2388 ( .A(\u_decoder/fir_filter/n878 ), .Q(n2548) );
  AOI221 U2389 ( .A(\u_decoder/fir_filter/I_data_add_2 [13]), .B(n1096), .C(
        \u_decoder/fir_filter/I_data_add_2_buff [13]), .D(n1159), .Q(
        \u_decoder/fir_filter/n878 ) );
  INV3 U2390 ( .A(\u_decoder/fir_filter/n877 ), .Q(n2547) );
  AOI221 U2391 ( .A(\u_decoder/fir_filter/I_data_add_2 [14]), .B(n1096), .C(
        \u_decoder/fir_filter/I_data_add_2_buff [14]), .D(n1157), .Q(
        \u_decoder/fir_filter/n877 ) );
  INV3 U2392 ( .A(\u_decoder/fir_filter/n857 ), .Q(n2524) );
  AOI221 U2393 ( .A(\u_decoder/fir_filter/I_data_add_1 [13]), .B(n1097), .C(
        \u_decoder/fir_filter/I_data_add_1_buff [13]), .D(n1161), .Q(
        \u_decoder/fir_filter/n857 ) );
  INV3 U2394 ( .A(\u_decoder/fir_filter/n856 ), .Q(n2523) );
  AOI221 U2395 ( .A(\u_decoder/fir_filter/I_data_add_1 [14]), .B(n1097), .C(
        \u_decoder/fir_filter/I_data_add_1_buff [14]), .D(n1156), .Q(
        \u_decoder/fir_filter/n856 ) );
  INV3 U2396 ( .A(\u_decoder/fir_filter/n853 ), .Q(n2520) );
  AOI221 U2397 ( .A(\u_decoder/fir_filter/I_data_add_0 [13]), .B(n1097), .C(
        sig_decod_outI[2]), .D(n1156), .Q(\u_decoder/fir_filter/n853 ) );
  INV3 U2398 ( .A(\u_decoder/fir_filter/n852 ), .Q(n2519) );
  AOI221 U2399 ( .A(\u_decoder/fir_filter/I_data_add_0 [14]), .B(n1149), .C(
        sig_decod_outI[3]), .D(n1152), .Q(\u_decoder/fir_filter/n852 ) );
  INV3 U2400 ( .A(\u_decoder/fir_filter/n685 ), .Q(n2503) );
  AOI221 U2401 ( .A(\u_decoder/fir_filter/Q_data_add_7 [13]), .B(n1085), .C(
        \u_decoder/fir_filter/Q_data_add_7_buff [13]), .D(n1165), .Q(
        \u_decoder/fir_filter/n685 ) );
  INV3 U2402 ( .A(\u_decoder/fir_filter/n684 ), .Q(n2502) );
  AOI221 U2403 ( .A(\u_decoder/fir_filter/Q_data_add_7 [14]), .B(n1087), .C(
        \u_decoder/fir_filter/Q_data_add_7_buff [14]), .D(n1166), .Q(
        \u_decoder/fir_filter/n684 ) );
  INV3 U2404 ( .A(\u_decoder/fir_filter/n664 ), .Q(n2488) );
  AOI221 U2405 ( .A(\u_decoder/fir_filter/Q_data_add_6 [13]), .B(n1086), .C(
        \u_decoder/fir_filter/Q_data_add_6_buff [13]), .D(n1163), .Q(
        \u_decoder/fir_filter/n664 ) );
  INV3 U2406 ( .A(\u_decoder/fir_filter/n663 ), .Q(n2487) );
  AOI221 U2407 ( .A(\u_decoder/fir_filter/Q_data_add_6 [14]), .B(n1086), .C(
        \u_decoder/fir_filter/Q_data_add_6_buff [14]), .D(n1164), .Q(
        \u_decoder/fir_filter/n663 ) );
  INV3 U2408 ( .A(\u_decoder/fir_filter/n643 ), .Q(n2473) );
  AOI221 U2409 ( .A(\u_decoder/fir_filter/Q_data_add_5 [13]), .B(n1086), .C(
        \u_decoder/fir_filter/Q_data_add_5_buff [13]), .D(n1157), .Q(
        \u_decoder/fir_filter/n643 ) );
  INV3 U2410 ( .A(\u_decoder/fir_filter/n642 ), .Q(n2472) );
  AOI221 U2411 ( .A(\u_decoder/fir_filter/Q_data_add_5 [14]), .B(n1086), .C(
        \u_decoder/fir_filter/Q_data_add_5_buff [14]), .D(n1159), .Q(
        \u_decoder/fir_filter/n642 ) );
  INV3 U2412 ( .A(\u_decoder/fir_filter/n601 ), .Q(n2443) );
  AOI221 U2413 ( .A(\u_decoder/fir_filter/Q_data_add_3 [13]), .B(n1088), .C(
        \u_decoder/fir_filter/Q_data_add_3_buff [13]), .D(n1161), .Q(
        \u_decoder/fir_filter/n601 ) );
  INV3 U2414 ( .A(\u_decoder/fir_filter/n600 ), .Q(n2442) );
  AOI221 U2415 ( .A(\u_decoder/fir_filter/Q_data_add_3 [14]), .B(n1088), .C(
        \u_decoder/fir_filter/Q_data_add_3_buff [14]), .D(n1161), .Q(
        \u_decoder/fir_filter/n600 ) );
  INV3 U2416 ( .A(\u_decoder/fir_filter/n580 ), .Q(n2428) );
  AOI221 U2417 ( .A(\u_decoder/fir_filter/Q_data_add_2 [13]), .B(n1089), .C(
        \u_decoder/fir_filter/Q_data_add_2_buff [13]), .D(n1162), .Q(
        \u_decoder/fir_filter/n580 ) );
  INV3 U2418 ( .A(\u_decoder/fir_filter/n579 ), .Q(n2427) );
  AOI221 U2419 ( .A(\u_decoder/fir_filter/Q_data_add_2 [14]), .B(n1089), .C(
        \u_decoder/fir_filter/Q_data_add_2_buff [14]), .D(n1161), .Q(
        \u_decoder/fir_filter/n579 ) );
  INV3 U2420 ( .A(\u_decoder/fir_filter/n559 ), .Q(n2404) );
  AOI221 U2421 ( .A(\u_decoder/fir_filter/Q_data_add_1 [13]), .B(n1090), .C(
        \u_decoder/fir_filter/Q_data_add_1_buff [13]), .D(n1158), .Q(
        \u_decoder/fir_filter/n559 ) );
  INV3 U2422 ( .A(\u_decoder/fir_filter/n558 ), .Q(n2403) );
  AOI221 U2423 ( .A(\u_decoder/fir_filter/Q_data_add_1 [14]), .B(n1090), .C(
        \u_decoder/fir_filter/Q_data_add_1_buff [14]), .D(n1161), .Q(
        \u_decoder/fir_filter/n558 ) );
  INV3 U2424 ( .A(\u_decoder/fir_filter/n555 ), .Q(n2400) );
  AOI221 U2425 ( .A(\u_decoder/fir_filter/Q_data_add_0 [13]), .B(n1090), .C(
        sig_decod_outQ[2]), .D(n1151), .Q(\u_decoder/fir_filter/n555 ) );
  INV3 U2426 ( .A(\u_decoder/fir_filter/n553 ), .Q(n2399) );
  AOI221 U2427 ( .A(\u_decoder/fir_filter/Q_data_add_0 [14]), .B(n1090), .C(
        sig_decod_outQ[3]), .D(n1163), .Q(\u_decoder/fir_filter/n553 ) );
  NOR21 U2428 ( .A(\u_decoder/iq_demod/sin_out [1]), .B(
        \u_decoder/iq_demod/Q_if_buff[3] ), .Q(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/ab[3][1] ) );
  NOR21 U2429 ( .A(\u_decoder/iq_demod/cos_out [1]), .B(
        \u_decoder/iq_demod/Q_if_buff[3] ), .Q(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/ab[3][1] ) );
  NOR21 U2430 ( .A(\u_decoder/iq_demod/sin_out [1]), .B(
        \u_decoder/iq_demod/I_if_buff[3] ), .Q(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/ab[3][1] ) );
  NOR21 U2431 ( .A(\u_decoder/iq_demod/cos_out [1]), .B(
        \u_decoder/iq_demod/I_if_buff[3] ), .Q(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/ab[3][1] ) );
  NOR21 U2432 ( .A(\u_decoder/iq_demod/Q_if_signed [2]), .B(n23), .Q(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/ab[2][3] ) );
  NOR21 U2433 ( .A(\u_decoder/iq_demod/sin_out [2]), .B(
        \u_decoder/iq_demod/Q_if_buff[3] ), .Q(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/ab[3][2] ) );
  NOR21 U2434 ( .A(\u_decoder/iq_demod/Q_if_signed [2]), .B(n22), .Q(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/ab[2][3] ) );
  NOR21 U2435 ( .A(\u_decoder/iq_demod/cos_out [2]), .B(
        \u_decoder/iq_demod/Q_if_buff[3] ), .Q(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/ab[3][2] ) );
  NOR21 U2436 ( .A(\u_decoder/iq_demod/I_if_signed [2]), .B(n23), .Q(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/ab[2][3] ) );
  NOR21 U2437 ( .A(\u_decoder/iq_demod/sin_out [2]), .B(
        \u_decoder/iq_demod/I_if_buff[3] ), .Q(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/ab[3][2] ) );
  NOR21 U2438 ( .A(\u_decoder/iq_demod/I_if_signed [2]), .B(n22), .Q(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/ab[2][3] ) );
  NOR21 U2439 ( .A(\u_decoder/iq_demod/cos_out [2]), .B(
        \u_decoder/iq_demod/I_if_buff[3] ), .Q(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/ab[3][2] ) );
  INV3 U2440 ( .A(\u_decoder/fir_filter/n1079 ), .Q(n2267) );
  AOI221 U2441 ( .A(\u_decoder/fir_filter/I_data_mult_4 [9]), .B(n1091), .C(
        \u_decoder/fir_filter/I_data_mult_4_buff [9]), .D(n1163), .Q(
        \u_decoder/fir_filter/n1079 ) );
  INV3 U2442 ( .A(\u_decoder/fir_filter/n782 ), .Q(n2338) );
  AOI221 U2443 ( .A(\u_decoder/fir_filter/Q_data_mult_4 [9]), .B(n1083), .C(
        \u_decoder/fir_filter/Q_data_mult_4_buff [9]), .D(n1164), .Q(
        \u_decoder/fir_filter/n782 ) );
  INV3 U2444 ( .A(\u_coder/n268 ), .Q(n1929) );
  AOI221 U2445 ( .A(\u_coder/n263 ), .B(\u_coder/j [13]), .C(n2169), .D(
        \u_coder/N1026 ), .Q(\u_coder/n268 ) );
  INV3 U2446 ( .A(\u_coder/n290 ), .Q(n1949) );
  AOI221 U2447 ( .A(n891), .B(\u_coder/i [13]), .C(n2156), .D(\u_coder/N720 ), 
        .Q(\u_coder/n290 ) );
  INV3 U2448 ( .A(\u_coder/n269 ), .Q(n1928) );
  AOI221 U2449 ( .A(n890), .B(\u_coder/j [12]), .C(n2169), .D(\u_coder/N1025 ), 
        .Q(\u_coder/n269 ) );
  INV3 U2450 ( .A(\u_coder/n291 ), .Q(n1948) );
  AOI221 U2451 ( .A(n892), .B(\u_coder/i [12]), .C(n2156), .D(\u_coder/N719 ), 
        .Q(\u_coder/n291 ) );
  INV3 U2452 ( .A(\u_decoder/fir_filter/n625 ), .Q(n2461) );
  AOI221 U2453 ( .A(\u_decoder/fir_filter/Q_data_add_4 [10]), .B(n1087), .C(
        \u_decoder/fir_filter/Q_data_add_4_buff [10]), .D(n1162), .Q(
        \u_decoder/fir_filter/n625 ) );
  INV3 U2454 ( .A(\u_decoder/fir_filter/n923 ), .Q(n2581) );
  AOI221 U2455 ( .A(\u_decoder/fir_filter/I_data_add_4 [10]), .B(n1094), .C(
        \u_decoder/fir_filter/I_data_add_4_buff [10]), .D(n1160), .Q(
        \u_decoder/fir_filter/n923 ) );
  NOR21 U2456 ( .A(\u_decoder/iq_demod/Q_if_signed [0]), .B(n23), .Q(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/ab[0][3] ) );
  NOR21 U2457 ( .A(\u_decoder/iq_demod/Q_if_signed [0]), .B(n22), .Q(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/ab[0][3] ) );
  NOR21 U2458 ( .A(\u_decoder/iq_demod/I_if_signed [0]), .B(n23), .Q(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/ab[0][3] ) );
  NOR21 U2459 ( .A(\u_decoder/iq_demod/I_if_signed [0]), .B(n22), .Q(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/ab[0][3] ) );
  NOR21 U2460 ( .A(\u_decoder/iq_demod/Q_if_signed [1]), .B(n23), .Q(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/ab[1][3] ) );
  NOR21 U2461 ( .A(n124), .B(n45), .Q(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/ab[2][2] ) );
  NOR21 U2462 ( .A(n698), .B(n699), .Q(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/CARRYB[1][2] ) );
  NOR21 U2463 ( .A(\u_decoder/iq_demod/Q_if_signed [1]), .B(n22), .Q(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/ab[1][3] ) );
  NOR21 U2464 ( .A(n124), .B(n43), .Q(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/ab[2][2] ) );
  NOR21 U2465 ( .A(n722), .B(n723), .Q(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/CARRYB[1][2] ) );
  NOR21 U2466 ( .A(\u_decoder/iq_demod/I_if_signed [1]), .B(n23), .Q(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/ab[1][3] ) );
  NOR21 U2467 ( .A(n125), .B(n45), .Q(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/ab[2][2] ) );
  NOR21 U2468 ( .A(n734), .B(n735), .Q(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/CARRYB[1][2] ) );
  NOR21 U2469 ( .A(\u_decoder/iq_demod/I_if_signed [1]), .B(n22), .Q(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/ab[1][3] ) );
  NOR21 U2470 ( .A(n125), .B(n43), .Q(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/ab[2][2] ) );
  NOR21 U2471 ( .A(n710), .B(n711), .Q(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/CARRYB[1][2] ) );
  NOR21 U2472 ( .A(\u_decoder/iq_demod/sin_out [0]), .B(
        \u_decoder/iq_demod/Q_if_buff[3] ), .Q(
        \u_decoder/iq_demod/dp_cluster_0/mult_151/ab[3][0] ) );
  NOR21 U2473 ( .A(\u_decoder/iq_demod/cos_out [0]), .B(
        \u_decoder/iq_demod/Q_if_buff[3] ), .Q(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/ab[3][0] ) );
  NOR21 U2474 ( .A(\u_decoder/iq_demod/sin_out [0]), .B(
        \u_decoder/iq_demod/I_if_buff[3] ), .Q(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/ab[3][0] ) );
  NOR21 U2475 ( .A(\u_decoder/iq_demod/cos_out [0]), .B(
        \u_decoder/iq_demod/I_if_buff[3] ), .Q(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/ab[3][0] ) );
  NAND22 U2476 ( .A(\u_decoder/fir_filter/I_data_mult_1_buff [11]), .B(n1160), 
        .Q(\u_decoder/fir_filter/n1129 ) );
  NAND22 U2477 ( .A(\u_decoder/fir_filter/I_data_mult_1_buff [10]), .B(n1160), 
        .Q(\u_decoder/fir_filter/n1128 ) );
  NAND22 U2478 ( .A(\u_decoder/fir_filter/I_data_mult_1_buff [9]), .B(n1160), 
        .Q(\u_decoder/fir_filter/n1127 ) );
  NAND22 U2479 ( .A(\u_decoder/fir_filter/I_data_mult_2_buff [10]), .B(n1159), 
        .Q(\u_decoder/fir_filter/n1112 ) );
  NAND22 U2480 ( .A(\u_decoder/fir_filter/I_data_mult_2_buff [9]), .B(n1159), 
        .Q(\u_decoder/fir_filter/n1111 ) );
  NAND22 U2481 ( .A(\u_decoder/fir_filter/I_data_mult_6_buff [10]), .B(n1157), 
        .Q(\u_decoder/fir_filter/n1047 ) );
  NAND22 U2482 ( .A(\u_decoder/fir_filter/I_data_mult_6_buff [9]), .B(n1157), 
        .Q(\u_decoder/fir_filter/n1046 ) );
  NAND22 U2483 ( .A(\u_decoder/fir_filter/I_data_mult_7_buff [11]), .B(n1156), 
        .Q(\u_decoder/fir_filter/n1031 ) );
  NAND22 U2484 ( .A(\u_decoder/fir_filter/I_data_mult_7_buff [10]), .B(n1156), 
        .Q(\u_decoder/fir_filter/n1030 ) );
  NAND22 U2485 ( .A(\u_decoder/fir_filter/I_data_mult_7_buff [9]), .B(n1156), 
        .Q(\u_decoder/fir_filter/n1029 ) );
  NAND22 U2486 ( .A(\u_decoder/fir_filter/Q_data_mult_1_buff [11]), .B(n1152), 
        .Q(\u_decoder/fir_filter/n832 ) );
  NAND22 U2487 ( .A(\u_decoder/fir_filter/Q_data_mult_1_buff [10]), .B(n1152), 
        .Q(\u_decoder/fir_filter/n831 ) );
  NAND22 U2488 ( .A(\u_decoder/fir_filter/Q_data_mult_1_buff [9]), .B(n1152), 
        .Q(\u_decoder/fir_filter/n830 ) );
  NAND22 U2489 ( .A(\u_decoder/fir_filter/Q_data_mult_2_buff [10]), .B(n1152), 
        .Q(\u_decoder/fir_filter/n815 ) );
  NAND22 U2490 ( .A(\u_decoder/fir_filter/Q_data_mult_2_buff [9]), .B(n1157), 
        .Q(\u_decoder/fir_filter/n814 ) );
  NAND22 U2491 ( .A(\u_decoder/fir_filter/Q_data_mult_6_buff [10]), .B(n1154), 
        .Q(\u_decoder/fir_filter/n750 ) );
  NAND22 U2492 ( .A(\u_decoder/fir_filter/Q_data_mult_6_buff [9]), .B(n1156), 
        .Q(\u_decoder/fir_filter/n749 ) );
  NAND22 U2493 ( .A(\u_decoder/fir_filter/Q_data_mult_7_buff [11]), .B(n1154), 
        .Q(\u_decoder/fir_filter/n734 ) );
  NAND22 U2494 ( .A(\u_decoder/fir_filter/Q_data_mult_7_buff [10]), .B(n1154), 
        .Q(\u_decoder/fir_filter/n733 ) );
  NAND22 U2495 ( .A(\u_decoder/fir_filter/Q_data_mult_7_buff [9]), .B(n1154), 
        .Q(\u_decoder/fir_filter/n732 ) );
  NAND22 U2496 ( .A(\u_decoder/fir_filter/I_data_mult_0_buff [10]), .B(n1160), 
        .Q(\u_decoder/fir_filter/n1144 ) );
  NAND22 U2497 ( .A(\u_decoder/fir_filter/I_data_mult_0_buff [9]), .B(n1153), 
        .Q(\u_decoder/fir_filter/n1143 ) );
  NAND22 U2498 ( .A(\u_decoder/fir_filter/Q_data_mult_0_buff [10]), .B(n1151), 
        .Q(\u_decoder/fir_filter/n847 ) );
  NAND22 U2499 ( .A(\u_decoder/fir_filter/Q_data_mult_0_buff [9]), .B(n1152), 
        .Q(\u_decoder/fir_filter/n846 ) );
  NAND22 U2500 ( .A(\u_decoder/fir_filter/I_data_mult_0_buff [8]), .B(n1160), 
        .Q(\u_decoder/fir_filter/n1142 ) );
  NAND22 U2501 ( .A(\u_decoder/fir_filter/Q_data_mult_0_buff [8]), .B(n1153), 
        .Q(\u_decoder/fir_filter/n845 ) );
  INV3 U2502 ( .A(\u_coder/n270 ), .Q(n1927) );
  AOI221 U2503 ( .A(\u_coder/n263 ), .B(\u_coder/j [11]), .C(n2169), .D(
        \u_coder/N1024 ), .Q(\u_coder/n270 ) );
  INV3 U2504 ( .A(\u_coder/n292 ), .Q(n1947) );
  AOI221 U2505 ( .A(n891), .B(\u_coder/i [11]), .C(n2156), .D(\u_coder/N718 ), 
        .Q(\u_coder/n292 ) );
  INV3 U2506 ( .A(\u_decoder/fir_filter/n1081 ), .Q(n2261) );
  AOI221 U2507 ( .A(\u_decoder/fir_filter/I_data_mult_4 [11]), .B(n1090), .C(
        \u_decoder/fir_filter/I_data_mult_4_buff [11]), .D(n1163), .Q(
        \u_decoder/fir_filter/n1081 ) );
  XNR21 U2508 ( .A(n2943), .B(n2944), .Q(
        \u_decoder/fir_filter/I_data_mult_4 [11]) );
  NAND22 U2509 ( .A(n2262), .B(n2945), .Q(n2944) );
  INV3 U2510 ( .A(\u_decoder/fir_filter/n784 ), .Q(n2332) );
  AOI221 U2511 ( .A(\u_decoder/fir_filter/Q_data_mult_4 [11]), .B(n1083), .C(
        \u_decoder/fir_filter/Q_data_mult_4_buff [11]), .D(n1165), .Q(
        \u_decoder/fir_filter/n784 ) );
  XNR21 U2512 ( .A(n2857), .B(n2858), .Q(
        \u_decoder/fir_filter/Q_data_mult_4 [11]) );
  NAND22 U2513 ( .A(n2333), .B(n2859), .Q(n2858) );
  INV3 U2514 ( .A(\u_decoder/fir_filter/n986 ), .Q(n2626) );
  AOI221 U2515 ( .A(\u_decoder/fir_filter/I_data_add_7 [10]), .B(n1092), .C(
        \u_decoder/fir_filter/I_data_add_7_buff [10]), .D(n1164), .Q(
        \u_decoder/fir_filter/n986 ) );
  INV3 U2516 ( .A(\u_decoder/fir_filter/n985 ), .Q(n2625) );
  AOI221 U2517 ( .A(\u_decoder/fir_filter/I_data_add_7 [11]), .B(n1092), .C(
        \u_decoder/fir_filter/I_data_add_7_buff [11]), .D(n1165), .Q(
        \u_decoder/fir_filter/n985 ) );
  INV3 U2518 ( .A(\u_decoder/fir_filter/n984 ), .Q(n2624) );
  AOI221 U2519 ( .A(\u_decoder/fir_filter/I_data_add_7 [12]), .B(n1092), .C(
        \u_decoder/fir_filter/I_data_add_7_buff [12]), .D(n1165), .Q(
        \u_decoder/fir_filter/n984 ) );
  INV3 U2520 ( .A(\u_decoder/fir_filter/n965 ), .Q(n2611) );
  AOI221 U2521 ( .A(\u_decoder/fir_filter/I_data_add_6 [10]), .B(n1093), .C(
        \u_decoder/fir_filter/I_data_add_6_buff [10]), .D(n1165), .Q(
        \u_decoder/fir_filter/n965 ) );
  INV3 U2522 ( .A(\u_decoder/fir_filter/n964 ), .Q(n2610) );
  AOI221 U2523 ( .A(\u_decoder/fir_filter/I_data_add_6 [11]), .B(n1093), .C(
        \u_decoder/fir_filter/I_data_add_6_buff [11]), .D(n1165), .Q(
        \u_decoder/fir_filter/n964 ) );
  INV3 U2524 ( .A(\u_decoder/fir_filter/n963 ), .Q(n2609) );
  AOI221 U2525 ( .A(\u_decoder/fir_filter/I_data_add_6 [12]), .B(n1093), .C(
        \u_decoder/fir_filter/I_data_add_6_buff [12]), .D(n1165), .Q(
        \u_decoder/fir_filter/n963 ) );
  INV3 U2526 ( .A(\u_decoder/fir_filter/n944 ), .Q(n2596) );
  AOI221 U2527 ( .A(\u_decoder/fir_filter/I_data_add_5 [10]), .B(n1093), .C(
        \u_decoder/fir_filter/I_data_add_5_buff [10]), .D(n1166), .Q(
        \u_decoder/fir_filter/n944 ) );
  INV3 U2528 ( .A(\u_decoder/fir_filter/n943 ), .Q(n2595) );
  AOI221 U2529 ( .A(\u_decoder/fir_filter/I_data_add_5 [11]), .B(n1094), .C(
        \u_decoder/fir_filter/I_data_add_5_buff [11]), .D(n1166), .Q(
        \u_decoder/fir_filter/n943 ) );
  INV3 U2530 ( .A(\u_decoder/fir_filter/n942 ), .Q(n2594) );
  AOI221 U2531 ( .A(\u_decoder/fir_filter/I_data_add_5 [12]), .B(n1094), .C(
        \u_decoder/fir_filter/I_data_add_5_buff [12]), .D(n1166), .Q(
        \u_decoder/fir_filter/n942 ) );
  INV3 U2532 ( .A(\u_decoder/fir_filter/n922 ), .Q(n2580) );
  AOI221 U2533 ( .A(\u_decoder/fir_filter/I_data_add_4 [11]), .B(n1094), .C(
        \u_decoder/fir_filter/I_data_add_4_buff [11]), .D(n1166), .Q(
        \u_decoder/fir_filter/n922 ) );
  INV3 U2534 ( .A(\u_decoder/fir_filter/n921 ), .Q(n2579) );
  AOI221 U2535 ( .A(\u_decoder/fir_filter/I_data_add_4 [12]), .B(n1095), .C(
        \u_decoder/fir_filter/I_data_add_4_buff [12]), .D(n1163), .Q(
        \u_decoder/fir_filter/n921 ) );
  INV3 U2536 ( .A(\u_decoder/fir_filter/n902 ), .Q(n2566) );
  AOI221 U2537 ( .A(\u_decoder/fir_filter/I_data_add_3 [10]), .B(n1095), .C(
        \u_decoder/fir_filter/I_data_add_3_buff [10]), .D(n1155), .Q(
        \u_decoder/fir_filter/n902 ) );
  INV3 U2538 ( .A(\u_decoder/fir_filter/n901 ), .Q(n2565) );
  AOI221 U2539 ( .A(\u_decoder/fir_filter/I_data_add_3 [11]), .B(n1095), .C(
        \u_decoder/fir_filter/I_data_add_3_buff [11]), .D(n1160), .Q(
        \u_decoder/fir_filter/n901 ) );
  INV3 U2540 ( .A(\u_decoder/fir_filter/n900 ), .Q(n2564) );
  AOI221 U2541 ( .A(\u_decoder/fir_filter/I_data_add_3 [12]), .B(n1095), .C(
        \u_decoder/fir_filter/I_data_add_3_buff [12]), .D(n1159), .Q(
        \u_decoder/fir_filter/n900 ) );
  INV3 U2542 ( .A(\u_decoder/fir_filter/n881 ), .Q(n2551) );
  AOI221 U2543 ( .A(\u_decoder/fir_filter/I_data_add_2 [10]), .B(n1096), .C(
        \u_decoder/fir_filter/I_data_add_2_buff [10]), .D(n1158), .Q(
        \u_decoder/fir_filter/n881 ) );
  INV3 U2544 ( .A(\u_decoder/fir_filter/n880 ), .Q(n2550) );
  AOI221 U2545 ( .A(\u_decoder/fir_filter/I_data_add_2 [11]), .B(n1096), .C(
        \u_decoder/fir_filter/I_data_add_2_buff [11]), .D(n1164), .Q(
        \u_decoder/fir_filter/n880 ) );
  INV3 U2546 ( .A(\u_decoder/fir_filter/n879 ), .Q(n2549) );
  AOI221 U2547 ( .A(\u_decoder/fir_filter/I_data_add_2 [12]), .B(n1096), .C(
        \u_decoder/fir_filter/I_data_add_2_buff [12]), .D(n1165), .Q(
        \u_decoder/fir_filter/n879 ) );
  INV3 U2548 ( .A(\u_decoder/fir_filter/n860 ), .Q(n2527) );
  AOI221 U2549 ( .A(\u_decoder/fir_filter/I_data_add_1 [10]), .B(n1097), .C(
        \u_decoder/fir_filter/I_data_add_1_buff [10]), .D(n1155), .Q(
        \u_decoder/fir_filter/n860 ) );
  INV3 U2550 ( .A(\u_decoder/fir_filter/n859 ), .Q(n2526) );
  AOI221 U2551 ( .A(\u_decoder/fir_filter/I_data_add_1 [11]), .B(n1097), .C(
        \u_decoder/fir_filter/I_data_add_1_buff [11]), .D(n1154), .Q(
        \u_decoder/fir_filter/n859 ) );
  INV3 U2552 ( .A(\u_decoder/fir_filter/n858 ), .Q(n2525) );
  AOI221 U2553 ( .A(\u_decoder/fir_filter/I_data_add_1 [12]), .B(n1097), .C(
        \u_decoder/fir_filter/I_data_add_1_buff [12]), .D(n1153), .Q(
        \u_decoder/fir_filter/n858 ) );
  INV3 U2554 ( .A(\u_decoder/fir_filter/n855 ), .Q(n2522) );
  AOI221 U2555 ( .A(\u_decoder/fir_filter/I_data_add_0 [11]), .B(n1097), .C(
        sig_decod_outI[0]), .D(n1159), .Q(\u_decoder/fir_filter/n855 ) );
  INV3 U2556 ( .A(\u_decoder/fir_filter/n854 ), .Q(n2521) );
  AOI221 U2557 ( .A(\u_decoder/fir_filter/I_data_add_0 [12]), .B(n1097), .C(
        sig_decod_outI[1]), .D(n1159), .Q(\u_decoder/fir_filter/n854 ) );
  INV3 U2558 ( .A(\u_decoder/fir_filter/n688 ), .Q(n2506) );
  AOI221 U2559 ( .A(\u_decoder/fir_filter/Q_data_add_7 [10]), .B(n1084), .C(
        \u_decoder/fir_filter/Q_data_add_7_buff [10]), .D(n1163), .Q(
        \u_decoder/fir_filter/n688 ) );
  INV3 U2560 ( .A(\u_decoder/fir_filter/n687 ), .Q(n2505) );
  AOI221 U2561 ( .A(\u_decoder/fir_filter/Q_data_add_7 [11]), .B(n1085), .C(
        \u_decoder/fir_filter/Q_data_add_7_buff [11]), .D(n1163), .Q(
        \u_decoder/fir_filter/n687 ) );
  INV3 U2562 ( .A(\u_decoder/fir_filter/n686 ), .Q(n2504) );
  AOI221 U2563 ( .A(\u_decoder/fir_filter/Q_data_add_7 [12]), .B(n1085), .C(
        \u_decoder/fir_filter/Q_data_add_7_buff [12]), .D(n1165), .Q(
        \u_decoder/fir_filter/n686 ) );
  INV3 U2564 ( .A(\u_decoder/fir_filter/n667 ), .Q(n2491) );
  AOI221 U2565 ( .A(\u_decoder/fir_filter/Q_data_add_6 [10]), .B(n1085), .C(
        \u_decoder/fir_filter/Q_data_add_6_buff [10]), .D(n1166), .Q(
        \u_decoder/fir_filter/n667 ) );
  INV3 U2566 ( .A(\u_decoder/fir_filter/n666 ), .Q(n2490) );
  AOI221 U2567 ( .A(\u_decoder/fir_filter/Q_data_add_6 [11]), .B(n1085), .C(
        \u_decoder/fir_filter/Q_data_add_6_buff [11]), .D(n1163), .Q(
        \u_decoder/fir_filter/n666 ) );
  INV3 U2568 ( .A(\u_decoder/fir_filter/n665 ), .Q(n2489) );
  AOI221 U2569 ( .A(\u_decoder/fir_filter/Q_data_add_6 [12]), .B(n1085), .C(
        \u_decoder/fir_filter/Q_data_add_6_buff [12]), .D(n1164), .Q(
        \u_decoder/fir_filter/n665 ) );
  INV3 U2570 ( .A(\u_decoder/fir_filter/n646 ), .Q(n2476) );
  AOI221 U2571 ( .A(\u_decoder/fir_filter/Q_data_add_5 [10]), .B(n1086), .C(
        \u_decoder/fir_filter/Q_data_add_5_buff [10]), .D(n1164), .Q(
        \u_decoder/fir_filter/n646 ) );
  INV3 U2572 ( .A(\u_decoder/fir_filter/n645 ), .Q(n2475) );
  AOI221 U2573 ( .A(\u_decoder/fir_filter/Q_data_add_5 [11]), .B(n1086), .C(
        \u_decoder/fir_filter/Q_data_add_5_buff [11]), .D(n1165), .Q(
        \u_decoder/fir_filter/n645 ) );
  INV3 U2574 ( .A(\u_decoder/fir_filter/n644 ), .Q(n2474) );
  AOI221 U2575 ( .A(\u_decoder/fir_filter/Q_data_add_5 [12]), .B(n1086), .C(
        \u_decoder/fir_filter/Q_data_add_5_buff [12]), .D(n1158), .Q(
        \u_decoder/fir_filter/n644 ) );
  INV3 U2576 ( .A(\u_decoder/fir_filter/n624 ), .Q(n2460) );
  AOI221 U2577 ( .A(\u_decoder/fir_filter/Q_data_add_4 [11]), .B(n1087), .C(
        \u_decoder/fir_filter/Q_data_add_4_buff [11]), .D(n1162), .Q(
        \u_decoder/fir_filter/n624 ) );
  INV3 U2578 ( .A(\u_decoder/fir_filter/n623 ), .Q(n2459) );
  AOI221 U2579 ( .A(\u_decoder/fir_filter/Q_data_add_4 [12]), .B(n1087), .C(
        \u_decoder/fir_filter/Q_data_add_4_buff [12]), .D(n1162), .Q(
        \u_decoder/fir_filter/n623 ) );
  INV3 U2580 ( .A(\u_decoder/fir_filter/n604 ), .Q(n2446) );
  AOI221 U2581 ( .A(\u_decoder/fir_filter/Q_data_add_3 [10]), .B(n1088), .C(
        \u_decoder/fir_filter/Q_data_add_3_buff [10]), .D(n1161), .Q(
        \u_decoder/fir_filter/n604 ) );
  INV3 U2582 ( .A(\u_decoder/fir_filter/n603 ), .Q(n2445) );
  AOI221 U2583 ( .A(\u_decoder/fir_filter/Q_data_add_3 [11]), .B(n1088), .C(
        \u_decoder/fir_filter/Q_data_add_3_buff [11]), .D(n1161), .Q(
        \u_decoder/fir_filter/n603 ) );
  INV3 U2584 ( .A(\u_decoder/fir_filter/n602 ), .Q(n2444) );
  AOI221 U2585 ( .A(\u_decoder/fir_filter/Q_data_add_3 [12]), .B(n1088), .C(
        \u_decoder/fir_filter/Q_data_add_3_buff [12]), .D(n1166), .Q(
        \u_decoder/fir_filter/n602 ) );
  INV3 U2586 ( .A(\u_decoder/fir_filter/n583 ), .Q(n2431) );
  AOI221 U2587 ( .A(\u_decoder/fir_filter/Q_data_add_2 [10]), .B(n1089), .C(
        \u_decoder/fir_filter/Q_data_add_2_buff [10]), .D(n1161), .Q(
        \u_decoder/fir_filter/n583 ) );
  INV3 U2588 ( .A(\u_decoder/fir_filter/n582 ), .Q(n2430) );
  AOI221 U2589 ( .A(\u_decoder/fir_filter/Q_data_add_2 [11]), .B(n1089), .C(
        \u_decoder/fir_filter/Q_data_add_2_buff [11]), .D(n1161), .Q(
        \u_decoder/fir_filter/n582 ) );
  INV3 U2590 ( .A(\u_decoder/fir_filter/n581 ), .Q(n2429) );
  AOI221 U2591 ( .A(\u_decoder/fir_filter/Q_data_add_2 [12]), .B(n1089), .C(
        \u_decoder/fir_filter/Q_data_add_2_buff [12]), .D(n1162), .Q(
        \u_decoder/fir_filter/n581 ) );
  INV3 U2592 ( .A(\u_decoder/fir_filter/n562 ), .Q(n2407) );
  AOI221 U2593 ( .A(\u_decoder/fir_filter/Q_data_add_1 [10]), .B(n1090), .C(
        \u_decoder/fir_filter/Q_data_add_1_buff [10]), .D(n1163), .Q(
        \u_decoder/fir_filter/n562 ) );
  INV3 U2594 ( .A(\u_decoder/fir_filter/n561 ), .Q(n2406) );
  AOI221 U2595 ( .A(\u_decoder/fir_filter/Q_data_add_1 [11]), .B(n1090), .C(
        \u_decoder/fir_filter/Q_data_add_1_buff [11]), .D(n1156), .Q(
        \u_decoder/fir_filter/n561 ) );
  INV3 U2596 ( .A(\u_decoder/fir_filter/n560 ), .Q(n2405) );
  AOI221 U2597 ( .A(\u_decoder/fir_filter/Q_data_add_1 [12]), .B(n1090), .C(
        \u_decoder/fir_filter/Q_data_add_1_buff [12]), .D(n1155), .Q(
        \u_decoder/fir_filter/n560 ) );
  INV3 U2598 ( .A(\u_decoder/fir_filter/n557 ), .Q(n2402) );
  AOI221 U2599 ( .A(\u_decoder/fir_filter/Q_data_add_0 [11]), .B(n1090), .C(
        sig_decod_outQ[0]), .D(n1162), .Q(\u_decoder/fir_filter/n557 ) );
  INV3 U2600 ( .A(\u_decoder/fir_filter/n556 ), .Q(n2401) );
  AOI221 U2601 ( .A(\u_decoder/fir_filter/Q_data_add_0 [12]), .B(n1090), .C(
        sig_decod_outQ[1]), .D(n1164), .Q(\u_decoder/fir_filter/n556 ) );
  AOI311 U2602 ( .A(n2706), .B(n2704), .C(n2703), .D(
        \u_inFIFO/outWriteCount[7] ), .Q(n2705) );
  OAI2111 U2603 ( .A(\u_inFIFO/outReadCount[5] ), .B(\u_inFIFO/n183 ), .C(
        n2702), .D(n2701), .Q(n2703) );
  NAND22 U2604 ( .A(\u_inFIFO/outWriteCount[4] ), .B(n162), .Q(n2701) );
  AOI221 U2605 ( .A(\sig_MUX_inMUX5[0] ), .B(n2131), .C(in_MUX_inSEL3), .D(
        sig_DEMUX_outDEMUX2[1]), .Q(n3113) );
  NOR31 U2606 ( .A(n3117), .B(in_DEMUX_inSEL2[2]), .C(in_DEMUX_inSEL2[1]), .Q(
        sig_DEMUX_outDEMUX2[1]) );
  AOI211 U2607 ( .A(\u_cordic/mycordic/present_I_table[4][1] ), .B(
        \u_cordic/mycordic/present_Q_table[4][4] ), .C(n2657), .Q(n3034) );
  INV3 U2608 ( .A(n3032), .Q(n2657) );
  OAI2111 U2609 ( .A(\u_cordic/mycordic/present_I_table[4][1] ), .B(
        \u_cordic/mycordic/present_Q_table[4][4] ), .C(
        \u_cordic/mycordic/present_I_table[4][0] ), .D(
        \u_cordic/mycordic/present_Q_table[4][3] ), .Q(n3032) );
  INV3 U2610 ( .A(n3016), .Q(n2648) );
  NAND22 U2611 ( .A(n197), .B(n3017), .Q(n3016) );
  AOI221 U2612 ( .A(n3015), .B(\u_cordic/mycordic/present_Q_table[5][1] ), .C(
        n46), .D(n2650), .Q(n3017) );
  NOR40 U2613 ( .A(n2710), .B(n2711), .C(n2150), .D(n2709), .Q(
        \sig_MUX_inMUX5[0] ) );
  INV3 U2614 ( .A(n2706), .Q(n2150) );
  NAND41 U2615 ( .A(n2704), .B(n2698), .C(n2697), .D(n2694), .Q(n2710) );
  AOI211 U2616 ( .A(\u_inFIFO/outWriteCount[1] ), .B(n2708), .C(n2149), .Q(
        n2709) );
  INV3 U2617 ( .A(n3013), .Q(n2641) );
  AOI211 U2618 ( .A(n3011), .B(\u_cordic/mycordic/present_Q_table[5][5] ), .C(
        n2642), .Q(n3013) );
  AOI221 U2619 ( .A(n3029), .B(\u_cordic/mycordic/present_I_table[4][2] ), .C(
        n227), .D(n2652), .Q(n3031) );
  INV3 U2620 ( .A(n3028), .Q(n2652) );
  NOR21 U2621 ( .A(\u_cordic/mycordic/present_I_table[4][2] ), .B(n3029), .Q(
        n3028) );
  NOR21 U2622 ( .A(n2103), .B(\u_coder/IorQ ), .Q(\u_coder/n213 ) );
  INV3 U2623 ( .A(n3113), .Q(n2103) );
  INV3 U2624 ( .A(n3034), .Q(n2656) );
  NOR31 U2625 ( .A(\u_coder/n209 ), .B(\u_coder/n210 ), .C(n1811), .Q(
        \u_coder/n179 ) );
  INV3 U2626 ( .A(\u_coder/n211 ), .Q(n1811) );
  AOI311 U2627 ( .A(\u_coder/n213 ), .B(\u_coder/n181 ), .C(\u_coder/n191 ), 
        .D(\u_coder/stateQ[0] ), .Q(\u_coder/n210 ) );
  AOI211 U2628 ( .A(n2185), .B(\u_coder/n212 ), .C(n1236), .Q(\u_coder/n211 )
         );
  INV3 U2629 ( .A(n3009), .Q(n2645) );
  AOI211 U2630 ( .A(n3007), .B(\u_cordic/mycordic/present_Q_table[5][3] ), .C(
        n2646), .Q(n3009) );
  INV3 U2631 ( .A(n3020), .Q(n2644) );
  AOI211 U2632 ( .A(n247), .B(n3021), .C(
        \u_cordic/mycordic/present_I_table[5][7] ), .Q(n3020) );
  AOI211 U2633 ( .A(n3019), .B(\u_cordic/mycordic/present_Q_table[5][3] ), .C(
        n2647), .Q(n3021) );
  INV3 U2634 ( .A(n3004), .Q(n2649) );
  OAI2111 U2635 ( .A(n2700), .B(n2699), .C(n2698), .D(n2697), .Q(n2702) );
  NOR21 U2636 ( .A(\u_inFIFO/outReadCount[3] ), .B(\u_inFIFO/n185 ), .Q(n2700)
         );
  OAI2111 U2637 ( .A(n2695), .B(n126), .C(n2147), .D(n2694), .Q(n2696) );
  OAI2111 U2638 ( .A(\u_cordic/mycordic/present_Q_table[5][1] ), .B(
        \u_cordic/mycordic/present_I_table[5][5] ), .C(
        \u_cordic/mycordic/present_Q_table[5][0] ), .D(
        \u_cordic/mycordic/present_I_table[5][4] ), .Q(n3003) );
  INV3 U2639 ( .A(\u_coder/n151 ), .Q(n1808) );
  AOI211 U2640 ( .A(sig_coder_outSinI[1]), .B(n1809), .C(\u_coder/n152 ), .Q(
        \u_coder/n151 ) );
  AOI221 U2641 ( .A(\u_coder/n149 ), .B(\u_coder/n157 ), .C(\u_coder/n137 ), 
        .D(\u_coder/n155 ), .Q(\u_coder/n153 ) );
  OAI2111 U2642 ( .A(n2152), .B(\u_coder/n182 ), .C(\u_coder/n207 ), .D(
        \u_coder/n208 ), .Q(\u_coder/n339 ) );
  INV3 U2643 ( .A(\u_coder/n219 ), .Q(n2152) );
  NAND31 U2644 ( .A(\u_coder/my_clk_10M ), .B(\u_coder/n214 ), .C(
        \u_coder/stateQ[0] ), .Q(\u_coder/n207 ) );
  NAND22 U2645 ( .A(sig_coder_outSinQ[0]), .B(\u_coder/n179 ), .Q(
        \u_coder/n208 ) );
  OAI2111 U2646 ( .A(\u_coder/n163 ), .B(\u_coder/n139 ), .C(\u_coder/n164 ), 
        .D(\u_coder/n165 ), .Q(\u_coder/n336 ) );
  AOI221 U2647 ( .A(\u_coder/n137 ), .B(\u_coder/n174 ), .C(\u_coder/n149 ), 
        .D(\u_coder/n174 ), .Q(\u_coder/n163 ) );
  NAND31 U2648 ( .A(\u_coder/stateI[0] ), .B(n2096), .C(\u_coder/my_clk_10M ), 
        .Q(\u_coder/n164 ) );
  NAND22 U2649 ( .A(sig_coder_outSinI[0]), .B(n1809), .Q(\u_coder/n165 ) );
  INV3 U2650 ( .A(\u_coder/n140 ), .Q(n1807) );
  AOI211 U2651 ( .A(sig_coder_outSinI[2]), .B(n1809), .C(\u_coder/n141 ), .Q(
        \u_coder/n140 ) );
  AOI221 U2652 ( .A(\u_coder/n149 ), .B(\u_coder/n150 ), .C(\u_coder/n137 ), 
        .D(\u_coder/n145 ), .Q(\u_coder/n142 ) );
  NAND22 U2653 ( .A(\u_coder/IorQ ), .B(n3113), .Q(\u_coder/n170 ) );
  XNR21 U2654 ( .A(\u_outFIFO/r98/carry [7]), .B(\u_outFIFO/outWriteCount[7] ), 
        .Q(\u_outFIFO/N150 ) );
  XNR21 U2655 ( .A(\u_inFIFO/r96/carry [7]), .B(\u_inFIFO/outWriteCount[7] ), 
        .Q(\u_inFIFO/N140 ) );
  INV3 U2656 ( .A(\u_cordic/mycordic/n549 ), .Q(n1545) );
  AOI221 U2657 ( .A(\u_cordic/mycordic/N395 ), .B(n778), .C(
        \u_cordic/mycordic/N427 ), .D(n1908), .Q(\u_cordic/mycordic/n549 ) );
  INV3 U2658 ( .A(\u_cordic/mycordic/n335 ), .Q(n1484) );
  AOI221 U2659 ( .A(\u_cordic/mycordic/N331 ), .B(\u_cordic/mycordic/n336 ), 
        .C(\u_cordic/mycordic/N363 ), .D(n1904), .Q(\u_cordic/mycordic/n335 )
         );
  INV3 U2660 ( .A(n3010), .Q(n2642) );
  INV3 U2661 ( .A(n3022), .Q(n2643) );
  INV3 U2662 ( .A(n3018), .Q(n2647) );
  INV3 U2663 ( .A(n3006), .Q(n2646) );
  INV3 U2664 ( .A(\u_cordic/mycordic/n362 ), .Q(n1540) );
  AOI221 U2665 ( .A(\u_cordic/mycordic/N447 ), .B(\u_cordic/mycordic/n363 ), 
        .C(\u_cordic/mycordic/N475 ), .D(n1907), .Q(\u_cordic/mycordic/n362 )
         );
  INV3 U2666 ( .A(\u_cordic/mycordic/n540 ), .Q(n1520) );
  AOI221 U2667 ( .A(\u_cordic/mycordic/N455 ), .B(\u_cordic/mycordic/n363 ), 
        .C(\u_cordic/mycordic/N483 ), .D(n1907), .Q(\u_cordic/mycordic/n540 )
         );
  INV3 U2668 ( .A(\u_cordic/mycordic/n473 ), .Q(n1535) );
  AOI221 U2669 ( .A(\u_cordic/mycordic/N470 ), .B(n777), .C(
        \u_cordic/mycordic/N498 ), .D(n1907), .Q(\u_cordic/mycordic/n473 ) );
  XNR21 U2670 ( .A(\u_cordic/mycordic/present_ANGLE_table[3][14] ), .B(
        \u_cordic/mycordic/sub_218/carry[14] ), .Q(\u_cordic/mycordic/N498 )
         );
  XOR21 U2671 ( .A(\u_cordic/mycordic/present_ANGLE_table[3][14] ), .B(
        \u_cordic/mycordic/add_213/carry[14] ), .Q(\u_cordic/mycordic/N470 )
         );
  INV3 U2672 ( .A(\u_coder/n300 ), .Q(n1939) );
  AOI221 U2673 ( .A(\u_coder/i [3]), .B(n894), .C(n2156), .D(\u_coder/N710 ), 
        .Q(\u_coder/n300 ) );
  INV3 U2674 ( .A(\u_coder/n277 ), .Q(n1920) );
  AOI221 U2675 ( .A(\u_coder/n263 ), .B(\u_coder/j [4]), .C(n2169), .D(
        \u_coder/N1017 ), .Q(\u_coder/n277 ) );
  INV3 U2676 ( .A(\u_coder/n276 ), .Q(n1921) );
  AOI221 U2677 ( .A(n890), .B(\u_coder/j [5]), .C(n2169), .D(\u_coder/N1018 ), 
        .Q(\u_coder/n276 ) );
  INV3 U2678 ( .A(\u_decoder/fir_filter/n628 ), .Q(n2464) );
  AOI221 U2679 ( .A(\u_decoder/fir_filter/Q_data_add_4 [7]), .B(n1087), .C(
        \u_decoder/fir_filter/Q_data_add_4_buff [7]), .D(n1162), .Q(
        \u_decoder/fir_filter/n628 ) );
  INV3 U2680 ( .A(\u_decoder/fir_filter/n626 ), .Q(n2462) );
  AOI221 U2681 ( .A(\u_decoder/fir_filter/Q_data_add_4 [9]), .B(n1087), .C(
        \u_decoder/fir_filter/Q_data_add_4_buff [9]), .D(n1162), .Q(
        \u_decoder/fir_filter/n626 ) );
  INV3 U2682 ( .A(\u_decoder/fir_filter/n926 ), .Q(n2584) );
  AOI221 U2683 ( .A(\u_decoder/fir_filter/I_data_add_4 [7]), .B(n1094), .C(
        \u_decoder/fir_filter/I_data_add_4_buff [7]), .D(n1157), .Q(
        \u_decoder/fir_filter/n926 ) );
  INV3 U2684 ( .A(\u_decoder/fir_filter/n924 ), .Q(n2582) );
  AOI221 U2685 ( .A(\u_decoder/fir_filter/I_data_add_4 [9]), .B(n1094), .C(
        \u_decoder/fir_filter/I_data_add_4_buff [9]), .D(n1159), .Q(
        \u_decoder/fir_filter/n924 ) );
  INV3 U2686 ( .A(\u_cordic/mycordic/n440 ), .Q(n1450) );
  AOI221 U2687 ( .A(\u_cordic/mycordic/N547 ), .B(n771), .C(
        \u_cordic/mycordic/N563 ), .D(n1903), .Q(\u_cordic/mycordic/n440 ) );
  XNR21 U2688 ( .A(\u_cordic/mycordic/present_ANGLE_table[5][13] ), .B(
        \u_cordic/mycordic/sub_236/carry [13]), .Q(\u_cordic/mycordic/N563 )
         );
  XOR21 U2689 ( .A(\u_cordic/mycordic/present_ANGLE_table[5][13] ), .B(
        \u_cordic/mycordic/add_233/carry [13]), .Q(\u_cordic/mycordic/N547 )
         );
  INV3 U2690 ( .A(\u_cordic/mycordic/n439 ), .Q(n1451) );
  AOI221 U2691 ( .A(\u_cordic/mycordic/N548 ), .B(n770), .C(
        \u_cordic/mycordic/N564 ), .D(n1903), .Q(\u_cordic/mycordic/n439 ) );
  XNR21 U2692 ( .A(\u_cordic/mycordic/present_ANGLE_table[5][14] ), .B(
        \u_cordic/mycordic/sub_236/carry [14]), .Q(\u_cordic/mycordic/N564 )
         );
  XOR21 U2693 ( .A(\u_cordic/mycordic/present_ANGLE_table[5][14] ), .B(
        \u_cordic/mycordic/add_233/carry [14]), .Q(\u_cordic/mycordic/N548 )
         );
  INV3 U2694 ( .A(\u_cordic/mycordic/n437 ), .Q(n1452) );
  AOI221 U2695 ( .A(\u_cordic/mycordic/N549 ), .B(n771), .C(
        \u_cordic/mycordic/N565 ), .D(n1903), .Q(\u_cordic/mycordic/n437 ) );
  XNR21 U2696 ( .A(\u_cordic/mycordic/sub_236/carry [15]), .B(
        \u_cordic/mycordic/present_ANGLE_table[5][15] ), .Q(
        \u_cordic/mycordic/N565 ) );
  XOR21 U2697 ( .A(\u_cordic/mycordic/add_233/carry [15]), .B(
        \u_cordic/mycordic/present_ANGLE_table[5][15] ), .Q(
        \u_cordic/mycordic/N549 ) );
  INV3 U2698 ( .A(n3037), .Q(n2654) );
  AOI211 U2699 ( .A(n3036), .B(\u_cordic/mycordic/present_I_table[4][3] ), .C(
        n2655), .Q(n3037) );
  INV3 U2700 ( .A(n3035), .Q(n2655) );
  INV3 U2701 ( .A(\u_coder/n302 ), .Q(n1937) );
  AOI221 U2702 ( .A(\u_coder/i [1]), .B(n893), .C(n2156), .D(\u_coder/N708 ), 
        .Q(\u_coder/n302 ) );
  INV3 U2703 ( .A(\u_cordic/mycordic/n538 ), .Q(n1496) );
  AOI221 U2704 ( .A(\u_cordic/mycordic/N500 ), .B(n776), .C(
        \u_cordic/mycordic/N517 ), .D(n1906), .Q(\u_cordic/mycordic/n538 ) );
  INV3 U2705 ( .A(\u_coder/n301 ), .Q(n1938) );
  AOI221 U2706 ( .A(\u_coder/i [2]), .B(n894), .C(n2156), .D(\u_coder/N709 ), 
        .Q(\u_coder/n301 ) );
  INV3 U2707 ( .A(n3024), .Q(n2640) );
  AOI211 U2708 ( .A(n286), .B(n3025), .C(
        \u_cordic/mycordic/present_I_table[5][7] ), .Q(n3024) );
  AOI211 U2709 ( .A(n3023), .B(\u_cordic/mycordic/present_Q_table[5][5] ), .C(
        n2643), .Q(n3025) );
  INV3 U2710 ( .A(n2693), .Q(n2147) );
  AOI211 U2711 ( .A(n126), .B(n2695), .C(\u_inFIFO/outWriteCount[1] ), .Q(
        n2693) );
  XNR21 U2712 ( .A(\u_cordic/mycordic/r173/carry [14]), .B(
        \u_cordic/mycordic/present_ANGLE_table[6][14] ), .Q(n374) );
  INV3 U2713 ( .A(\u_coder/n234 ), .Q(n1813) );
  OAI2111 U2714 ( .A(\u_coder/n213 ), .B(\u_coder/stateQ[0] ), .C(
        \u_coder/n235 ), .D(\u_coder/n236 ), .Q(\u_coder/n234 ) );
  NOR21 U2715 ( .A(n387), .B(n305), .Q(\u_cordic/mycordic/add_262/carry [5])
         );
  AOI211 U2716 ( .A(\u_outFIFO/n1145 ), .B(\u_outFIFO/n1146 ), .C(n1233), .Q(
        \u_outFIFO/N50 ) );
  AOI221 U2717 ( .A(n2218), .B(\u_outFIFO/currentState [1]), .C(n2224), .D(
        \u_outFIFO/n1147 ), .Q(\u_outFIFO/n1146 ) );
  AOI221 U2718 ( .A(\u_outFIFO/N1269 ), .B(\u_outFIFO/n1148 ), .C(
        \u_outFIFO/N1270 ), .D(\u_outFIFO/n1149 ), .Q(\u_outFIFO/n1145 ) );
  NOR21 U2719 ( .A(n297), .B(n97), .Q(\u_cordic/mycordic/sub_196/carry[2] ) );
  NOR21 U2720 ( .A(n402), .B(n98), .Q(\u_cordic/mycordic/add_191/carry[3] ) );
  NOR21 U2721 ( .A(n509), .B(n142), .Q(\u_cordic/mycordic/sub_196/carry[5] )
         );
  INV3 U2722 ( .A(\u_cordic/mycordic/sub_196/carry[4] ), .Q(n509) );
  NOR21 U2723 ( .A(n520), .B(n143), .Q(\u_cordic/mycordic/sub_207/carry [4])
         );
  INV3 U2724 ( .A(\u_cordic/mycordic/sub_207/carry [3]), .Q(n520) );
  NOR21 U2725 ( .A(n532), .B(n144), .Q(\u_cordic/mycordic/sub_218/carry[3] )
         );
  INV3 U2726 ( .A(\u_cordic/mycordic/sub_218/carry[2] ), .Q(n532) );
  NOR21 U2727 ( .A(n299), .B(n99), .Q(\u_cordic/mycordic/sub_229/carry[2] ) );
  NOR21 U2728 ( .A(n305), .B(n96), .Q(\u_cordic/mycordic/r173/carry [4]) );
  XOR21 U2729 ( .A(\u_cordic/mycordic/present_ANGLE_table[6][15] ), .B(
        \u_cordic/mycordic/add_262/carry [15]), .Q(\u_cordic/mycordic/N630 )
         );
  NOR21 U2730 ( .A(n268), .B(n561), .Q(\u_cordic/mycordic/add_262/carry [15])
         );
  XOR21 U2731 ( .A(\u_cordic/mycordic/add_262/carry [14]), .B(
        \u_cordic/mycordic/present_ANGLE_table[6][14] ), .Q(
        \u_cordic/mycordic/N629 ) );
  NOR21 U2732 ( .A(n389), .B(n475), .Q(\u_cordic/mycordic/add_262/carry [8])
         );
  NOR21 U2733 ( .A(n174), .B(n230), .Q(\u_cordic/mycordic/add_200/carry [1])
         );
  NOR21 U2734 ( .A(n176), .B(n231), .Q(\u_cordic/mycordic/add_206/carry [1])
         );
  NOR21 U2735 ( .A(n173), .B(n232), .Q(\u_cordic/mycordic/add_189/carry [1])
         );
  NOR21 U2736 ( .A(n175), .B(n233), .Q(\u_cordic/mycordic/add_195/carry [1])
         );
  NOR21 U2737 ( .A(n163), .B(n234), .Q(\u_cordic/mycordic/add_217/carry [1])
         );
  INV3 U2738 ( .A(n478), .Q(\u_outFIFO/r98/carry [1]) );
  NOR21 U2739 ( .A(n130), .B(\u_outFIFO/outWriteCount[0] ), .Q(n478) );
  NOR21 U2740 ( .A(n411), .B(n145), .Q(\u_cordic/mycordic/sub_196/carry[4] )
         );
  NOR21 U2741 ( .A(n404), .B(n146), .Q(\u_cordic/mycordic/add_191/carry[6] )
         );
  NOR21 U2742 ( .A(n500), .B(n147), .Q(\u_cordic/mycordic/add_191/carry[7] )
         );
  INV3 U2743 ( .A(\u_cordic/mycordic/add_191/carry[6] ), .Q(n500) );
  NOR21 U2744 ( .A(n501), .B(n183), .Q(\u_cordic/mycordic/add_191/carry[8] )
         );
  INV3 U2745 ( .A(\u_cordic/mycordic/add_191/carry[7] ), .Q(n501) );
  NOR21 U2746 ( .A(n502), .B(n184), .Q(\u_cordic/mycordic/add_191/carry[9] )
         );
  INV3 U2747 ( .A(\u_cordic/mycordic/add_191/carry[8] ), .Q(n502) );
  NOR21 U2748 ( .A(n503), .B(n235), .Q(\u_cordic/mycordic/add_191/carry[10] )
         );
  INV3 U2749 ( .A(\u_cordic/mycordic/add_191/carry[9] ), .Q(n503) );
  NOR21 U2750 ( .A(n504), .B(n236), .Q(\u_cordic/mycordic/add_191/carry[11] )
         );
  INV3 U2751 ( .A(\u_cordic/mycordic/add_191/carry[10] ), .Q(n504) );
  NOR21 U2752 ( .A(n505), .B(n269), .Q(\u_cordic/mycordic/add_191/carry[12] )
         );
  INV3 U2753 ( .A(\u_cordic/mycordic/add_191/carry[11] ), .Q(n505) );
  NOR21 U2754 ( .A(n506), .B(n270), .Q(\u_cordic/mycordic/add_191/carry[13] )
         );
  INV3 U2755 ( .A(\u_cordic/mycordic/add_191/carry[12] ), .Q(n506) );
  NOR21 U2756 ( .A(n507), .B(n271), .Q(\u_cordic/mycordic/add_191/carry[14] )
         );
  INV3 U2757 ( .A(\u_cordic/mycordic/add_191/carry[13] ), .Q(n507) );
  NOR21 U2758 ( .A(n298), .B(n148), .Q(\u_cordic/mycordic/sub_207/carry [3])
         );
  NOR21 U2759 ( .A(n419), .B(n149), .Q(\u_cordic/mycordic/add_202/carry [5])
         );
  NOR21 U2760 ( .A(n510), .B(n150), .Q(\u_cordic/mycordic/add_202/carry [6])
         );
  INV3 U2761 ( .A(\u_cordic/mycordic/add_202/carry [5]), .Q(n510) );
  NOR21 U2762 ( .A(n511), .B(n151), .Q(\u_cordic/mycordic/add_202/carry [7])
         );
  INV3 U2763 ( .A(\u_cordic/mycordic/add_202/carry [6]), .Q(n511) );
  NOR21 U2764 ( .A(n512), .B(n185), .Q(\u_cordic/mycordic/add_202/carry [8])
         );
  INV3 U2765 ( .A(\u_cordic/mycordic/add_202/carry [7]), .Q(n512) );
  NOR21 U2766 ( .A(n513), .B(n186), .Q(\u_cordic/mycordic/add_202/carry [9])
         );
  INV3 U2767 ( .A(\u_cordic/mycordic/add_202/carry [8]), .Q(n513) );
  NOR21 U2768 ( .A(n514), .B(n237), .Q(\u_cordic/mycordic/add_202/carry [10])
         );
  INV3 U2769 ( .A(\u_cordic/mycordic/add_202/carry [9]), .Q(n514) );
  NOR21 U2770 ( .A(n515), .B(n238), .Q(\u_cordic/mycordic/add_202/carry [11])
         );
  INV3 U2771 ( .A(\u_cordic/mycordic/add_202/carry [10]), .Q(n515) );
  NOR21 U2772 ( .A(n516), .B(n272), .Q(\u_cordic/mycordic/add_202/carry [12])
         );
  INV3 U2773 ( .A(\u_cordic/mycordic/add_202/carry [11]), .Q(n516) );
  NOR21 U2774 ( .A(n517), .B(n273), .Q(\u_cordic/mycordic/add_202/carry [13])
         );
  INV3 U2775 ( .A(\u_cordic/mycordic/add_202/carry [12]), .Q(n517) );
  NOR21 U2776 ( .A(n518), .B(n274), .Q(\u_cordic/mycordic/add_202/carry [14])
         );
  INV3 U2777 ( .A(\u_cordic/mycordic/add_202/carry [13]), .Q(n518) );
  NOR21 U2778 ( .A(n295), .B(n100), .Q(\u_cordic/mycordic/sub_218/carry[2] )
         );
  NOR21 U2779 ( .A(n434), .B(n101), .Q(\u_cordic/mycordic/add_213/carry[4] )
         );
  NOR21 U2780 ( .A(n521), .B(n152), .Q(\u_cordic/mycordic/add_213/carry[5] )
         );
  INV3 U2781 ( .A(\u_cordic/mycordic/add_213/carry[4] ), .Q(n521) );
  NOR21 U2782 ( .A(n522), .B(n153), .Q(\u_cordic/mycordic/add_213/carry[6] )
         );
  INV3 U2783 ( .A(\u_cordic/mycordic/add_213/carry[5] ), .Q(n522) );
  NOR21 U2784 ( .A(n523), .B(n154), .Q(\u_cordic/mycordic/add_213/carry[7] )
         );
  INV3 U2785 ( .A(\u_cordic/mycordic/add_213/carry[6] ), .Q(n523) );
  NOR21 U2786 ( .A(n524), .B(n187), .Q(\u_cordic/mycordic/add_213/carry[8] )
         );
  INV3 U2787 ( .A(\u_cordic/mycordic/add_213/carry[7] ), .Q(n524) );
  NOR21 U2788 ( .A(n525), .B(n188), .Q(\u_cordic/mycordic/add_213/carry[9] )
         );
  INV3 U2789 ( .A(\u_cordic/mycordic/add_213/carry[8] ), .Q(n525) );
  NOR21 U2790 ( .A(n526), .B(n239), .Q(\u_cordic/mycordic/add_213/carry[10] )
         );
  INV3 U2791 ( .A(\u_cordic/mycordic/add_213/carry[9] ), .Q(n526) );
  NOR21 U2792 ( .A(n527), .B(n240), .Q(\u_cordic/mycordic/add_213/carry[11] )
         );
  INV3 U2793 ( .A(\u_cordic/mycordic/add_213/carry[10] ), .Q(n527) );
  NOR21 U2794 ( .A(n528), .B(n275), .Q(\u_cordic/mycordic/add_213/carry[12] )
         );
  INV3 U2795 ( .A(\u_cordic/mycordic/add_213/carry[11] ), .Q(n528) );
  NOR21 U2796 ( .A(n529), .B(n276), .Q(\u_cordic/mycordic/add_213/carry[13] )
         );
  INV3 U2797 ( .A(\u_cordic/mycordic/add_213/carry[12] ), .Q(n529) );
  NOR21 U2798 ( .A(n530), .B(n277), .Q(\u_cordic/mycordic/add_213/carry[14] )
         );
  INV3 U2799 ( .A(\u_cordic/mycordic/add_213/carry[13] ), .Q(n530) );
  NOR21 U2800 ( .A(n447), .B(n102), .Q(\u_cordic/mycordic/add_224/carry[3] )
         );
  NOR21 U2801 ( .A(n533), .B(n103), .Q(\u_cordic/mycordic/add_224/carry[4] )
         );
  INV3 U2802 ( .A(\u_cordic/mycordic/add_224/carry[3] ), .Q(n533) );
  NOR21 U2803 ( .A(n534), .B(n155), .Q(\u_cordic/mycordic/add_224/carry[5] )
         );
  INV3 U2804 ( .A(\u_cordic/mycordic/add_224/carry[4] ), .Q(n534) );
  NOR21 U2805 ( .A(n535), .B(n156), .Q(\u_cordic/mycordic/add_224/carry[6] )
         );
  INV3 U2806 ( .A(\u_cordic/mycordic/add_224/carry[5] ), .Q(n535) );
  NOR21 U2807 ( .A(n536), .B(n157), .Q(\u_cordic/mycordic/add_224/carry[7] )
         );
  INV3 U2808 ( .A(\u_cordic/mycordic/add_224/carry[6] ), .Q(n536) );
  NOR21 U2809 ( .A(n537), .B(n189), .Q(\u_cordic/mycordic/add_224/carry[8] )
         );
  INV3 U2810 ( .A(\u_cordic/mycordic/add_224/carry[7] ), .Q(n537) );
  NOR21 U2811 ( .A(n538), .B(n190), .Q(\u_cordic/mycordic/add_224/carry[9] )
         );
  INV3 U2812 ( .A(\u_cordic/mycordic/add_224/carry[8] ), .Q(n538) );
  NOR21 U2813 ( .A(n539), .B(n241), .Q(\u_cordic/mycordic/add_224/carry[10] )
         );
  INV3 U2814 ( .A(\u_cordic/mycordic/add_224/carry[9] ), .Q(n539) );
  NOR21 U2815 ( .A(n540), .B(n242), .Q(\u_cordic/mycordic/add_224/carry[11] )
         );
  INV3 U2816 ( .A(\u_cordic/mycordic/add_224/carry[10] ), .Q(n540) );
  NOR21 U2817 ( .A(n541), .B(n278), .Q(\u_cordic/mycordic/add_224/carry[12] )
         );
  INV3 U2818 ( .A(\u_cordic/mycordic/add_224/carry[11] ), .Q(n541) );
  NOR21 U2819 ( .A(n542), .B(n279), .Q(\u_cordic/mycordic/add_224/carry[13] )
         );
  INV3 U2820 ( .A(\u_cordic/mycordic/add_224/carry[12] ), .Q(n542) );
  NOR21 U2821 ( .A(n543), .B(n280), .Q(\u_cordic/mycordic/add_224/carry[14] )
         );
  INV3 U2822 ( .A(\u_cordic/mycordic/add_224/carry[13] ), .Q(n543) );
  NOR21 U2823 ( .A(n296), .B(n104), .Q(\u_cordic/mycordic/add_233/carry [3])
         );
  NOR21 U2824 ( .A(n545), .B(n105), .Q(\u_cordic/mycordic/add_233/carry [4])
         );
  INV3 U2825 ( .A(\u_cordic/mycordic/add_233/carry [3]), .Q(n545) );
  NOR21 U2826 ( .A(n546), .B(n158), .Q(\u_cordic/mycordic/add_233/carry [5])
         );
  INV3 U2827 ( .A(\u_cordic/mycordic/add_233/carry [4]), .Q(n546) );
  NOR21 U2828 ( .A(n547), .B(n159), .Q(\u_cordic/mycordic/add_233/carry [6])
         );
  INV3 U2829 ( .A(\u_cordic/mycordic/add_233/carry [5]), .Q(n547) );
  NOR21 U2830 ( .A(n548), .B(n160), .Q(\u_cordic/mycordic/add_233/carry [7])
         );
  INV3 U2831 ( .A(\u_cordic/mycordic/add_233/carry [6]), .Q(n548) );
  NOR21 U2832 ( .A(n549), .B(n191), .Q(\u_cordic/mycordic/add_233/carry [8])
         );
  INV3 U2833 ( .A(\u_cordic/mycordic/add_233/carry [7]), .Q(n549) );
  NOR21 U2834 ( .A(n550), .B(n192), .Q(\u_cordic/mycordic/add_233/carry [9])
         );
  INV3 U2835 ( .A(\u_cordic/mycordic/add_233/carry [8]), .Q(n550) );
  NOR21 U2836 ( .A(n551), .B(n243), .Q(\u_cordic/mycordic/add_233/carry [10])
         );
  INV3 U2837 ( .A(\u_cordic/mycordic/add_233/carry [9]), .Q(n551) );
  NOR21 U2838 ( .A(n552), .B(n244), .Q(\u_cordic/mycordic/add_233/carry [11])
         );
  INV3 U2839 ( .A(\u_cordic/mycordic/add_233/carry [10]), .Q(n552) );
  NOR21 U2840 ( .A(n553), .B(n281), .Q(\u_cordic/mycordic/add_233/carry [12])
         );
  INV3 U2841 ( .A(\u_cordic/mycordic/add_233/carry [11]), .Q(n553) );
  NOR21 U2842 ( .A(n554), .B(n282), .Q(\u_cordic/mycordic/add_233/carry [13])
         );
  INV3 U2843 ( .A(\u_cordic/mycordic/add_233/carry [12]), .Q(n554) );
  NOR21 U2844 ( .A(n555), .B(n283), .Q(\u_cordic/mycordic/add_233/carry [14])
         );
  INV3 U2845 ( .A(\u_cordic/mycordic/add_233/carry [13]), .Q(n555) );
  AOI221 U2846 ( .A(\u_outFIFO/N126 ), .B(n1912), .C(\u_outFIFO/N150 ), .D(
        \u_outFIFO/n1131 ), .Q(\u_outFIFO/n1138 ) );
  XOR21 U2847 ( .A(\u_outFIFO/add_255/carry [7]), .B(
        \u_outFIFO/outWriteCount[7] ), .Q(\u_outFIFO/N126 ) );
  AOI211 U2848 ( .A(\u_coder/n246 ), .B(\u_coder/n126 ), .C(\u_coder/n247 ), 
        .Q(\u_coder/n243 ) );
  NAND22 U2849 ( .A(sig_coder_outSinIMasked[3]), .B(\u_coder/n245 ), .Q(
        \u_coder/n244 ) );
  INV3 U2850 ( .A(\u_cordic/mycordic/n507 ), .Q(n1465) );
  AOI221 U2851 ( .A(\u_cordic/mycordic/N344 ), .B(n772), .C(
        \u_cordic/mycordic/N376 ), .D(n1904), .Q(\u_cordic/mycordic/n507 ) );
  XNR21 U2852 ( .A(\u_cordic/mycordic/present_ANGLE_table[1][12] ), .B(
        \u_cordic/mycordic/sub_196/carry[12] ), .Q(\u_cordic/mycordic/N376 )
         );
  XOR21 U2853 ( .A(\u_cordic/mycordic/present_ANGLE_table[1][12] ), .B(
        \u_cordic/mycordic/add_191/carry[12] ), .Q(\u_cordic/mycordic/N344 )
         );
  INV3 U2854 ( .A(\u_cordic/mycordic/n475 ), .Q(n1533) );
  AOI221 U2855 ( .A(\u_cordic/mycordic/N468 ), .B(n777), .C(
        \u_cordic/mycordic/N496 ), .D(n1907), .Q(\u_cordic/mycordic/n475 ) );
  XNR21 U2856 ( .A(\u_cordic/mycordic/present_ANGLE_table[3][12] ), .B(
        \u_cordic/mycordic/sub_218/carry[12] ), .Q(\u_cordic/mycordic/N496 )
         );
  XOR21 U2857 ( .A(\u_cordic/mycordic/present_ANGLE_table[3][12] ), .B(
        \u_cordic/mycordic/add_213/carry[12] ), .Q(\u_cordic/mycordic/N468 )
         );
  AOI221 U2858 ( .A(\u_inFIFO/N149 ), .B(\u_inFIFO/n533 ), .C(\u_inFIFO/N140 ), 
        .D(\u_inFIFO/n534 ), .Q(\u_inFIFO/n548 ) );
  XOR21 U2859 ( .A(\u_inFIFO/add_263/carry [7]), .B(
        \u_inFIFO/outWriteCount[7] ), .Q(\u_inFIFO/N149 ) );
  AOI211 U2860 ( .A(n2174), .B(\u_coder/n127 ), .C(\u_coder/n228 ), .Q(
        \u_coder/n226 ) );
  NAND22 U2861 ( .A(sig_coder_outSinQMasked[3]), .B(n1813), .Q(\u_coder/n227 )
         );
  NAND22 U2862 ( .A(\u_inFIFO/outReadCount[3] ), .B(\u_inFIFO/n185 ), .Q(n2697) );
  AOI221 U2863 ( .A(\u_coder/n137 ), .B(n2104), .C(n2168), .D(\u_coder/n138 ), 
        .Q(\u_coder/n136 ) );
  INV3 U2864 ( .A(\u_coder/n139 ), .Q(n2104) );
  NAND22 U2865 ( .A(\u_decoder/fir_filter/I_data_mult_3_buff [9]), .B(n1158), 
        .Q(\u_decoder/fir_filter/n1095 ) );
  NAND22 U2866 ( .A(\u_decoder/fir_filter/I_data_mult_5_buff [9]), .B(n1164), 
        .Q(\u_decoder/fir_filter/n1063 ) );
  NAND22 U2867 ( .A(\u_decoder/fir_filter/Q_data_mult_3_buff [9]), .B(n1151), 
        .Q(\u_decoder/fir_filter/n798 ) );
  NAND22 U2868 ( .A(\u_decoder/fir_filter/Q_data_mult_5_buff [9]), .B(n1155), 
        .Q(\u_decoder/fir_filter/n766 ) );
  NAND22 U2869 ( .A(\u_decoder/fir_filter/I_data_mult_2_buff [8]), .B(n1159), 
        .Q(\u_decoder/fir_filter/n1110 ) );
  NAND22 U2870 ( .A(\u_decoder/fir_filter/I_data_mult_6_buff [8]), .B(n1157), 
        .Q(\u_decoder/fir_filter/n1045 ) );
  NAND22 U2871 ( .A(\u_decoder/fir_filter/Q_data_mult_2_buff [8]), .B(n1159), 
        .Q(\u_decoder/fir_filter/n813 ) );
  NAND22 U2872 ( .A(\u_decoder/fir_filter/Q_data_mult_6_buff [8]), .B(n1155), 
        .Q(\u_decoder/fir_filter/n748 ) );
  NAND22 U2873 ( .A(\u_decoder/fir_filter/I_data_mult_2_buff [7]), .B(n1159), 
        .Q(\u_decoder/fir_filter/n1109 ) );
  NAND22 U2874 ( .A(\u_decoder/fir_filter/I_data_mult_3_buff [7]), .B(n1159), 
        .Q(\u_decoder/fir_filter/n1093 ) );
  NAND22 U2875 ( .A(\u_decoder/fir_filter/I_data_mult_5_buff [7]), .B(n1165), 
        .Q(\u_decoder/fir_filter/n1061 ) );
  NAND22 U2876 ( .A(\u_decoder/fir_filter/I_data_mult_6_buff [7]), .B(n1157), 
        .Q(\u_decoder/fir_filter/n1044 ) );
  NAND22 U2877 ( .A(\u_decoder/fir_filter/Q_data_mult_2_buff [7]), .B(n1159), 
        .Q(\u_decoder/fir_filter/n812 ) );
  NAND22 U2878 ( .A(\u_decoder/fir_filter/Q_data_mult_3_buff [7]), .B(n1162), 
        .Q(\u_decoder/fir_filter/n796 ) );
  NAND22 U2879 ( .A(\u_decoder/fir_filter/Q_data_mult_5_buff [7]), .B(n1155), 
        .Q(\u_decoder/fir_filter/n764 ) );
  NAND22 U2880 ( .A(\u_decoder/fir_filter/Q_data_mult_6_buff [7]), .B(n1154), 
        .Q(\u_decoder/fir_filter/n747 ) );
  NAND22 U2881 ( .A(\u_decoder/fir_filter/I_data_mult_3_buff [8]), .B(n1158), 
        .Q(\u_decoder/fir_filter/n1094 ) );
  NAND22 U2882 ( .A(\u_decoder/fir_filter/I_data_mult_5_buff [8]), .B(n1154), 
        .Q(\u_decoder/fir_filter/n1062 ) );
  NAND22 U2883 ( .A(\u_decoder/fir_filter/Q_data_mult_3_buff [8]), .B(n1161), 
        .Q(\u_decoder/fir_filter/n797 ) );
  NAND22 U2884 ( .A(\u_decoder/fir_filter/Q_data_mult_5_buff [8]), .B(n1155), 
        .Q(\u_decoder/fir_filter/n765 ) );
  NAND22 U2885 ( .A(\u_decoder/fir_filter/I_data_mult_1_buff [8]), .B(n1160), 
        .Q(\u_decoder/fir_filter/n1126 ) );
  NAND22 U2886 ( .A(\u_decoder/fir_filter/I_data_mult_7_buff [8]), .B(n1156), 
        .Q(\u_decoder/fir_filter/n1028 ) );
  NAND22 U2887 ( .A(\u_decoder/fir_filter/Q_data_mult_1_buff [8]), .B(n1152), 
        .Q(\u_decoder/fir_filter/n829 ) );
  NAND22 U2888 ( .A(\u_decoder/fir_filter/Q_data_mult_7_buff [8]), .B(n1154), 
        .Q(\u_decoder/fir_filter/n731 ) );
  NAND22 U2889 ( .A(\u_inFIFO/outReadCount[2] ), .B(\u_inFIFO/n186 ), .Q(n2694) );
  NAND22 U2890 ( .A(\u_decoder/fir_filter/I_data_mult_0_buff [7]), .B(n1153), 
        .Q(\u_decoder/fir_filter/n1141 ) );
  NAND22 U2891 ( .A(\u_decoder/fir_filter/Q_data_mult_0_buff [7]), .B(n1151), 
        .Q(\u_decoder/fir_filter/n844 ) );
  NOR21 U2892 ( .A(\u_inFIFO/n188 ), .B(\u_inFIFO/outReadCount[0] ), .Q(n2695)
         );
  INV3 U2893 ( .A(\u_cordic/mycordic/n400 ), .Q(n1869) );
  NAND22 U2894 ( .A(\u_cordic/mycordic/next_ANGLE_table[6][14] ), .B(n1215), 
        .Q(\u_cordic/mycordic/n400 ) );
  NAND22 U2895 ( .A(\u_inFIFO/outReadCount[4] ), .B(\u_inFIFO/n184 ), .Q(n2698) );
  NOR21 U2896 ( .A(n179), .B(\u_cordic/mycordic/present_I_table[4][0] ), .Q(
        n3027) );
  AOI211 U2897 ( .A(\u_inFIFO/n558 ), .B(\u_inFIFO/n559 ), .C(n1240), .Q(
        \u_inFIFO/N50 ) );
  NAND22 U2898 ( .A(n2145), .B(\u_inFIFO/n560 ), .Q(\u_inFIFO/n559 ) );
  AOI221 U2899 ( .A(\u_inFIFO/currentState [0]), .B(\u_inFIFO/n215 ), .C(
        \u_inFIFO/N375 ), .D(\u_inFIFO/n561 ), .Q(\u_inFIFO/n558 ) );
  INV3 U2900 ( .A(n2711), .Q(n2145) );
  INV3 U2901 ( .A(n399), .Q(\u_cordic/mycordic/r173/carry [6]) );
  NOR21 U2902 ( .A(\u_cordic/mycordic/present_ANGLE_table[6][5] ), .B(
        \u_cordic/mycordic/r173/carry [5]), .Q(n399) );
  INV3 U2903 ( .A(n474), .Q(\u_cordic/mycordic/add_262/carry [6]) );
  NOR21 U2904 ( .A(\u_cordic/mycordic/present_ANGLE_table[6][5] ), .B(
        \u_cordic/mycordic/add_262/carry [5]), .Q(n474) );
  NAND22 U2905 ( .A(\u_coder/n185 ), .B(\u_coder/n186 ), .Q(\u_coder/n337 ) );
  AOI221 U2906 ( .A(n2185), .B(\u_coder/n187 ), .C(n2102), .D(\u_coder/n188 ), 
        .Q(\u_coder/n185 ) );
  NAND22 U2907 ( .A(sig_coder_outSinQ[2]), .B(\u_coder/n179 ), .Q(
        \u_coder/n186 ) );
  NAND22 U2908 ( .A(\u_coder/n196 ), .B(\u_coder/n197 ), .Q(\u_coder/n338 ) );
  AOI221 U2909 ( .A(n2185), .B(\u_coder/n198 ), .C(n2102), .D(\u_coder/n199 ), 
        .Q(\u_coder/n196 ) );
  NAND22 U2910 ( .A(sig_coder_outSinQ[1]), .B(\u_coder/n179 ), .Q(
        \u_coder/n197 ) );
  INV3 U2911 ( .A(n475), .Q(\u_cordic/mycordic/add_262/carry [7]) );
  NOR21 U2912 ( .A(\u_cordic/mycordic/present_ANGLE_table[6][6] ), .B(
        \u_cordic/mycordic/add_262/carry [6]), .Q(n475) );
  INV3 U2913 ( .A(n400), .Q(\u_cordic/mycordic/r173/carry [8]) );
  NOR21 U2914 ( .A(\u_cordic/mycordic/present_ANGLE_table[6][7] ), .B(
        \u_cordic/mycordic/r173/carry [7]), .Q(n400) );
  INV3 U2915 ( .A(n476), .Q(\u_cordic/mycordic/add_262/carry [9]) );
  NOR21 U2916 ( .A(\u_cordic/mycordic/present_ANGLE_table[6][8] ), .B(
        \u_cordic/mycordic/add_262/carry [8]), .Q(n476) );
  INV3 U2917 ( .A(n402), .Q(\u_cordic/mycordic/add_191/carry[2] ) );
  NOR21 U2918 ( .A(\u_cordic/mycordic/present_ANGLE_table[1][0] ), .B(
        \u_cordic/mycordic/present_ANGLE_table[1][1] ), .Q(n402) );
  INV3 U2919 ( .A(n418), .Q(\u_cordic/mycordic/add_202/carry [3]) );
  NOR21 U2920 ( .A(\u_cordic/mycordic/present_ANGLE_table[2][1] ), .B(
        \u_cordic/mycordic/present_ANGLE_table[2][2] ), .Q(n418) );
  INV3 U2921 ( .A(n433), .Q(\u_cordic/mycordic/add_213/carry[2] ) );
  NOR21 U2922 ( .A(\u_cordic/mycordic/present_ANGLE_table[3][0] ), .B(
        \u_cordic/mycordic/present_ANGLE_table[3][1] ), .Q(n433) );
  INV3 U2923 ( .A(n447), .Q(\u_cordic/mycordic/add_224/carry[2] ) );
  NOR21 U2924 ( .A(\u_cordic/mycordic/present_ANGLE_table[4][0] ), .B(
        \u_cordic/mycordic/present_ANGLE_table[4][1] ), .Q(n447) );
  INV3 U2925 ( .A(n466), .Q(\u_cordic/mycordic/sub_236/carry [3]) );
  NOR21 U2926 ( .A(\u_cordic/mycordic/present_ANGLE_table[5][1] ), .B(
        \u_cordic/mycordic/present_ANGLE_table[5][2] ), .Q(n466) );
  NAND22 U2927 ( .A(\u_coder/n229 ), .B(\u_coder/n230 ), .Q(\u_coder/n342 ) );
  NAND22 U2928 ( .A(sig_coder_outSinQMasked[2]), .B(n1813), .Q(\u_coder/n230 )
         );
  NAND22 U2929 ( .A(\u_coder/n229 ), .B(\u_coder/n231 ), .Q(\u_coder/n343 ) );
  NAND22 U2930 ( .A(sig_coder_outSinQMasked[1]), .B(n1813), .Q(\u_coder/n231 )
         );
  INV3 U2931 ( .A(n479), .Q(\u_inFIFO/r96/carry [1]) );
  NOR21 U2932 ( .A(n129), .B(\u_inFIFO/outWriteCount[0] ), .Q(n479) );
  INV3 U2933 ( .A(\u_cordic/mycordic/n367 ), .Q(n1569) );
  AOI221 U2934 ( .A(\u_cordic/mycordic/N387 ), .B(n778), .C(
        \u_cordic/mycordic/N419 ), .D(n1908), .Q(\u_cordic/mycordic/n367 ) );
  INV3 U2935 ( .A(\u_cordic/mycordic/n375 ), .Q(n1476) );
  AOI221 U2936 ( .A(\u_cordic/mycordic/N323 ), .B(\u_cordic/mycordic/n336 ), 
        .C(\u_cordic/mycordic/N355 ), .D(n1904), .Q(\u_cordic/mycordic/n375 )
         );
  INV3 U2937 ( .A(n420), .Q(\u_cordic/mycordic/sub_205/carry [1]) );
  NOR21 U2938 ( .A(n174), .B(\u_cordic/mycordic/present_I_table[3][0] ), .Q(
        n420) );
  INV3 U2939 ( .A(n417), .Q(\u_cordic/mycordic/sub_201/carry [1]) );
  NOR21 U2940 ( .A(n176), .B(\u_cordic/mycordic/present_Q_table[3][0] ), .Q(
        n417) );
  INV3 U2941 ( .A(n405), .Q(\u_cordic/mycordic/sub_194/carry [1]) );
  NOR21 U2942 ( .A(n173), .B(\u_cordic/mycordic/present_I_table[2][0] ), .Q(
        n405) );
  INV3 U2943 ( .A(n401), .Q(\u_cordic/mycordic/sub_190/carry [1]) );
  NOR21 U2944 ( .A(n175), .B(\u_cordic/mycordic/present_Q_table[2][0] ), .Q(
        n401) );
  INV3 U2945 ( .A(n432), .Q(\u_cordic/mycordic/sub_212/carry [1]) );
  NOR21 U2946 ( .A(n163), .B(\u_cordic/mycordic/present_Q_table[4][0] ), .Q(
        n432) );
  INV3 U2947 ( .A(n411), .Q(\u_cordic/mycordic/sub_196/carry[3] ) );
  NOR21 U2948 ( .A(\u_cordic/mycordic/sub_196/carry[2] ), .B(
        \u_cordic/mycordic/present_ANGLE_table[1][2] ), .Q(n411) );
  INV3 U2949 ( .A(\u_cordic/mycordic/n401 ), .Q(n1870) );
  NAND22 U2950 ( .A(\u_cordic/mycordic/next_ANGLE_table[6][13] ), .B(n1215), 
        .Q(\u_cordic/mycordic/n401 ) );
  INV3 U2951 ( .A(n3014), .Q(n2650) );
  NOR21 U2952 ( .A(\u_cordic/mycordic/present_Q_table[5][1] ), .B(n3015), .Q(
        n3014) );
  INV3 U2953 ( .A(n398), .Q(\u_cordic/mycordic/r173/carry [5]) );
  NOR21 U2954 ( .A(\u_cordic/mycordic/present_ANGLE_table[6][4] ), .B(
        \u_cordic/mycordic/r173/carry [4]), .Q(n398) );
  NOR21 U2955 ( .A(n508), .B(n308), .Q(\u_cordic/mycordic/add_191/carry[15] )
         );
  INV3 U2956 ( .A(\u_cordic/mycordic/add_191/carry[14] ), .Q(n508) );
  NOR21 U2957 ( .A(n519), .B(n309), .Q(\u_cordic/mycordic/add_202/carry [15])
         );
  INV3 U2958 ( .A(\u_cordic/mycordic/add_202/carry [14]), .Q(n519) );
  NOR21 U2959 ( .A(n531), .B(n310), .Q(\u_cordic/mycordic/add_213/carry[15] )
         );
  INV3 U2960 ( .A(\u_cordic/mycordic/add_213/carry[14] ), .Q(n531) );
  NOR21 U2961 ( .A(n544), .B(n311), .Q(\u_cordic/mycordic/add_224/carry[15] )
         );
  INV3 U2962 ( .A(\u_cordic/mycordic/add_224/carry[14] ), .Q(n544) );
  NOR21 U2963 ( .A(n556), .B(n312), .Q(\u_cordic/mycordic/add_233/carry [15])
         );
  INV3 U2964 ( .A(\u_cordic/mycordic/add_233/carry [14]), .Q(n556) );
  INV3 U2965 ( .A(n403), .Q(\u_cordic/mycordic/add_191/carry[4] ) );
  NOR21 U2966 ( .A(\u_cordic/mycordic/add_191/carry[3] ), .B(
        \u_cordic/mycordic/present_ANGLE_table[1][3] ), .Q(n403) );
  INV3 U2967 ( .A(n412), .Q(\u_cordic/mycordic/sub_196/carry[6] ) );
  NOR21 U2968 ( .A(\u_cordic/mycordic/sub_196/carry[5] ), .B(
        \u_cordic/mycordic/present_ANGLE_table[1][5] ), .Q(n412) );
  INV3 U2969 ( .A(n413), .Q(\u_cordic/mycordic/sub_196/carry[7] ) );
  NOR21 U2970 ( .A(\u_cordic/mycordic/sub_196/carry[6] ), .B(
        \u_cordic/mycordic/present_ANGLE_table[1][6] ), .Q(n413) );
  INV3 U2971 ( .A(n414), .Q(\u_cordic/mycordic/sub_196/carry[8] ) );
  NOR21 U2972 ( .A(\u_cordic/mycordic/sub_196/carry[7] ), .B(
        \u_cordic/mycordic/present_ANGLE_table[1][7] ), .Q(n414) );
  INV3 U2973 ( .A(n415), .Q(\u_cordic/mycordic/sub_196/carry[9] ) );
  NOR21 U2974 ( .A(\u_cordic/mycordic/sub_196/carry[8] ), .B(
        \u_cordic/mycordic/present_ANGLE_table[1][8] ), .Q(n415) );
  INV3 U2975 ( .A(n416), .Q(\u_cordic/mycordic/sub_196/carry[10] ) );
  NOR21 U2976 ( .A(\u_cordic/mycordic/sub_196/carry[9] ), .B(
        \u_cordic/mycordic/present_ANGLE_table[1][9] ), .Q(n416) );
  INV3 U2977 ( .A(n406), .Q(\u_cordic/mycordic/sub_196/carry[11] ) );
  NOR21 U2978 ( .A(\u_cordic/mycordic/sub_196/carry[10] ), .B(
        \u_cordic/mycordic/present_ANGLE_table[1][10] ), .Q(n406) );
  INV3 U2979 ( .A(n407), .Q(\u_cordic/mycordic/sub_196/carry[12] ) );
  NOR21 U2980 ( .A(\u_cordic/mycordic/sub_196/carry[11] ), .B(
        \u_cordic/mycordic/present_ANGLE_table[1][11] ), .Q(n407) );
  INV3 U2981 ( .A(n408), .Q(\u_cordic/mycordic/sub_196/carry[13] ) );
  NOR21 U2982 ( .A(\u_cordic/mycordic/sub_196/carry[12] ), .B(
        \u_cordic/mycordic/present_ANGLE_table[1][12] ), .Q(n408) );
  INV3 U2983 ( .A(n409), .Q(\u_cordic/mycordic/sub_196/carry[14] ) );
  NOR21 U2984 ( .A(\u_cordic/mycordic/sub_196/carry[13] ), .B(
        \u_cordic/mycordic/present_ANGLE_table[1][13] ), .Q(n409) );
  INV3 U2985 ( .A(n426), .Q(\u_cordic/mycordic/sub_207/carry [5]) );
  NOR21 U2986 ( .A(\u_cordic/mycordic/sub_207/carry [4]), .B(
        \u_cordic/mycordic/present_ANGLE_table[2][4] ), .Q(n426) );
  INV3 U2987 ( .A(n427), .Q(\u_cordic/mycordic/sub_207/carry [6]) );
  NOR21 U2988 ( .A(\u_cordic/mycordic/sub_207/carry [5]), .B(
        \u_cordic/mycordic/present_ANGLE_table[2][5] ), .Q(n427) );
  INV3 U2989 ( .A(n428), .Q(\u_cordic/mycordic/sub_207/carry [7]) );
  NOR21 U2990 ( .A(\u_cordic/mycordic/sub_207/carry [6]), .B(
        \u_cordic/mycordic/present_ANGLE_table[2][6] ), .Q(n428) );
  INV3 U2991 ( .A(n429), .Q(\u_cordic/mycordic/sub_207/carry [8]) );
  NOR21 U2992 ( .A(\u_cordic/mycordic/sub_207/carry [7]), .B(
        \u_cordic/mycordic/present_ANGLE_table[2][7] ), .Q(n429) );
  INV3 U2993 ( .A(n430), .Q(\u_cordic/mycordic/sub_207/carry [9]) );
  NOR21 U2994 ( .A(\u_cordic/mycordic/sub_207/carry [8]), .B(
        \u_cordic/mycordic/present_ANGLE_table[2][8] ), .Q(n430) );
  INV3 U2995 ( .A(n431), .Q(\u_cordic/mycordic/sub_207/carry [10]) );
  NOR21 U2996 ( .A(\u_cordic/mycordic/sub_207/carry [9]), .B(
        \u_cordic/mycordic/present_ANGLE_table[2][9] ), .Q(n431) );
  INV3 U2997 ( .A(n421), .Q(\u_cordic/mycordic/sub_207/carry [11]) );
  NOR21 U2998 ( .A(\u_cordic/mycordic/sub_207/carry [10]), .B(
        \u_cordic/mycordic/present_ANGLE_table[2][10] ), .Q(n421) );
  INV3 U2999 ( .A(n422), .Q(\u_cordic/mycordic/sub_207/carry [12]) );
  NOR21 U3000 ( .A(\u_cordic/mycordic/sub_207/carry [11]), .B(
        \u_cordic/mycordic/present_ANGLE_table[2][11] ), .Q(n422) );
  INV3 U3001 ( .A(n423), .Q(\u_cordic/mycordic/sub_207/carry [13]) );
  NOR21 U3002 ( .A(\u_cordic/mycordic/sub_207/carry [12]), .B(
        \u_cordic/mycordic/present_ANGLE_table[2][12] ), .Q(n423) );
  INV3 U3003 ( .A(n424), .Q(\u_cordic/mycordic/sub_207/carry [14]) );
  NOR21 U3004 ( .A(\u_cordic/mycordic/sub_207/carry [13]), .B(
        \u_cordic/mycordic/present_ANGLE_table[2][13] ), .Q(n424) );
  INV3 U3005 ( .A(n440), .Q(\u_cordic/mycordic/sub_218/carry[4] ) );
  NOR21 U3006 ( .A(\u_cordic/mycordic/sub_218/carry[3] ), .B(
        \u_cordic/mycordic/present_ANGLE_table[3][3] ), .Q(n440) );
  INV3 U3007 ( .A(n441), .Q(\u_cordic/mycordic/sub_218/carry[5] ) );
  NOR21 U3008 ( .A(\u_cordic/mycordic/sub_218/carry[4] ), .B(
        \u_cordic/mycordic/present_ANGLE_table[3][4] ), .Q(n441) );
  INV3 U3009 ( .A(n442), .Q(\u_cordic/mycordic/sub_218/carry[6] ) );
  NOR21 U3010 ( .A(\u_cordic/mycordic/sub_218/carry[5] ), .B(
        \u_cordic/mycordic/present_ANGLE_table[3][5] ), .Q(n442) );
  INV3 U3011 ( .A(n443), .Q(\u_cordic/mycordic/sub_218/carry[7] ) );
  NOR21 U3012 ( .A(\u_cordic/mycordic/sub_218/carry[6] ), .B(
        \u_cordic/mycordic/present_ANGLE_table[3][6] ), .Q(n443) );
  INV3 U3013 ( .A(n444), .Q(\u_cordic/mycordic/sub_218/carry[8] ) );
  NOR21 U3014 ( .A(\u_cordic/mycordic/sub_218/carry[7] ), .B(
        \u_cordic/mycordic/present_ANGLE_table[3][7] ), .Q(n444) );
  INV3 U3015 ( .A(n445), .Q(\u_cordic/mycordic/sub_218/carry[9] ) );
  NOR21 U3016 ( .A(\u_cordic/mycordic/sub_218/carry[8] ), .B(
        \u_cordic/mycordic/present_ANGLE_table[3][8] ), .Q(n445) );
  INV3 U3017 ( .A(n446), .Q(\u_cordic/mycordic/sub_218/carry[10] ) );
  NOR21 U3018 ( .A(\u_cordic/mycordic/sub_218/carry[9] ), .B(
        \u_cordic/mycordic/present_ANGLE_table[3][9] ), .Q(n446) );
  INV3 U3019 ( .A(n435), .Q(\u_cordic/mycordic/sub_218/carry[11] ) );
  NOR21 U3020 ( .A(\u_cordic/mycordic/sub_218/carry[10] ), .B(
        \u_cordic/mycordic/present_ANGLE_table[3][10] ), .Q(n435) );
  INV3 U3021 ( .A(n436), .Q(\u_cordic/mycordic/sub_218/carry[12] ) );
  NOR21 U3022 ( .A(\u_cordic/mycordic/sub_218/carry[11] ), .B(
        \u_cordic/mycordic/present_ANGLE_table[3][11] ), .Q(n436) );
  INV3 U3023 ( .A(n437), .Q(\u_cordic/mycordic/sub_218/carry[13] ) );
  NOR21 U3024 ( .A(\u_cordic/mycordic/sub_218/carry[12] ), .B(
        \u_cordic/mycordic/present_ANGLE_table[3][12] ), .Q(n437) );
  INV3 U3025 ( .A(n438), .Q(\u_cordic/mycordic/sub_218/carry[14] ) );
  NOR21 U3026 ( .A(\u_cordic/mycordic/sub_218/carry[13] ), .B(
        \u_cordic/mycordic/present_ANGLE_table[3][13] ), .Q(n438) );
  INV3 U3027 ( .A(n453), .Q(\u_cordic/mycordic/sub_229/carry[3] ) );
  NOR21 U3028 ( .A(\u_cordic/mycordic/sub_229/carry[2] ), .B(
        \u_cordic/mycordic/present_ANGLE_table[4][2] ), .Q(n453) );
  INV3 U3029 ( .A(n454), .Q(\u_cordic/mycordic/sub_229/carry[4] ) );
  NOR21 U3030 ( .A(\u_cordic/mycordic/sub_229/carry[3] ), .B(
        \u_cordic/mycordic/present_ANGLE_table[4][3] ), .Q(n454) );
  INV3 U3031 ( .A(n455), .Q(\u_cordic/mycordic/sub_229/carry[5] ) );
  NOR21 U3032 ( .A(\u_cordic/mycordic/sub_229/carry[4] ), .B(
        \u_cordic/mycordic/present_ANGLE_table[4][4] ), .Q(n455) );
  INV3 U3033 ( .A(n456), .Q(\u_cordic/mycordic/sub_229/carry[6] ) );
  NOR21 U3034 ( .A(\u_cordic/mycordic/sub_229/carry[5] ), .B(
        \u_cordic/mycordic/present_ANGLE_table[4][5] ), .Q(n456) );
  INV3 U3035 ( .A(n457), .Q(\u_cordic/mycordic/sub_229/carry[7] ) );
  NOR21 U3036 ( .A(\u_cordic/mycordic/sub_229/carry[6] ), .B(
        \u_cordic/mycordic/present_ANGLE_table[4][6] ), .Q(n457) );
  INV3 U3037 ( .A(n458), .Q(\u_cordic/mycordic/sub_229/carry[8] ) );
  NOR21 U3038 ( .A(\u_cordic/mycordic/sub_229/carry[7] ), .B(
        \u_cordic/mycordic/present_ANGLE_table[4][7] ), .Q(n458) );
  INV3 U3039 ( .A(n459), .Q(\u_cordic/mycordic/sub_229/carry[9] ) );
  NOR21 U3040 ( .A(\u_cordic/mycordic/sub_229/carry[8] ), .B(
        \u_cordic/mycordic/present_ANGLE_table[4][8] ), .Q(n459) );
  INV3 U3041 ( .A(n460), .Q(\u_cordic/mycordic/sub_229/carry[10] ) );
  NOR21 U3042 ( .A(\u_cordic/mycordic/sub_229/carry[9] ), .B(
        \u_cordic/mycordic/present_ANGLE_table[4][9] ), .Q(n460) );
  INV3 U3043 ( .A(n448), .Q(\u_cordic/mycordic/sub_229/carry[11] ) );
  NOR21 U3044 ( .A(\u_cordic/mycordic/sub_229/carry[10] ), .B(
        \u_cordic/mycordic/present_ANGLE_table[4][10] ), .Q(n448) );
  INV3 U3045 ( .A(n449), .Q(\u_cordic/mycordic/sub_229/carry[12] ) );
  NOR21 U3046 ( .A(\u_cordic/mycordic/sub_229/carry[11] ), .B(
        \u_cordic/mycordic/present_ANGLE_table[4][11] ), .Q(n449) );
  INV3 U3047 ( .A(n450), .Q(\u_cordic/mycordic/sub_229/carry[13] ) );
  NOR21 U3048 ( .A(\u_cordic/mycordic/sub_229/carry[12] ), .B(
        \u_cordic/mycordic/present_ANGLE_table[4][12] ), .Q(n450) );
  INV3 U3049 ( .A(n451), .Q(\u_cordic/mycordic/sub_229/carry[14] ) );
  NOR21 U3050 ( .A(\u_cordic/mycordic/sub_229/carry[13] ), .B(
        \u_cordic/mycordic/present_ANGLE_table[4][13] ), .Q(n451) );
  INV3 U3051 ( .A(n467), .Q(\u_cordic/mycordic/sub_236/carry [4]) );
  NOR21 U3052 ( .A(\u_cordic/mycordic/sub_236/carry [3]), .B(
        \u_cordic/mycordic/present_ANGLE_table[5][3] ), .Q(n467) );
  INV3 U3053 ( .A(n468), .Q(\u_cordic/mycordic/sub_236/carry [5]) );
  NOR21 U3054 ( .A(\u_cordic/mycordic/sub_236/carry [4]), .B(
        \u_cordic/mycordic/present_ANGLE_table[5][4] ), .Q(n468) );
  INV3 U3055 ( .A(n469), .Q(\u_cordic/mycordic/sub_236/carry [6]) );
  NOR21 U3056 ( .A(\u_cordic/mycordic/sub_236/carry [5]), .B(
        \u_cordic/mycordic/present_ANGLE_table[5][5] ), .Q(n469) );
  INV3 U3057 ( .A(n470), .Q(\u_cordic/mycordic/sub_236/carry [7]) );
  NOR21 U3058 ( .A(\u_cordic/mycordic/sub_236/carry [6]), .B(
        \u_cordic/mycordic/present_ANGLE_table[5][6] ), .Q(n470) );
  INV3 U3059 ( .A(n471), .Q(\u_cordic/mycordic/sub_236/carry [8]) );
  NOR21 U3060 ( .A(\u_cordic/mycordic/sub_236/carry [7]), .B(
        \u_cordic/mycordic/present_ANGLE_table[5][7] ), .Q(n471) );
  INV3 U3061 ( .A(n472), .Q(\u_cordic/mycordic/sub_236/carry [9]) );
  NOR21 U3062 ( .A(\u_cordic/mycordic/sub_236/carry [8]), .B(
        \u_cordic/mycordic/present_ANGLE_table[5][8] ), .Q(n472) );
  INV3 U3063 ( .A(n473), .Q(\u_cordic/mycordic/sub_236/carry [10]) );
  NOR21 U3064 ( .A(\u_cordic/mycordic/sub_236/carry [9]), .B(
        \u_cordic/mycordic/present_ANGLE_table[5][9] ), .Q(n473) );
  INV3 U3065 ( .A(n461), .Q(\u_cordic/mycordic/sub_236/carry [11]) );
  NOR21 U3066 ( .A(\u_cordic/mycordic/sub_236/carry [10]), .B(
        \u_cordic/mycordic/present_ANGLE_table[5][10] ), .Q(n461) );
  INV3 U3067 ( .A(n462), .Q(\u_cordic/mycordic/sub_236/carry [12]) );
  NOR21 U3068 ( .A(\u_cordic/mycordic/sub_236/carry [11]), .B(
        \u_cordic/mycordic/present_ANGLE_table[5][11] ), .Q(n462) );
  INV3 U3069 ( .A(n463), .Q(\u_cordic/mycordic/sub_236/carry [13]) );
  NOR21 U3070 ( .A(\u_cordic/mycordic/sub_236/carry [12]), .B(
        \u_cordic/mycordic/present_ANGLE_table[5][12] ), .Q(n463) );
  INV3 U3071 ( .A(n464), .Q(\u_cordic/mycordic/sub_236/carry [14]) );
  NOR21 U3072 ( .A(\u_cordic/mycordic/sub_236/carry [13]), .B(
        \u_cordic/mycordic/present_ANGLE_table[5][13] ), .Q(n464) );
  NAND22 U3073 ( .A(\u_coder/n232 ), .B(\u_coder/n233 ), .Q(\u_coder/n344 ) );
  NAND22 U3074 ( .A(sig_coder_outSinQMasked[0]), .B(n1813), .Q(\u_coder/n232 )
         );
  INV3 U3075 ( .A(\u_coder/n218 ), .Q(n2172) );
  INV3 U3076 ( .A(n404), .Q(\u_cordic/mycordic/add_191/carry[5] ) );
  NOR21 U3077 ( .A(\u_cordic/mycordic/add_191/carry[4] ), .B(
        \u_cordic/mycordic/present_ANGLE_table[1][4] ), .Q(n404) );
  INV3 U3078 ( .A(n419), .Q(\u_cordic/mycordic/add_202/carry [4]) );
  NOR21 U3079 ( .A(\u_cordic/mycordic/add_202/carry [3]), .B(
        \u_cordic/mycordic/present_ANGLE_table[2][3] ), .Q(n419) );
  INV3 U3080 ( .A(n434), .Q(\u_cordic/mycordic/add_213/carry[3] ) );
  NOR21 U3081 ( .A(\u_cordic/mycordic/add_213/carry[2] ), .B(
        \u_cordic/mycordic/present_ANGLE_table[3][2] ), .Q(n434) );
  NOR21 U3082 ( .A(\u_cordic/mycordic/present_I_table[4][3] ), .B(n2651), .Q(
        n3030) );
  INV3 U3083 ( .A(n3031), .Q(n2651) );
  NAND22 U3084 ( .A(\u_coder/n248 ), .B(\u_coder/n249 ), .Q(\u_coder/n348 ) );
  NAND22 U3085 ( .A(sig_coder_outSinIMasked[2]), .B(\u_coder/n245 ), .Q(
        \u_coder/n249 ) );
  NAND22 U3086 ( .A(\u_coder/n248 ), .B(\u_coder/n250 ), .Q(\u_coder/n349 ) );
  NAND22 U3087 ( .A(sig_coder_outSinIMasked[1]), .B(\u_coder/n245 ), .Q(
        \u_coder/n250 ) );
  NAND22 U3088 ( .A(\u_coder/n252 ), .B(\u_coder/n253 ), .Q(\u_coder/n350 ) );
  NAND22 U3089 ( .A(sig_coder_outSinIMasked[0]), .B(\u_coder/n245 ), .Q(
        \u_coder/n252 ) );
  NAND22 U3090 ( .A(\u_cordic/mycordic/present_I_table[5][4] ), .B(n180), .Q(
        n3015) );
  NOR21 U3091 ( .A(n181), .B(n494), .Q(\u_cordic/mycordic/r173/carry [10]) );
  INV3 U3092 ( .A(\u_cordic/mycordic/r173/carry [9]), .Q(n494) );
  NOR21 U3093 ( .A(n228), .B(n495), .Q(\u_cordic/mycordic/r173/carry [11]) );
  INV3 U3094 ( .A(\u_cordic/mycordic/r173/carry [10]), .Q(n495) );
  NOR21 U3095 ( .A(n228), .B(n557), .Q(\u_cordic/mycordic/add_262/carry [11])
         );
  INV3 U3096 ( .A(\u_cordic/mycordic/add_262/carry [10]), .Q(n557) );
  NOR21 U3097 ( .A(n229), .B(n496), .Q(\u_cordic/mycordic/r173/carry [12]) );
  INV3 U3098 ( .A(\u_cordic/mycordic/r173/carry [11]), .Q(n496) );
  NOR21 U3099 ( .A(n229), .B(n558), .Q(\u_cordic/mycordic/add_262/carry [12])
         );
  INV3 U3100 ( .A(\u_cordic/mycordic/add_262/carry [11]), .Q(n558) );
  NOR21 U3101 ( .A(n266), .B(n497), .Q(\u_cordic/mycordic/r173/carry [13]) );
  INV3 U3102 ( .A(\u_cordic/mycordic/r173/carry [12]), .Q(n497) );
  NOR21 U3103 ( .A(n266), .B(n559), .Q(\u_cordic/mycordic/add_262/carry [13])
         );
  INV3 U3104 ( .A(\u_cordic/mycordic/add_262/carry [12]), .Q(n559) );
  NOR21 U3105 ( .A(n267), .B(n498), .Q(\u_cordic/mycordic/r173/carry [14]) );
  INV3 U3106 ( .A(\u_cordic/mycordic/r173/carry [13]), .Q(n498) );
  NOR21 U3107 ( .A(n267), .B(n560), .Q(\u_cordic/mycordic/add_262/carry [14])
         );
  INV3 U3108 ( .A(\u_cordic/mycordic/add_262/carry [13]), .Q(n560) );
  NOR21 U3109 ( .A(\u_cordic/mycordic/present_I_table[4][1] ), .B(n2653), .Q(
        n3026) );
  INV3 U3110 ( .A(n3027), .Q(n2653) );
  INV3 U3111 ( .A(n410), .Q(\u_cordic/mycordic/sub_196/carry[15] ) );
  NOR21 U3112 ( .A(\u_cordic/mycordic/sub_196/carry[14] ), .B(
        \u_cordic/mycordic/present_ANGLE_table[1][14] ), .Q(n410) );
  INV3 U3113 ( .A(n425), .Q(\u_cordic/mycordic/sub_207/carry [15]) );
  NOR21 U3114 ( .A(\u_cordic/mycordic/sub_207/carry [14]), .B(
        \u_cordic/mycordic/present_ANGLE_table[2][14] ), .Q(n425) );
  INV3 U3115 ( .A(n439), .Q(\u_cordic/mycordic/sub_218/carry[15] ) );
  NOR21 U3116 ( .A(\u_cordic/mycordic/sub_218/carry[14] ), .B(
        \u_cordic/mycordic/present_ANGLE_table[3][14] ), .Q(n439) );
  INV3 U3117 ( .A(n452), .Q(\u_cordic/mycordic/sub_229/carry[15] ) );
  NOR21 U3118 ( .A(\u_cordic/mycordic/sub_229/carry[14] ), .B(
        \u_cordic/mycordic/present_ANGLE_table[4][14] ), .Q(n452) );
  INV3 U3119 ( .A(n465), .Q(\u_cordic/mycordic/sub_236/carry [15]) );
  NOR21 U3120 ( .A(\u_cordic/mycordic/sub_236/carry [14]), .B(
        \u_cordic/mycordic/present_ANGLE_table[5][14] ), .Q(n465) );
  NOR21 U3121 ( .A(n141), .B(n399), .Q(\u_cordic/mycordic/r173/carry [7]) );
  NOR21 U3122 ( .A(n182), .B(n400), .Q(\u_cordic/mycordic/r173/carry [9]) );
  NOR21 U3123 ( .A(n181), .B(n476), .Q(\u_cordic/mycordic/add_262/carry [10])
         );
  NOR21 U3124 ( .A(n268), .B(n499), .Q(\u_cordic/mycordic/r173/carry [15]) );
  XNR21 U3125 ( .A(\u_cordic/mycordic/r173/carry [13]), .B(
        \u_cordic/mycordic/present_ANGLE_table[6][13] ), .Q(n375) );
  INV3 U3126 ( .A(\u_cordic/mycordic/n399 ), .Q(n1868) );
  NAND22 U3127 ( .A(\u_cordic/mycordic/next_ANGLE_table[6][15] ), .B(n1215), 
        .Q(\u_cordic/mycordic/n399 ) );
  INV3 U3128 ( .A(\u_coder/n272 ), .Q(n1925) );
  AOI221 U3129 ( .A(\u_coder/n263 ), .B(\u_coder/j [9]), .C(n2169), .D(
        \u_coder/N1022 ), .Q(\u_coder/n272 ) );
  INV3 U3130 ( .A(\u_coder/n294 ), .Q(n1945) );
  AOI221 U3131 ( .A(n894), .B(\u_coder/i [9]), .C(n2156), .D(\u_coder/N716 ), 
        .Q(\u_coder/n294 ) );
  INV3 U3132 ( .A(\u_coder/n275 ), .Q(n1922) );
  AOI221 U3133 ( .A(n890), .B(\u_coder/j [6]), .C(n2169), .D(\u_coder/N1019 ), 
        .Q(\u_coder/n275 ) );
  INV3 U3134 ( .A(\u_coder/n271 ), .Q(n1926) );
  AOI221 U3135 ( .A(n890), .B(\u_coder/j [10]), .C(n2169), .D(\u_coder/N1023 ), 
        .Q(\u_coder/n271 ) );
  INV3 U3136 ( .A(\u_coder/n297 ), .Q(n1942) );
  AOI221 U3137 ( .A(n893), .B(\u_coder/i [6]), .C(n2156), .D(\u_coder/N713 ), 
        .Q(\u_coder/n297 ) );
  INV3 U3138 ( .A(\u_coder/n293 ), .Q(n1946) );
  AOI221 U3139 ( .A(n894), .B(\u_coder/i [10]), .C(n2156), .D(\u_coder/N717 ), 
        .Q(\u_coder/n293 ) );
  INV3 U3140 ( .A(\u_coder/n274 ), .Q(n1923) );
  AOI221 U3141 ( .A(n890), .B(\u_coder/j [7]), .C(n2169), .D(\u_coder/N1020 ), 
        .Q(\u_coder/n274 ) );
  INV3 U3142 ( .A(\u_coder/n273 ), .Q(n1924) );
  AOI221 U3143 ( .A(n890), .B(\u_coder/j [8]), .C(n2169), .D(\u_coder/N1021 ), 
        .Q(\u_coder/n273 ) );
  INV3 U3144 ( .A(\u_coder/n296 ), .Q(n1943) );
  AOI221 U3145 ( .A(n893), .B(\u_coder/i [7]), .C(n2156), .D(\u_coder/N714 ), 
        .Q(\u_coder/n296 ) );
  INV3 U3146 ( .A(\u_coder/n295 ), .Q(n1944) );
  AOI221 U3147 ( .A(n894), .B(\u_coder/i [8]), .C(n2156), .D(\u_coder/N715 ), 
        .Q(\u_coder/n295 ) );
  INV3 U3148 ( .A(\u_coder/n299 ), .Q(n1940) );
  AOI221 U3149 ( .A(n892), .B(\u_coder/i [4]), .C(n2156), .D(\u_coder/N711 ), 
        .Q(\u_coder/n299 ) );
  INV3 U3150 ( .A(\u_coder/n298 ), .Q(n1941) );
  AOI221 U3151 ( .A(n893), .B(\u_coder/i [5]), .C(n2156), .D(\u_coder/N712 ), 
        .Q(\u_coder/n298 ) );
  INV3 U3152 ( .A(\u_coder/n279 ), .Q(n1918) );
  AOI221 U3153 ( .A(\u_coder/N1015 ), .B(n2169), .C(\u_coder/n263 ), .D(
        \u_coder/j [2]), .Q(\u_coder/n279 ) );
  INV3 U3154 ( .A(\u_coder/n178 ), .Q(n1810) );
  AOI211 U3155 ( .A(\u_coder/n179 ), .B(sig_coder_outSinQ[3]), .C(
        \u_coder/n180 ), .Q(\u_coder/n178 ) );
  INV3 U3156 ( .A(\u_cordic/mycordic/n506 ), .Q(n1466) );
  AOI221 U3157 ( .A(\u_cordic/mycordic/N345 ), .B(\u_cordic/mycordic/n336 ), 
        .C(\u_cordic/mycordic/N377 ), .D(n1904), .Q(\u_cordic/mycordic/n506 )
         );
  XNR21 U3158 ( .A(\u_cordic/mycordic/present_ANGLE_table[1][13] ), .B(
        \u_cordic/mycordic/sub_196/carry[13] ), .Q(\u_cordic/mycordic/N377 )
         );
  XOR21 U3159 ( .A(\u_cordic/mycordic/present_ANGLE_table[1][13] ), .B(
        \u_cordic/mycordic/add_191/carry[13] ), .Q(\u_cordic/mycordic/N345 )
         );
  INV3 U3160 ( .A(\u_cordic/mycordic/n505 ), .Q(n1467) );
  AOI221 U3161 ( .A(\u_cordic/mycordic/N346 ), .B(n772), .C(
        \u_cordic/mycordic/N378 ), .D(n1904), .Q(\u_cordic/mycordic/n505 ) );
  XNR21 U3162 ( .A(\u_cordic/mycordic/present_ANGLE_table[1][14] ), .B(
        \u_cordic/mycordic/sub_196/carry[14] ), .Q(\u_cordic/mycordic/N378 )
         );
  XOR21 U3163 ( .A(\u_cordic/mycordic/present_ANGLE_table[1][14] ), .B(
        \u_cordic/mycordic/add_191/carry[14] ), .Q(\u_cordic/mycordic/N346 )
         );
  INV3 U3164 ( .A(\u_cordic/mycordic/n490 ), .Q(n1559) );
  AOI221 U3165 ( .A(\u_cordic/mycordic/N409 ), .B(n778), .C(
        \u_cordic/mycordic/N441 ), .D(n1908), .Q(\u_cordic/mycordic/n490 ) );
  XNR21 U3166 ( .A(\u_cordic/mycordic/present_ANGLE_table[2][13] ), .B(
        \u_cordic/mycordic/sub_207/carry [13]), .Q(\u_cordic/mycordic/N441 )
         );
  XOR21 U3167 ( .A(\u_cordic/mycordic/present_ANGLE_table[2][13] ), .B(
        \u_cordic/mycordic/add_202/carry [13]), .Q(\u_cordic/mycordic/N409 )
         );
  INV3 U3168 ( .A(\u_cordic/mycordic/n489 ), .Q(n1560) );
  AOI221 U3169 ( .A(\u_cordic/mycordic/N410 ), .B(\u_cordic/mycordic/n332 ), 
        .C(\u_cordic/mycordic/N442 ), .D(n1908), .Q(\u_cordic/mycordic/n489 )
         );
  XNR21 U3170 ( .A(\u_cordic/mycordic/present_ANGLE_table[2][14] ), .B(
        \u_cordic/mycordic/sub_207/carry [14]), .Q(\u_cordic/mycordic/N442 )
         );
  XOR21 U3171 ( .A(\u_cordic/mycordic/present_ANGLE_table[2][14] ), .B(
        \u_cordic/mycordic/add_202/carry [14]), .Q(\u_cordic/mycordic/N410 )
         );
  INV3 U3172 ( .A(\u_cordic/mycordic/n474 ), .Q(n1534) );
  AOI221 U3173 ( .A(\u_cordic/mycordic/N469 ), .B(\u_cordic/mycordic/n363 ), 
        .C(\u_cordic/mycordic/N497 ), .D(n1907), .Q(\u_cordic/mycordic/n474 )
         );
  XNR21 U3174 ( .A(\u_cordic/mycordic/present_ANGLE_table[3][13] ), .B(
        \u_cordic/mycordic/sub_218/carry[13] ), .Q(\u_cordic/mycordic/N497 )
         );
  XOR21 U3175 ( .A(\u_cordic/mycordic/present_ANGLE_table[3][13] ), .B(
        \u_cordic/mycordic/add_213/carry[13] ), .Q(\u_cordic/mycordic/N469 )
         );
  INV3 U3176 ( .A(\u_cordic/mycordic/n459 ), .Q(n1509) );
  AOI221 U3177 ( .A(\u_cordic/mycordic/N513 ), .B(\u_cordic/mycordic/n456 ), 
        .C(\u_cordic/mycordic/N530 ), .D(n1906), .Q(\u_cordic/mycordic/n459 )
         );
  XNR21 U3178 ( .A(\u_cordic/mycordic/present_ANGLE_table[4][12] ), .B(
        \u_cordic/mycordic/sub_229/carry[12] ), .Q(\u_cordic/mycordic/N530 )
         );
  XOR21 U3179 ( .A(\u_cordic/mycordic/present_ANGLE_table[4][12] ), .B(
        \u_cordic/mycordic/add_224/carry[12] ), .Q(\u_cordic/mycordic/N513 )
         );
  INV3 U3180 ( .A(\u_cordic/mycordic/n458 ), .Q(n1510) );
  AOI221 U3181 ( .A(\u_cordic/mycordic/N514 ), .B(n776), .C(
        \u_cordic/mycordic/N531 ), .D(n1906), .Q(\u_cordic/mycordic/n458 ) );
  XNR21 U3182 ( .A(\u_cordic/mycordic/present_ANGLE_table[4][13] ), .B(
        \u_cordic/mycordic/sub_229/carry[13] ), .Q(\u_cordic/mycordic/N531 )
         );
  XOR21 U3183 ( .A(\u_cordic/mycordic/present_ANGLE_table[4][13] ), .B(
        \u_cordic/mycordic/add_224/carry[13] ), .Q(\u_cordic/mycordic/N514 )
         );
  INV3 U3184 ( .A(\u_cordic/mycordic/n457 ), .Q(n1511) );
  AOI221 U3185 ( .A(\u_cordic/mycordic/N515 ), .B(n776), .C(
        \u_cordic/mycordic/N532 ), .D(n1906), .Q(\u_cordic/mycordic/n457 ) );
  XNR21 U3186 ( .A(\u_cordic/mycordic/present_ANGLE_table[4][14] ), .B(
        \u_cordic/mycordic/sub_229/carry[14] ), .Q(\u_cordic/mycordic/N532 )
         );
  XOR21 U3187 ( .A(\u_cordic/mycordic/present_ANGLE_table[4][14] ), .B(
        \u_cordic/mycordic/add_224/carry[14] ), .Q(\u_cordic/mycordic/N515 )
         );
  INV3 U3188 ( .A(\u_decoder/fir_filter/n1078 ), .Q(n2268) );
  AOI221 U3189 ( .A(\u_decoder/fir_filter/I_data_mult_4 [8]), .B(n1091), .C(
        \u_decoder/fir_filter/I_data_mult_4_buff [8]), .D(n1163), .Q(
        \u_decoder/fir_filter/n1078 ) );
  AOI211 U3190 ( .A(n365), .B(n347), .C(n2951), .Q(
        \u_decoder/fir_filter/I_data_mult_4 [8]) );
  INV3 U3191 ( .A(\u_decoder/fir_filter/n781 ), .Q(n2339) );
  AOI221 U3192 ( .A(\u_decoder/fir_filter/Q_data_mult_4 [8]), .B(n1083), .C(
        \u_decoder/fir_filter/Q_data_mult_4_buff [8]), .D(n1166), .Q(
        \u_decoder/fir_filter/n781 ) );
  AOI211 U3193 ( .A(n366), .B(n348), .C(n2865), .Q(
        \u_decoder/fir_filter/Q_data_mult_4 [8]) );
  INV3 U3194 ( .A(\u_cordic/mycordic/n504 ), .Q(n1468) );
  AOI221 U3195 ( .A(\u_cordic/mycordic/N347 ), .B(\u_cordic/mycordic/n336 ), 
        .C(\u_cordic/mycordic/N379 ), .D(n1904), .Q(\u_cordic/mycordic/n504 )
         );
  XNR21 U3196 ( .A(\u_cordic/mycordic/sub_196/carry[15] ), .B(
        \u_cordic/mycordic/present_ANGLE_table[1][15] ), .Q(
        \u_cordic/mycordic/N379 ) );
  XOR21 U3197 ( .A(\u_cordic/mycordic/add_191/carry[15] ), .B(
        \u_cordic/mycordic/present_ANGLE_table[1][15] ), .Q(
        \u_cordic/mycordic/N347 ) );
  INV3 U3198 ( .A(\u_cordic/mycordic/n488 ), .Q(n1561) );
  AOI221 U3199 ( .A(\u_cordic/mycordic/N411 ), .B(n778), .C(
        \u_cordic/mycordic/N443 ), .D(n1908), .Q(\u_cordic/mycordic/n488 ) );
  XNR21 U3200 ( .A(\u_cordic/mycordic/sub_207/carry [15]), .B(
        \u_cordic/mycordic/present_ANGLE_table[2][15] ), .Q(
        \u_cordic/mycordic/N443 ) );
  XOR21 U3201 ( .A(\u_cordic/mycordic/add_202/carry [15]), .B(
        \u_cordic/mycordic/present_ANGLE_table[2][15] ), .Q(
        \u_cordic/mycordic/N411 ) );
  INV3 U3202 ( .A(\u_cordic/mycordic/n472 ), .Q(n1536) );
  AOI221 U3203 ( .A(\u_cordic/mycordic/N471 ), .B(\u_cordic/mycordic/n363 ), 
        .C(\u_cordic/mycordic/N499 ), .D(n1907), .Q(\u_cordic/mycordic/n472 )
         );
  XNR21 U3204 ( .A(\u_cordic/mycordic/sub_218/carry[15] ), .B(
        \u_cordic/mycordic/present_ANGLE_table[3][15] ), .Q(
        \u_cordic/mycordic/N499 ) );
  XOR21 U3205 ( .A(\u_cordic/mycordic/add_213/carry[15] ), .B(
        \u_cordic/mycordic/present_ANGLE_table[3][15] ), .Q(
        \u_cordic/mycordic/N471 ) );
  INV3 U3206 ( .A(\u_cordic/mycordic/n455 ), .Q(n1512) );
  AOI221 U3207 ( .A(\u_cordic/mycordic/N516 ), .B(\u_cordic/mycordic/n456 ), 
        .C(\u_cordic/mycordic/N533 ), .D(n1906), .Q(\u_cordic/mycordic/n455 )
         );
  XNR21 U3208 ( .A(\u_cordic/mycordic/sub_229/carry[15] ), .B(
        \u_cordic/mycordic/present_ANGLE_table[4][15] ), .Q(
        \u_cordic/mycordic/N533 ) );
  XOR21 U3209 ( .A(\u_cordic/mycordic/add_224/carry[15] ), .B(
        \u_cordic/mycordic/present_ANGLE_table[4][15] ), .Q(
        \u_cordic/mycordic/N516 ) );
  INV3 U3210 ( .A(\u_decoder/fir_filter/n989 ), .Q(n2629) );
  AOI221 U3211 ( .A(\u_decoder/fir_filter/I_data_add_7 [7]), .B(n1092), .C(
        \u_decoder/fir_filter/I_data_add_7_buff [7]), .D(n1164), .Q(
        \u_decoder/fir_filter/n989 ) );
  INV3 U3212 ( .A(\u_decoder/fir_filter/n988 ), .Q(n2628) );
  AOI221 U3213 ( .A(\u_decoder/fir_filter/I_data_add_7 [8]), .B(n1092), .C(
        \u_decoder/fir_filter/I_data_add_7_buff [8]), .D(n1164), .Q(
        \u_decoder/fir_filter/n988 ) );
  INV3 U3214 ( .A(\u_decoder/fir_filter/n987 ), .Q(n2627) );
  AOI221 U3215 ( .A(\u_decoder/fir_filter/I_data_add_7 [9]), .B(n1092), .C(
        \u_decoder/fir_filter/I_data_add_7_buff [9]), .D(n1164), .Q(
        \u_decoder/fir_filter/n987 ) );
  INV3 U3216 ( .A(\u_decoder/fir_filter/n968 ), .Q(n2614) );
  AOI221 U3217 ( .A(\u_decoder/fir_filter/I_data_add_6 [7]), .B(n1092), .C(
        \u_decoder/fir_filter/I_data_add_6_buff [7]), .D(n1165), .Q(
        \u_decoder/fir_filter/n968 ) );
  INV3 U3218 ( .A(\u_decoder/fir_filter/n967 ), .Q(n2613) );
  AOI221 U3219 ( .A(\u_decoder/fir_filter/I_data_add_6 [8]), .B(n1092), .C(
        \u_decoder/fir_filter/I_data_add_6_buff [8]), .D(n1165), .Q(
        \u_decoder/fir_filter/n967 ) );
  INV3 U3220 ( .A(\u_decoder/fir_filter/n966 ), .Q(n2612) );
  AOI221 U3221 ( .A(\u_decoder/fir_filter/I_data_add_6 [9]), .B(n1093), .C(
        \u_decoder/fir_filter/I_data_add_6_buff [9]), .D(n1165), .Q(
        \u_decoder/fir_filter/n966 ) );
  INV3 U3222 ( .A(\u_decoder/fir_filter/n947 ), .Q(n2599) );
  AOI221 U3223 ( .A(\u_decoder/fir_filter/I_data_add_5 [7]), .B(n1093), .C(
        \u_decoder/fir_filter/I_data_add_5_buff [7]), .D(n1166), .Q(
        \u_decoder/fir_filter/n947 ) );
  INV3 U3224 ( .A(\u_decoder/fir_filter/n946 ), .Q(n2598) );
  AOI221 U3225 ( .A(\u_decoder/fir_filter/I_data_add_5 [8]), .B(n1093), .C(
        \u_decoder/fir_filter/I_data_add_5_buff [8]), .D(n1166), .Q(
        \u_decoder/fir_filter/n946 ) );
  INV3 U3226 ( .A(\u_decoder/fir_filter/n945 ), .Q(n2597) );
  AOI221 U3227 ( .A(\u_decoder/fir_filter/I_data_add_5 [9]), .B(n1093), .C(
        \u_decoder/fir_filter/I_data_add_5_buff [9]), .D(n1166), .Q(
        \u_decoder/fir_filter/n945 ) );
  INV3 U3228 ( .A(\u_decoder/fir_filter/n925 ), .Q(n2583) );
  AOI221 U3229 ( .A(\u_decoder/fir_filter/I_data_add_4 [8]), .B(n1094), .C(
        \u_decoder/fir_filter/I_data_add_4_buff [8]), .D(n1158), .Q(
        \u_decoder/fir_filter/n925 ) );
  INV3 U3230 ( .A(\u_decoder/fir_filter/n905 ), .Q(n2569) );
  AOI221 U3231 ( .A(\u_decoder/fir_filter/I_data_add_3 [7]), .B(n1095), .C(
        \u_decoder/fir_filter/I_data_add_3_buff [7]), .D(n1157), .Q(
        \u_decoder/fir_filter/n905 ) );
  INV3 U3232 ( .A(\u_decoder/fir_filter/n904 ), .Q(n2568) );
  AOI221 U3233 ( .A(\u_decoder/fir_filter/I_data_add_3 [8]), .B(n1095), .C(
        \u_decoder/fir_filter/I_data_add_3_buff [8]), .D(n1158), .Q(
        \u_decoder/fir_filter/n904 ) );
  INV3 U3234 ( .A(\u_decoder/fir_filter/n903 ), .Q(n2567) );
  AOI221 U3235 ( .A(\u_decoder/fir_filter/I_data_add_3 [9]), .B(n1095), .C(
        \u_decoder/fir_filter/I_data_add_3_buff [9]), .D(n1151), .Q(
        \u_decoder/fir_filter/n903 ) );
  INV3 U3236 ( .A(\u_decoder/fir_filter/n884 ), .Q(n2554) );
  AOI221 U3237 ( .A(\u_decoder/fir_filter/I_data_add_2 [7]), .B(n1096), .C(
        \u_decoder/fir_filter/I_data_add_2_buff [7]), .D(n1166), .Q(
        \u_decoder/fir_filter/n884 ) );
  INV3 U3238 ( .A(\u_decoder/fir_filter/n883 ), .Q(n2553) );
  AOI221 U3239 ( .A(\u_decoder/fir_filter/I_data_add_2 [8]), .B(n1096), .C(
        \u_decoder/fir_filter/I_data_add_2_buff [8]), .D(n1166), .Q(
        \u_decoder/fir_filter/n883 ) );
  INV3 U3240 ( .A(\u_decoder/fir_filter/n882 ), .Q(n2552) );
  AOI221 U3241 ( .A(\u_decoder/fir_filter/I_data_add_2 [9]), .B(n1096), .C(
        \u_decoder/fir_filter/I_data_add_2_buff [9]), .D(n1163), .Q(
        \u_decoder/fir_filter/n882 ) );
  INV3 U3242 ( .A(\u_decoder/fir_filter/n863 ), .Q(n2534) );
  AOI221 U3243 ( .A(\u_decoder/fir_filter/I_data_add_1 [7]), .B(n1097), .C(
        \u_decoder/fir_filter/I_data_add_1_buff [7]), .D(n1160), .Q(
        \u_decoder/fir_filter/n863 ) );
  INV3 U3244 ( .A(\u_decoder/fir_filter/n862 ), .Q(n2531) );
  AOI221 U3245 ( .A(\u_decoder/fir_filter/I_data_add_1 [8]), .B(n1097), .C(
        \u_decoder/fir_filter/I_data_add_1_buff [8]), .D(n1162), .Q(
        \u_decoder/fir_filter/n862 ) );
  INV3 U3246 ( .A(\u_decoder/fir_filter/n861 ), .Q(n2530) );
  AOI221 U3247 ( .A(\u_decoder/fir_filter/I_data_add_1 [9]), .B(n1097), .C(
        \u_decoder/fir_filter/I_data_add_1_buff [9]), .D(n1161), .Q(
        \u_decoder/fir_filter/n861 ) );
  INV3 U3248 ( .A(\u_decoder/fir_filter/n691 ), .Q(n2509) );
  AOI221 U3249 ( .A(\u_decoder/fir_filter/Q_data_add_7 [7]), .B(n1084), .C(
        \u_decoder/fir_filter/Q_data_add_7_buff [7]), .D(n1163), .Q(
        \u_decoder/fir_filter/n691 ) );
  INV3 U3250 ( .A(\u_decoder/fir_filter/n690 ), .Q(n2508) );
  AOI221 U3251 ( .A(\u_decoder/fir_filter/Q_data_add_7 [8]), .B(n1084), .C(
        \u_decoder/fir_filter/Q_data_add_7_buff [8]), .D(n1163), .Q(
        \u_decoder/fir_filter/n690 ) );
  INV3 U3252 ( .A(\u_decoder/fir_filter/n689 ), .Q(n2507) );
  AOI221 U3253 ( .A(\u_decoder/fir_filter/Q_data_add_7 [9]), .B(n1085), .C(
        \u_decoder/fir_filter/Q_data_add_7_buff [9]), .D(n1163), .Q(
        \u_decoder/fir_filter/n689 ) );
  INV3 U3254 ( .A(\u_decoder/fir_filter/n670 ), .Q(n2494) );
  AOI221 U3255 ( .A(\u_decoder/fir_filter/Q_data_add_6 [7]), .B(n1085), .C(
        \u_decoder/fir_filter/Q_data_add_6_buff [7]), .D(n1165), .Q(
        \u_decoder/fir_filter/n670 ) );
  INV3 U3256 ( .A(\u_decoder/fir_filter/n669 ), .Q(n2493) );
  AOI221 U3257 ( .A(\u_decoder/fir_filter/Q_data_add_6 [8]), .B(n1085), .C(
        \u_decoder/fir_filter/Q_data_add_6_buff [8]), .D(n1166), .Q(
        \u_decoder/fir_filter/n669 ) );
  INV3 U3258 ( .A(\u_decoder/fir_filter/n668 ), .Q(n2492) );
  AOI221 U3259 ( .A(\u_decoder/fir_filter/Q_data_add_6 [9]), .B(n1085), .C(
        \u_decoder/fir_filter/Q_data_add_6_buff [9]), .D(n1163), .Q(
        \u_decoder/fir_filter/n668 ) );
  INV3 U3260 ( .A(\u_decoder/fir_filter/n649 ), .Q(n2479) );
  AOI221 U3261 ( .A(\u_decoder/fir_filter/Q_data_add_5 [7]), .B(n1086), .C(
        \u_decoder/fir_filter/Q_data_add_5_buff [7]), .D(n1166), .Q(
        \u_decoder/fir_filter/n649 ) );
  INV3 U3262 ( .A(\u_decoder/fir_filter/n648 ), .Q(n2478) );
  AOI221 U3263 ( .A(\u_decoder/fir_filter/Q_data_add_5 [8]), .B(n1086), .C(
        \u_decoder/fir_filter/Q_data_add_5_buff [8]), .D(n1163), .Q(
        \u_decoder/fir_filter/n648 ) );
  INV3 U3264 ( .A(\u_decoder/fir_filter/n647 ), .Q(n2477) );
  AOI221 U3265 ( .A(\u_decoder/fir_filter/Q_data_add_5 [9]), .B(n1086), .C(
        \u_decoder/fir_filter/Q_data_add_5_buff [9]), .D(n1163), .Q(
        \u_decoder/fir_filter/n647 ) );
  INV3 U3266 ( .A(\u_decoder/fir_filter/n627 ), .Q(n2463) );
  AOI221 U3267 ( .A(\u_decoder/fir_filter/Q_data_add_4 [8]), .B(n1087), .C(
        \u_decoder/fir_filter/Q_data_add_4_buff [8]), .D(n1162), .Q(
        \u_decoder/fir_filter/n627 ) );
  INV3 U3268 ( .A(\u_decoder/fir_filter/n607 ), .Q(n2449) );
  AOI221 U3269 ( .A(\u_decoder/fir_filter/Q_data_add_3 [7]), .B(n1088), .C(
        \u_decoder/fir_filter/Q_data_add_3_buff [7]), .D(n1162), .Q(
        \u_decoder/fir_filter/n607 ) );
  INV3 U3270 ( .A(\u_decoder/fir_filter/n606 ), .Q(n2448) );
  AOI221 U3271 ( .A(\u_decoder/fir_filter/Q_data_add_3 [8]), .B(n1088), .C(
        \u_decoder/fir_filter/Q_data_add_3_buff [8]), .D(n1161), .Q(
        \u_decoder/fir_filter/n606 ) );
  INV3 U3272 ( .A(\u_decoder/fir_filter/n605 ), .Q(n2447) );
  AOI221 U3273 ( .A(\u_decoder/fir_filter/Q_data_add_3 [9]), .B(n1088), .C(
        \u_decoder/fir_filter/Q_data_add_3_buff [9]), .D(n1161), .Q(
        \u_decoder/fir_filter/n605 ) );
  INV3 U3274 ( .A(\u_decoder/fir_filter/n586 ), .Q(n2434) );
  AOI221 U3275 ( .A(\u_decoder/fir_filter/Q_data_add_2 [7]), .B(n1089), .C(
        \u_decoder/fir_filter/Q_data_add_2_buff [7]), .D(n1161), .Q(
        \u_decoder/fir_filter/n586 ) );
  INV3 U3276 ( .A(\u_decoder/fir_filter/n585 ), .Q(n2433) );
  AOI221 U3277 ( .A(\u_decoder/fir_filter/Q_data_add_2 [8]), .B(n1089), .C(
        \u_decoder/fir_filter/Q_data_add_2_buff [8]), .D(n1161), .Q(
        \u_decoder/fir_filter/n585 ) );
  INV3 U3278 ( .A(\u_decoder/fir_filter/n584 ), .Q(n2432) );
  AOI221 U3279 ( .A(\u_decoder/fir_filter/Q_data_add_2 [9]), .B(n1089), .C(
        \u_decoder/fir_filter/Q_data_add_2_buff [9]), .D(n1161), .Q(
        \u_decoder/fir_filter/n584 ) );
  INV3 U3280 ( .A(\u_decoder/fir_filter/n565 ), .Q(n2414) );
  AOI221 U3281 ( .A(\u_decoder/fir_filter/Q_data_add_1 [7]), .B(n1090), .C(
        \u_decoder/fir_filter/Q_data_add_1_buff [7]), .D(n1162), .Q(
        \u_decoder/fir_filter/n565 ) );
  INV3 U3282 ( .A(\u_decoder/fir_filter/n564 ), .Q(n2411) );
  AOI221 U3283 ( .A(\u_decoder/fir_filter/Q_data_add_1 [8]), .B(n1090), .C(
        \u_decoder/fir_filter/Q_data_add_1_buff [8]), .D(n1161), .Q(
        \u_decoder/fir_filter/n564 ) );
  INV3 U3284 ( .A(\u_decoder/fir_filter/n563 ), .Q(n2410) );
  AOI221 U3285 ( .A(\u_decoder/fir_filter/Q_data_add_1 [9]), .B(n1090), .C(
        \u_decoder/fir_filter/Q_data_add_1_buff [9]), .D(n1161), .Q(
        \u_decoder/fir_filter/n563 ) );
  NAND41 U3286 ( .A(\u_coder/n331 ), .B(\u_coder/n332 ), .C(\u_coder/n333 ), 
        .D(\u_coder/n334 ), .Q(\u_coder/n256 ) );
  NOR40 U3287 ( .A(\u_coder/i [9]), .B(\u_coder/i [8]), .C(\u_coder/i [7]), 
        .D(\u_coder/i [6]), .Q(\u_coder/n334 ) );
  NOR40 U3288 ( .A(\u_coder/i [5]), .B(\u_coder/i [4]), .C(\u_coder/i [19]), 
        .D(\u_coder/i [18]), .Q(\u_coder/n333 ) );
  NOR40 U3289 ( .A(\u_coder/i [17]), .B(\u_coder/i [16]), .C(\u_coder/i [15]), 
        .D(\u_coder/i [14]), .Q(\u_coder/n332 ) );
  NOR40 U3290 ( .A(n2763), .B(n2764), .C(n2225), .D(n2762), .Q(
        \u_outFIFO/N1270 ) );
  INV3 U3291 ( .A(n2759), .Q(n2225) );
  NAND41 U3292 ( .A(n2757), .B(n2751), .C(n2750), .D(n2747), .Q(n2763) );
  AOI211 U3293 ( .A(\u_outFIFO/outWriteCount[1] ), .B(n2761), .C(n2227), .Q(
        n2762) );
  AOI311 U3294 ( .A(n2759), .B(n2757), .C(n2756), .D(
        \u_outFIFO/outWriteCount[7] ), .Q(n2758) );
  OAI2111 U3295 ( .A(\u_outFIFO/outReadCount[5] ), .B(\u_outFIFO/n261 ), .C(
        n2755), .D(n2754), .Q(n2756) );
  NAND22 U3296 ( .A(\u_outFIFO/outWriteCount[4] ), .B(n196), .Q(n2754) );
  NAND41 U3297 ( .A(n2743), .B(n2742), .C(n2741), .D(n2740), .Q(\u_coder/N668 ) );
  NOR21 U3298 ( .A(\u_coder/i [10]), .B(n763), .Q(n2743) );
  NOR31 U3299 ( .A(\u_coder/i [11]), .B(\u_coder/i [13]), .C(\u_coder/i [12]), 
        .Q(n2742) );
  NOR40 U3300 ( .A(\u_coder/i [16]), .B(n2158), .C(\u_coder/i [15]), .D(
        \u_coder/i [14]), .Q(n2741) );
  NAND41 U3301 ( .A(n2734), .B(n2733), .C(n2732), .D(n2731), .Q(\u_coder/N974 ) );
  NOR21 U3302 ( .A(\u_coder/j [10]), .B(\u_coder/j [0]), .Q(n2734) );
  NOR31 U3303 ( .A(\u_coder/j [11]), .B(\u_coder/j [13]), .C(\u_coder/j [12]), 
        .Q(n2733) );
  NOR40 U3304 ( .A(\u_coder/j [16]), .B(n2171), .C(\u_coder/j [15]), .D(
        \u_coder/j [14]), .Q(n2732) );
  INV3 U3305 ( .A(\u_coder/n326 ), .Q(n2177) );
  NAND41 U3306 ( .A(\u_coder/n327 ), .B(\u_coder/n328 ), .C(\u_coder/n329 ), 
        .D(\u_coder/n330 ), .Q(\u_coder/n326 ) );
  NOR40 U3307 ( .A(\u_coder/j [9]), .B(\u_coder/j [8]), .C(\u_coder/j [7]), 
        .D(\u_coder/j [6]), .Q(\u_coder/n330 ) );
  NOR40 U3308 ( .A(\u_coder/j [5]), .B(\u_coder/j [4]), .C(\u_coder/j [19]), 
        .D(\u_coder/j [18]), .Q(\u_coder/n329 ) );
  NOR40 U3309 ( .A(\u_coder/j [13]), .B(\u_coder/j [12]), .C(\u_coder/j [11]), 
        .D(\u_coder/j [10]), .Q(\u_coder/n327 ) );
  NOR40 U3310 ( .A(\u_coder/i [13]), .B(\u_coder/i [12]), .C(\u_coder/i [11]), 
        .D(\u_coder/i [10]), .Q(\u_coder/n331 ) );
  NAND31 U3311 ( .A(\u_cdr/div1/n7 ), .B(\u_cdr/w_nb_P [4]), .C(n1242), .Q(
        n1243) );
  OAI311 U3312 ( .A(n1243), .B(\u_cdr/div1/n8 ), .C(\u_cdr/w_nb_P [2]), .D(
        \u_cdr/w_sE ), .Q(n1261) );
  NAND22 U3313 ( .A(\u_coder/N668 ), .B(\u_coder/isPositiveI ), .Q(
        \u_coder/n147 ) );
  NAND22 U3314 ( .A(\u_coder/N974 ), .B(\u_coder/n127 ), .Q(\u_coder/n192 ) );
  OAI311 U3315 ( .A(n1243), .B(\u_cdr/div1/n9 ), .C(\u_cdr/w_nb_P [3]), .D(
        n221), .Q(n1257) );
  NOR31 U3316 ( .A(\u_coder/n103 ), .B(\u_coder/n256 ), .C(\u_coder/n312 ), 
        .Q(\u_coder/n246 ) );
  NAND31 U3317 ( .A(\u_coder/n105 ), .B(\u_coder/n101 ), .C(\u_coder/n104 ), 
        .Q(\u_coder/n312 ) );
  NOR40 U3318 ( .A(n2739), .B(n2164), .C(\u_coder/i [1]), .D(\u_coder/i [19]), 
        .Q(n2740) );
  INV3 U3319 ( .A(n2738), .Q(n2164) );
  NAND22 U3320 ( .A(n2737), .B(n2736), .Q(n2739) );
  NOR31 U3321 ( .A(\u_coder/i [2]), .B(\u_coder/i [4]), .C(\u_coder/i [3]), 
        .Q(n2738) );
  NAND22 U3322 ( .A(\u_inFIFO/n215 ), .B(\u_inFIFO/n176 ), .Q(\u_inFIFO/n520 )
         );
  NOR40 U3323 ( .A(n2730), .B(n2179), .C(n762), .D(\u_coder/j [19]), .Q(n2731)
         );
  NAND22 U3324 ( .A(n2728), .B(n2727), .Q(n2730) );
  INV3 U3325 ( .A(n2729), .Q(n2179) );
  NOR21 U3326 ( .A(\u_coder/j [6]), .B(\u_coder/j [5]), .Q(n2728) );
  NOR21 U3327 ( .A(\u_decoder/fir_filter/state [1]), .B(
        \u_decoder/fir_filter/state [0]), .Q(\u_decoder/fir_filter/n1149 ) );
  INV3 U3328 ( .A(\u_inFIFO/n554 ), .Q(n1821) );
  AOI221 U3329 ( .A(\u_inFIFO/N124 ), .B(n2094), .C(\u_inFIFO/outReadCount[6] ), .D(\u_inFIFO/n542 ), .Q(\u_inFIFO/n554 ) );
  XOR21 U3330 ( .A(\u_inFIFO/add_252/carry [6]), .B(\u_inFIFO/outReadCount[6] ), .Q(\u_inFIFO/N124 ) );
  INV3 U3331 ( .A(\u_inFIFO/n541 ), .Q(n1827) );
  AOI221 U3332 ( .A(\u_inFIFO/N123 ), .B(n2094), .C(\u_inFIFO/outReadCount[5] ), .D(\u_inFIFO/n542 ), .Q(\u_inFIFO/n541 ) );
  INV3 U3333 ( .A(\u_inFIFO/n512 ), .Q(n1965) );
  AOI221 U3334 ( .A(\u_inFIFO/N217 ), .B(\u_inFIFO/n513 ), .C(n1211), .D(
        \u_inFIFO/j_FIFO [6]), .Q(\u_inFIFO/n512 ) );
  XOR21 U3335 ( .A(\u_inFIFO/add_357/carry [6]), .B(\u_inFIFO/j_FIFO [6]), .Q(
        \u_inFIFO/N217 ) );
  INV3 U3336 ( .A(\u_outFIFO/n676 ), .Q(n1588) );
  INV3 U3337 ( .A(\u_outFIFO/n673 ), .Q(n1587) );
  INV3 U3338 ( .A(\u_inFIFO/n515 ), .Q(n1963) );
  AOI221 U3339 ( .A(\u_inFIFO/N215 ), .B(\u_inFIFO/n513 ), .C(n1211), .D(
        \u_inFIFO/j_FIFO [4]), .Q(\u_inFIFO/n515 ) );
  INV3 U3340 ( .A(\u_outFIFO/n1121 ), .Q(n1803) );
  AOI221 U3341 ( .A(\u_outFIFO/N140 ), .B(\u_outFIFO/n1119 ), .C(
        \u_outFIFO/outReadCount[5] ), .D(\u_outFIFO/n1120 ), .Q(
        \u_outFIFO/n1121 ) );
  INV3 U3342 ( .A(\u_inFIFO/n519 ), .Q(n1959) );
  AOI221 U3343 ( .A(\u_inFIFO/n207 ), .B(\u_inFIFO/n513 ), .C(n1211), .D(
        \u_inFIFO/j_FIFO [0]), .Q(\u_inFIFO/n519 ) );
  INV3 U3344 ( .A(\u_cordic/mycordic/n479 ), .Q(n1529) );
  AOI221 U3345 ( .A(\u_cordic/mycordic/N464 ), .B(n777), .C(
        \u_cordic/mycordic/N492 ), .D(n1907), .Q(\u_cordic/mycordic/n479 ) );
  XNR21 U3346 ( .A(\u_cordic/mycordic/present_ANGLE_table[3][8] ), .B(
        \u_cordic/mycordic/sub_218/carry[8] ), .Q(\u_cordic/mycordic/N492 ) );
  XOR21 U3347 ( .A(\u_cordic/mycordic/present_ANGLE_table[3][8] ), .B(
        \u_cordic/mycordic/add_213/carry[8] ), .Q(\u_cordic/mycordic/N464 ) );
  INV3 U3348 ( .A(\u_cordic/mycordic/n478 ), .Q(n1530) );
  AOI221 U3349 ( .A(\u_cordic/mycordic/N465 ), .B(\u_cordic/mycordic/n363 ), 
        .C(\u_cordic/mycordic/N493 ), .D(n1907), .Q(\u_cordic/mycordic/n478 )
         );
  XNR21 U3350 ( .A(\u_cordic/mycordic/present_ANGLE_table[3][9] ), .B(
        \u_cordic/mycordic/sub_218/carry[9] ), .Q(\u_cordic/mycordic/N493 ) );
  XOR21 U3351 ( .A(\u_cordic/mycordic/present_ANGLE_table[3][9] ), .B(
        \u_cordic/mycordic/add_213/carry[9] ), .Q(\u_cordic/mycordic/N465 ) );
  INV3 U3352 ( .A(\u_decoder/fir_filter/n1076 ), .Q(n2270) );
  AOI221 U3353 ( .A(\u_decoder/fir_filter/I_data_mult_4 [6]), .B(n1091), .C(
        \u_decoder/fir_filter/I_data_mult_4_buff [6]), .D(n1164), .Q(
        \u_decoder/fir_filter/n1076 ) );
  INV3 U3354 ( .A(\u_decoder/fir_filter/n1073 ), .Q(n2273) );
  AOI221 U3355 ( .A(\u_decoder/fir_filter/I_data_mult_4 [3]), .B(n1091), .C(
        \u_decoder/fir_filter/I_data_mult_4_buff [3]), .D(n1164), .Q(
        \u_decoder/fir_filter/n1073 ) );
  XOR21 U3356 ( .A(n8), .B(\u_decoder/fir_filter/I_data_mult_0 [0]), .Q(
        \u_decoder/fir_filter/I_data_mult_4 [3]) );
  INV3 U3357 ( .A(\u_decoder/fir_filter/n1071 ), .Q(n2298) );
  AOI221 U3358 ( .A(n12), .B(n1091), .C(
        \u_decoder/fir_filter/I_data_mult_4_buff [1]), .D(n1164), .Q(
        \u_decoder/fir_filter/n1071 ) );
  INV3 U3359 ( .A(\u_decoder/fir_filter/n1070 ), .Q(n2255) );
  AOI221 U3360 ( .A(\u_decoder/fir_filter/I_data_mult_0 [0]), .B(n1091), .C(
        \u_decoder/fir_filter/I_data_mult_4_buff [0]), .D(n1164), .Q(
        \u_decoder/fir_filter/n1070 ) );
  INV3 U3361 ( .A(\u_decoder/fir_filter/n996 ), .Q(n2636) );
  AOI221 U3362 ( .A(\u_decoder/fir_filter/I_data_add_7 [0]), .B(n1091), .C(
        \u_decoder/fir_filter/I_data_add_7_buff [0]), .D(n1164), .Q(
        \u_decoder/fir_filter/n996 ) );
  XOR21 U3363 ( .A(\u_decoder/fir_filter/I_data_mult_7_buff [0]), .B(
        \u_decoder/fir_filter/I_data_mult_8_buff [0]), .Q(
        \u_decoder/fir_filter/I_data_add_7 [0]) );
  INV3 U3364 ( .A(\u_decoder/fir_filter/n975 ), .Q(n2621) );
  AOI221 U3365 ( .A(\u_decoder/fir_filter/I_data_add_6 [0]), .B(n1092), .C(
        \u_decoder/fir_filter/I_data_add_6_buff [0]), .D(n1165), .Q(
        \u_decoder/fir_filter/n975 ) );
  XOR21 U3366 ( .A(\u_decoder/fir_filter/I_data_mult_6_buff [0]), .B(
        \u_decoder/fir_filter/I_data_add_7_buff [0]), .Q(
        \u_decoder/fir_filter/I_data_add_6 [0]) );
  INV3 U3367 ( .A(\u_decoder/fir_filter/n954 ), .Q(n2606) );
  AOI221 U3368 ( .A(\u_decoder/fir_filter/I_data_add_5 [0]), .B(n1093), .C(
        \u_decoder/fir_filter/I_data_add_5_buff [0]), .D(n1166), .Q(
        \u_decoder/fir_filter/n954 ) );
  XOR21 U3369 ( .A(\u_decoder/fir_filter/I_data_mult_5_buff [0]), .B(
        \u_decoder/fir_filter/I_data_add_6_buff [0]), .Q(
        \u_decoder/fir_filter/I_data_add_5 [0]) );
  INV3 U3370 ( .A(\u_decoder/fir_filter/n933 ), .Q(n2591) );
  AOI221 U3371 ( .A(\u_decoder/fir_filter/I_data_add_4 [0]), .B(n1094), .C(
        \u_decoder/fir_filter/I_data_add_4_buff [0]), .D(n1166), .Q(
        \u_decoder/fir_filter/n933 ) );
  XOR21 U3372 ( .A(\u_decoder/fir_filter/I_data_mult_4_buff [0]), .B(
        \u_decoder/fir_filter/I_data_add_5_buff [0]), .Q(
        \u_decoder/fir_filter/I_data_add_4 [0]) );
  INV3 U3373 ( .A(\u_decoder/fir_filter/n932 ), .Q(n2590) );
  AOI221 U3374 ( .A(\u_decoder/fir_filter/I_data_add_4 [1]), .B(n1094), .C(
        \u_decoder/fir_filter/I_data_add_4_buff [1]), .D(n1166), .Q(
        \u_decoder/fir_filter/n932 ) );
  INV3 U3375 ( .A(\u_decoder/fir_filter/n677 ), .Q(n2501) );
  AOI221 U3376 ( .A(\u_decoder/fir_filter/Q_data_add_6 [0]), .B(n1085), .C(
        \u_decoder/fir_filter/Q_data_add_6_buff [0]), .D(n1161), .Q(
        \u_decoder/fir_filter/n677 ) );
  XOR21 U3377 ( .A(\u_decoder/fir_filter/Q_data_mult_6_buff [0]), .B(
        \u_decoder/fir_filter/Q_data_add_7_buff [0]), .Q(
        \u_decoder/fir_filter/Q_data_add_6 [0]) );
  INV3 U3378 ( .A(\u_decoder/fir_filter/n656 ), .Q(n2486) );
  AOI221 U3379 ( .A(\u_decoder/fir_filter/Q_data_add_5 [0]), .B(n1086), .C(
        \u_decoder/fir_filter/Q_data_add_5_buff [0]), .D(n1157), .Q(
        \u_decoder/fir_filter/n656 ) );
  XOR21 U3380 ( .A(\u_decoder/fir_filter/Q_data_mult_5_buff [0]), .B(
        \u_decoder/fir_filter/Q_data_add_6_buff [0]), .Q(
        \u_decoder/fir_filter/Q_data_add_5 [0]) );
  INV3 U3381 ( .A(\u_decoder/fir_filter/n635 ), .Q(n2471) );
  AOI221 U3382 ( .A(\u_decoder/fir_filter/Q_data_add_4 [0]), .B(n1087), .C(
        \u_decoder/fir_filter/Q_data_add_4_buff [0]), .D(n1165), .Q(
        \u_decoder/fir_filter/n635 ) );
  XOR21 U3383 ( .A(\u_decoder/fir_filter/Q_data_mult_4_buff [0]), .B(
        \u_decoder/fir_filter/Q_data_add_5_buff [0]), .Q(
        \u_decoder/fir_filter/Q_data_add_4 [0]) );
  INV3 U3384 ( .A(\u_decoder/fir_filter/n634 ), .Q(n2470) );
  AOI221 U3385 ( .A(\u_decoder/fir_filter/Q_data_add_4 [1]), .B(n1087), .C(
        \u_decoder/fir_filter/Q_data_add_4_buff [1]), .D(n1160), .Q(
        \u_decoder/fir_filter/n634 ) );
  INV3 U3386 ( .A(\u_decoder/fir_filter/n633 ), .Q(n2469) );
  AOI221 U3387 ( .A(\u_decoder/fir_filter/Q_data_add_4 [2]), .B(n1087), .C(
        \u_decoder/fir_filter/Q_data_add_4_buff [2]), .D(n1154), .Q(
        \u_decoder/fir_filter/n633 ) );
  INV3 U3388 ( .A(\u_decoder/fir_filter/n632 ), .Q(n2468) );
  AOI221 U3389 ( .A(\u_decoder/fir_filter/Q_data_add_4 [3]), .B(n1087), .C(
        \u_decoder/fir_filter/Q_data_add_4_buff [3]), .D(n1153), .Q(
        \u_decoder/fir_filter/n632 ) );
  INV3 U3390 ( .A(\u_decoder/fir_filter/n631 ), .Q(n2467) );
  AOI221 U3391 ( .A(\u_decoder/fir_filter/Q_data_add_4 [4]), .B(n1087), .C(
        \u_decoder/fir_filter/Q_data_add_4_buff [4]), .D(n1152), .Q(
        \u_decoder/fir_filter/n631 ) );
  INV3 U3392 ( .A(\u_decoder/fir_filter/n630 ), .Q(n2466) );
  AOI221 U3393 ( .A(\u_decoder/fir_filter/Q_data_add_4 [5]), .B(n1087), .C(
        \u_decoder/fir_filter/Q_data_add_4_buff [5]), .D(n1162), .Q(
        \u_decoder/fir_filter/n630 ) );
  INV3 U3394 ( .A(\u_decoder/fir_filter/n629 ), .Q(n2465) );
  AOI221 U3395 ( .A(\u_decoder/fir_filter/Q_data_add_4 [6]), .B(n1087), .C(
        \u_decoder/fir_filter/Q_data_add_4_buff [6]), .D(n1162), .Q(
        \u_decoder/fir_filter/n629 ) );
  INV3 U3396 ( .A(\u_decoder/fir_filter/n614 ), .Q(n2456) );
  AOI221 U3397 ( .A(\u_decoder/fir_filter/Q_data_add_3 [0]), .B(n1087), .C(
        \u_decoder/fir_filter/Q_data_add_3_buff [0]), .D(n1162), .Q(
        \u_decoder/fir_filter/n614 ) );
  XOR21 U3398 ( .A(\u_decoder/fir_filter/Q_data_mult_3_buff [0]), .B(
        \u_decoder/fir_filter/Q_data_add_4_buff [0]), .Q(
        \u_decoder/fir_filter/Q_data_add_3 [0]) );
  INV3 U3399 ( .A(\u_decoder/fir_filter/n593 ), .Q(n2441) );
  AOI221 U3400 ( .A(\u_decoder/fir_filter/Q_data_add_2 [0]), .B(n1088), .C(
        \u_decoder/fir_filter/Q_data_add_2_buff [0]), .D(n1161), .Q(
        \u_decoder/fir_filter/n593 ) );
  XOR21 U3401 ( .A(\u_decoder/fir_filter/Q_data_mult_2_buff [0]), .B(
        \u_decoder/fir_filter/Q_data_add_3_buff [0]), .Q(
        \u_decoder/fir_filter/Q_data_add_2 [0]) );
  INV3 U3402 ( .A(\u_decoder/fir_filter/n931 ), .Q(n2589) );
  AOI221 U3403 ( .A(\u_decoder/fir_filter/I_data_add_4 [2]), .B(n1094), .C(
        \u_decoder/fir_filter/I_data_add_4_buff [2]), .D(n1156), .Q(
        \u_decoder/fir_filter/n931 ) );
  INV3 U3404 ( .A(\u_decoder/fir_filter/n930 ), .Q(n2588) );
  AOI221 U3405 ( .A(\u_decoder/fir_filter/I_data_add_4 [3]), .B(n1094), .C(
        \u_decoder/fir_filter/I_data_add_4_buff [3]), .D(n1155), .Q(
        \u_decoder/fir_filter/n930 ) );
  INV3 U3406 ( .A(\u_decoder/fir_filter/n929 ), .Q(n2587) );
  AOI221 U3407 ( .A(\u_decoder/fir_filter/I_data_add_4 [4]), .B(n1094), .C(
        \u_decoder/fir_filter/I_data_add_4_buff [4]), .D(n1158), .Q(
        \u_decoder/fir_filter/n929 ) );
  INV3 U3408 ( .A(\u_decoder/fir_filter/n928 ), .Q(n2586) );
  AOI221 U3409 ( .A(\u_decoder/fir_filter/I_data_add_4 [5]), .B(n1094), .C(
        \u_decoder/fir_filter/I_data_add_4_buff [5]), .D(n1154), .Q(
        \u_decoder/fir_filter/n928 ) );
  INV3 U3410 ( .A(\u_decoder/fir_filter/n927 ), .Q(n2585) );
  AOI221 U3411 ( .A(\u_decoder/fir_filter/I_data_add_4 [6]), .B(n1094), .C(
        \u_decoder/fir_filter/I_data_add_4_buff [6]), .D(n1153), .Q(
        \u_decoder/fir_filter/n927 ) );
  INV3 U3412 ( .A(\u_decoder/fir_filter/n912 ), .Q(n2576) );
  AOI221 U3413 ( .A(\u_decoder/fir_filter/I_data_add_3 [0]), .B(n1095), .C(
        \u_decoder/fir_filter/I_data_add_3_buff [0]), .D(n1162), .Q(
        \u_decoder/fir_filter/n912 ) );
  XOR21 U3414 ( .A(\u_decoder/fir_filter/I_data_mult_3_buff [0]), .B(
        \u_decoder/fir_filter/I_data_add_4_buff [0]), .Q(
        \u_decoder/fir_filter/I_data_add_3 [0]) );
  INV3 U3415 ( .A(\u_decoder/fir_filter/n891 ), .Q(n2561) );
  AOI221 U3416 ( .A(\u_decoder/fir_filter/I_data_add_2 [0]), .B(n1096), .C(
        \u_decoder/fir_filter/I_data_add_2_buff [0]), .D(n1158), .Q(
        \u_decoder/fir_filter/n891 ) );
  XOR21 U3417 ( .A(\u_decoder/fir_filter/I_data_mult_2_buff [0]), .B(
        \u_decoder/fir_filter/I_data_add_3_buff [0]), .Q(
        \u_decoder/fir_filter/I_data_add_2 [0]) );
  INV3 U3418 ( .A(\u_decoder/fir_filter/n870 ), .Q(n2546) );
  AOI221 U3419 ( .A(\u_decoder/fir_filter/I_data_add_1 [0]), .B(n1096), .C(
        \u_decoder/fir_filter/I_data_add_1_buff [0]), .D(n1156), .Q(
        \u_decoder/fir_filter/n870 ) );
  XOR21 U3420 ( .A(\u_decoder/fir_filter/I_data_mult_1_buff [0]), .B(
        \u_decoder/fir_filter/I_data_add_2_buff [0]), .Q(
        \u_decoder/fir_filter/I_data_add_1 [0]) );
  INV3 U3421 ( .A(\u_decoder/fir_filter/n779 ), .Q(n2341) );
  AOI221 U3422 ( .A(\u_decoder/fir_filter/Q_data_mult_4 [6]), .B(n1083), .C(
        \u_decoder/fir_filter/Q_data_mult_4_buff [6]), .D(n1164), .Q(
        \u_decoder/fir_filter/n779 ) );
  NOR31 U3423 ( .A(\u_coder/j [2]), .B(\u_coder/j [4]), .C(\u_coder/j [3]), 
        .Q(n2729) );
  INV3 U3424 ( .A(\u_decoder/fir_filter/n698 ), .Q(n2516) );
  AOI221 U3425 ( .A(\u_decoder/fir_filter/Q_data_add_7 [0]), .B(n1084), .C(
        \u_decoder/fir_filter/Q_data_add_7_buff [0]), .D(n1161), .Q(
        \u_decoder/fir_filter/n698 ) );
  XOR21 U3426 ( .A(\u_decoder/fir_filter/Q_data_mult_7_buff [0]), .B(
        \u_decoder/fir_filter/Q_data_mult_8_buff [0]), .Q(
        \u_decoder/fir_filter/Q_data_add_7 [0]) );
  INV3 U3427 ( .A(\u_decoder/fir_filter/n572 ), .Q(n2426) );
  AOI221 U3428 ( .A(\u_decoder/fir_filter/Q_data_add_1 [0]), .B(n1089), .C(
        \u_decoder/fir_filter/Q_data_add_1_buff [0]), .D(n1160), .Q(
        \u_decoder/fir_filter/n572 ) );
  XOR21 U3429 ( .A(\u_decoder/fir_filter/Q_data_mult_1_buff [0]), .B(
        \u_decoder/fir_filter/Q_data_add_2_buff [0]), .Q(
        \u_decoder/fir_filter/Q_data_add_1 [0]) );
  INV3 U3430 ( .A(\u_cordic/mycordic/n441 ), .Q(n1449) );
  AOI221 U3431 ( .A(\u_cordic/mycordic/N546 ), .B(n770), .C(
        \u_cordic/mycordic/N562 ), .D(n1903), .Q(\u_cordic/mycordic/n441 ) );
  XNR21 U3432 ( .A(\u_cordic/mycordic/present_ANGLE_table[5][12] ), .B(
        \u_cordic/mycordic/sub_236/carry [12]), .Q(\u_cordic/mycordic/N562 )
         );
  XOR21 U3433 ( .A(\u_cordic/mycordic/present_ANGLE_table[5][12] ), .B(
        \u_cordic/mycordic/add_233/carry [12]), .Q(\u_cordic/mycordic/N546 )
         );
  INV3 U3434 ( .A(\u_decoder/fir_filter/n776 ), .Q(n2344) );
  AOI221 U3435 ( .A(\u_decoder/fir_filter/Q_data_mult_4 [3]), .B(n1084), .C(
        \u_decoder/fir_filter/Q_data_mult_4_buff [3]), .D(n1157), .Q(
        \u_decoder/fir_filter/n776 ) );
  XOR21 U3436 ( .A(n7), .B(\u_decoder/fir_filter/Q_data_mult_0 [0]), .Q(
        \u_decoder/fir_filter/Q_data_mult_4 [3]) );
  INV3 U3437 ( .A(\u_decoder/fir_filter/n774 ), .Q(n2369) );
  AOI221 U3438 ( .A(n11), .B(n1084), .C(
        \u_decoder/fir_filter/Q_data_mult_4_buff [1]), .D(n1159), .Q(
        \u_decoder/fir_filter/n774 ) );
  INV3 U3439 ( .A(\u_outFIFO/n681 ), .Q(n1590) );
  INV3 U3440 ( .A(\u_outFIFO/n671 ), .Q(n1586) );
  INV3 U3441 ( .A(\u_outFIFO/n1101 ), .Q(n1789) );
  INV3 U3442 ( .A(\u_outFIFO/n1093 ), .Q(n1785) );
  INV3 U3443 ( .A(\u_outFIFO/n1108 ), .Q(n1792) );
  INV3 U3444 ( .A(\u_outFIFO/n852 ), .Q(n1671) );
  INV3 U3445 ( .A(\u_outFIFO/n723 ), .Q(n1609) );
  INV3 U3446 ( .A(\u_outFIFO/n721 ), .Q(n1608) );
  INV3 U3447 ( .A(\u_outFIFO/n719 ), .Q(n1607) );
  INV3 U3448 ( .A(\u_outFIFO/n900 ), .Q(n1695) );
  INV3 U3449 ( .A(\u_outFIFO/n1084 ), .Q(n1781) );
  INV3 U3450 ( .A(\u_outFIFO/n944 ), .Q(n1717) );
  INV3 U3451 ( .A(\u_outFIFO/n1051 ), .Q(n1765) );
  INV3 U3452 ( .A(\u_outFIFO/n1068 ), .Q(n1773) );
  INV3 U3453 ( .A(\u_outFIFO/n1066 ), .Q(n1772) );
  INV3 U3454 ( .A(\u_outFIFO/n1060 ), .Q(n1769) );
  INV3 U3455 ( .A(\u_outFIFO/n1058 ), .Q(n1768) );
  INV3 U3456 ( .A(\u_outFIFO/n1027 ), .Q(n1753) );
  INV3 U3457 ( .A(\u_outFIFO/n1025 ), .Q(n1752) );
  INV3 U3458 ( .A(\u_outFIFO/n896 ), .Q(n1693) );
  INV3 U3459 ( .A(\u_outFIFO/n894 ), .Q(n1692) );
  INV3 U3460 ( .A(\u_outFIFO/n888 ), .Q(n1689) );
  INV3 U3461 ( .A(\u_outFIFO/n886 ), .Q(n1688) );
  INV3 U3462 ( .A(\u_outFIFO/n967 ), .Q(n1728) );
  INV3 U3463 ( .A(\u_outFIFO/n958 ), .Q(n1724) );
  INV3 U3464 ( .A(\u_outFIFO/n950 ), .Q(n1720) );
  INV3 U3465 ( .A(\u_outFIFO/n942 ), .Q(n1716) );
  INV3 U3466 ( .A(\u_outFIFO/n834 ), .Q(n1664) );
  INV3 U3467 ( .A(\u_outFIFO/n825 ), .Q(n1660) );
  INV3 U3468 ( .A(\u_outFIFO/n817 ), .Q(n1656) );
  INV3 U3469 ( .A(\u_outFIFO/n809 ), .Q(n1652) );
  INV3 U3470 ( .A(\u_cordic/mycordic/n344 ), .Q(n1495) );
  AOI221 U3471 ( .A(n1905), .B(\u_cordic/mycordic/N259 ), .C(n774), .D(
        \u_cordic/mycordic/N267 ), .Q(\u_cordic/mycordic/n344 ) );
  INV3 U3472 ( .A(\u_outFIFO/n1000 ), .Q(n1741) );
  INV3 U3473 ( .A(\u_outFIFO/n998 ), .Q(n1740) );
  INV3 U3474 ( .A(\u_outFIFO/n731 ), .Q(n1613) );
  INV3 U3475 ( .A(\u_outFIFO/n1007 ), .Q(n1744) );
  INV3 U3476 ( .A(\u_outFIFO/n977 ), .Q(n1732) );
  INV3 U3477 ( .A(\u_outFIFO/n870 ), .Q(n1680) );
  INV3 U3478 ( .A(\u_outFIFO/n868 ), .Q(n1679) );
  INV3 U3479 ( .A(\u_outFIFO/n844 ), .Q(n1668) );
  INV3 U3480 ( .A(\u_outFIFO/n841 ), .Q(n1667) );
  INV3 U3481 ( .A(\u_outFIFO/n737 ), .Q(n1616) );
  INV3 U3482 ( .A(\u_outFIFO/n735 ), .Q(n1615) );
  INV3 U3483 ( .A(\u_outFIFO/n711 ), .Q(n1604) );
  INV3 U3484 ( .A(\u_outFIFO/n708 ), .Q(n1603) );
  NAND22 U3485 ( .A(\u_decoder/fir_filter/state [1]), .B(
        \u_decoder/fir_filter/n410 ), .Q(\u_decoder/fir_filter/n1153 ) );
  INV3 U3486 ( .A(\u_outFIFO/N219 ), .Q(n2213) );
  INV3 U3487 ( .A(\u_outFIFO/N220 ), .Q(n2212) );
  NAND22 U3488 ( .A(\u_coder/N668 ), .B(\u_coder/n126 ), .Q(\u_coder/n158 ) );
  INV3 U3489 ( .A(\u_outFIFO/N132 ), .Q(n2232) );
  XNR21 U3490 ( .A(\u_outFIFO/add_256/carry [6]), .B(\u_outFIFO/i_FIFO [6]), 
        .Q(n376) );
  NAND22 U3491 ( .A(\u_outFIFO/currentState [0]), .B(\u_outFIFO/n256 ), .Q(
        \u_outFIFO/n308 ) );
  XNR21 U3492 ( .A(\u_cordic/mycordic/r173/carry [10]), .B(
        \u_cordic/mycordic/present_ANGLE_table[6][10] ), .Q(n377) );
  XNR21 U3493 ( .A(\u_cordic/mycordic/r173/carry [11]), .B(
        \u_cordic/mycordic/present_ANGLE_table[6][11] ), .Q(n378) );
  OAI2111 U3494 ( .A(n2753), .B(n2752), .C(n2751), .D(n2750), .Q(n2755) );
  NOR21 U3495 ( .A(\u_outFIFO/outReadCount[3] ), .B(\u_outFIFO/n263 ), .Q(
        n2753) );
  OAI2111 U3496 ( .A(n2748), .B(n161), .C(n2226), .D(n2747), .Q(n2749) );
  NAND22 U3497 ( .A(\u_coder/N974 ), .B(\u_coder/isPositiveQ ), .Q(
        \u_coder/n217 ) );
  NOR21 U3498 ( .A(\u_inFIFO/n173 ), .B(\u_inFIFO/currentState [3]), .Q(
        \u_inFIFO/n215 ) );
  NAND22 U3499 ( .A(\u_outFIFO/currentState [2]), .B(\u_outFIFO/n253 ), .Q(
        \u_outFIFO/n1159 ) );
  NOR31 U3500 ( .A(\u_coder/i [7]), .B(\u_coder/i [9]), .C(\u_coder/i [8]), 
        .Q(n2736) );
  NOR31 U3501 ( .A(\u_coder/j [7]), .B(\u_coder/j [9]), .C(\u_coder/j [8]), 
        .Q(n2727) );
  XOR21 U3502 ( .A(\u_cordic/mycordic/add_262/carry [10]), .B(
        \u_cordic/mycordic/present_ANGLE_table[6][10] ), .Q(
        \u_cordic/mycordic/N625 ) );
  XOR21 U3503 ( .A(\u_cordic/mycordic/add_262/carry [11]), .B(
        \u_cordic/mycordic/present_ANGLE_table[6][11] ), .Q(
        \u_cordic/mycordic/N626 ) );
  XOR21 U3504 ( .A(\u_cordic/mycordic/add_262/carry [13]), .B(
        \u_cordic/mycordic/present_ANGLE_table[6][13] ), .Q(
        \u_cordic/mycordic/N628 ) );
  NAND22 U3505 ( .A(\u_inFIFO/outReadCount[0] ), .B(\u_inFIFO/n188 ), .Q(n2708) );
  NAND22 U3506 ( .A(\u_inFIFO/outReadCount[6] ), .B(\u_inFIFO/n182 ), .Q(n2706) );
  NAND22 U3507 ( .A(\u_inFIFO/outReadCount[5] ), .B(\u_inFIFO/n183 ), .Q(n2704) );
  NAND22 U3508 ( .A(\u_decoder/fir_filter/I_data_mult_1_buff [5]), .B(n1160), 
        .Q(\u_decoder/fir_filter/n1123 ) );
  NAND22 U3509 ( .A(\u_decoder/fir_filter/I_data_mult_7_buff [5]), .B(n1156), 
        .Q(\u_decoder/fir_filter/n1025 ) );
  NAND22 U3510 ( .A(\u_decoder/fir_filter/Q_data_mult_1_buff [5]), .B(n1152), 
        .Q(\u_decoder/fir_filter/n826 ) );
  NAND22 U3511 ( .A(\u_decoder/fir_filter/Q_data_mult_7_buff [5]), .B(n1153), 
        .Q(\u_decoder/fir_filter/n728 ) );
  NAND22 U3512 ( .A(\u_decoder/fir_filter/I_data_mult_0_buff [4]), .B(n1160), 
        .Q(\u_decoder/fir_filter/n1138 ) );
  NAND22 U3513 ( .A(\u_decoder/fir_filter/Q_data_mult_0_buff [4]), .B(n1152), 
        .Q(\u_decoder/fir_filter/n841 ) );
  NAND22 U3514 ( .A(\u_decoder/fir_filter/I_data_mult_0_buff [1]), .B(n1160), 
        .Q(\u_decoder/fir_filter/n1135 ) );
  NAND22 U3515 ( .A(\u_decoder/fir_filter/I_data_mult_1_buff [1]), .B(n1159), 
        .Q(\u_decoder/fir_filter/n1119 ) );
  NAND22 U3516 ( .A(\u_decoder/fir_filter/I_data_mult_2_buff [2]), .B(n1158), 
        .Q(\u_decoder/fir_filter/n1104 ) );
  NAND22 U3517 ( .A(\u_decoder/fir_filter/I_data_mult_6_buff [2]), .B(n1157), 
        .Q(\u_decoder/fir_filter/n1039 ) );
  NAND22 U3518 ( .A(\u_decoder/fir_filter/I_data_mult_7_buff [1]), .B(n1166), 
        .Q(\u_decoder/fir_filter/n1021 ) );
  NAND22 U3519 ( .A(\u_decoder/fir_filter/Q_data_mult_0_buff [1]), .B(n1162), 
        .Q(\u_decoder/fir_filter/n838 ) );
  NAND22 U3520 ( .A(\u_decoder/fir_filter/Q_data_mult_1_buff [1]), .B(n1152), 
        .Q(\u_decoder/fir_filter/n822 ) );
  NAND22 U3521 ( .A(\u_decoder/fir_filter/Q_data_mult_2_buff [2]), .B(n1156), 
        .Q(\u_decoder/fir_filter/n807 ) );
  NAND22 U3522 ( .A(\u_decoder/fir_filter/Q_data_mult_6_buff [2]), .B(n1156), 
        .Q(\u_decoder/fir_filter/n742 ) );
  NAND22 U3523 ( .A(\u_decoder/fir_filter/Q_data_mult_7_buff [1]), .B(n1153), 
        .Q(\u_decoder/fir_filter/n724 ) );
  AOI221 U3524 ( .A(\u_outFIFO/N125 ), .B(n1912), .C(\u_outFIFO/N149 ), .D(
        \u_outFIFO/n1131 ), .Q(\u_outFIFO/n1130 ) );
  AOI221 U3525 ( .A(\u_outFIFO/N123 ), .B(n1912), .C(\u_outFIFO/N147 ), .D(
        \u_outFIFO/n1131 ), .Q(\u_outFIFO/n1133 ) );
  AOI221 U3526 ( .A(\u_outFIFO/N124 ), .B(n1912), .C(\u_outFIFO/N148 ), .D(
        \u_outFIFO/n1131 ), .Q(\u_outFIFO/n1132 ) );
  INV3 U3527 ( .A(\u_cordic/mycordic/n508 ), .Q(n1464) );
  AOI221 U3528 ( .A(\u_cordic/mycordic/N343 ), .B(\u_cordic/mycordic/n336 ), 
        .C(\u_cordic/mycordic/N375 ), .D(n1904), .Q(\u_cordic/mycordic/n508 )
         );
  XNR21 U3529 ( .A(\u_cordic/mycordic/present_ANGLE_table[1][11] ), .B(
        \u_cordic/mycordic/sub_196/carry[11] ), .Q(\u_cordic/mycordic/N375 )
         );
  XOR21 U3530 ( .A(\u_cordic/mycordic/present_ANGLE_table[1][11] ), .B(
        \u_cordic/mycordic/add_191/carry[11] ), .Q(\u_cordic/mycordic/N343 )
         );
  INV3 U3531 ( .A(\u_cordic/mycordic/n477 ), .Q(n1531) );
  AOI221 U3532 ( .A(\u_cordic/mycordic/N466 ), .B(n777), .C(
        \u_cordic/mycordic/N494 ), .D(n1907), .Q(\u_cordic/mycordic/n477 ) );
  XNR21 U3533 ( .A(\u_cordic/mycordic/present_ANGLE_table[3][10] ), .B(
        \u_cordic/mycordic/sub_218/carry[10] ), .Q(\u_cordic/mycordic/N494 )
         );
  XOR21 U3534 ( .A(\u_cordic/mycordic/present_ANGLE_table[3][10] ), .B(
        \u_cordic/mycordic/add_213/carry[10] ), .Q(\u_cordic/mycordic/N466 )
         );
  INV3 U3535 ( .A(\u_cordic/mycordic/n476 ), .Q(n1532) );
  AOI221 U3536 ( .A(\u_cordic/mycordic/N467 ), .B(\u_cordic/mycordic/n363 ), 
        .C(\u_cordic/mycordic/N495 ), .D(n1907), .Q(\u_cordic/mycordic/n476 )
         );
  XNR21 U3537 ( .A(\u_cordic/mycordic/present_ANGLE_table[3][11] ), .B(
        \u_cordic/mycordic/sub_218/carry[11] ), .Q(\u_cordic/mycordic/N495 )
         );
  XOR21 U3538 ( .A(\u_cordic/mycordic/present_ANGLE_table[3][11] ), .B(
        \u_cordic/mycordic/add_213/carry[11] ), .Q(\u_cordic/mycordic/N467 )
         );
  INV3 U3539 ( .A(\u_cordic/mycordic/n444 ), .Q(n1446) );
  AOI221 U3540 ( .A(\u_cordic/mycordic/N543 ), .B(n771), .C(
        \u_cordic/mycordic/N559 ), .D(n1903), .Q(\u_cordic/mycordic/n444 ) );
  XNR21 U3541 ( .A(\u_cordic/mycordic/present_ANGLE_table[5][9] ), .B(
        \u_cordic/mycordic/sub_236/carry [9]), .Q(\u_cordic/mycordic/N559 ) );
  XOR21 U3542 ( .A(\u_cordic/mycordic/present_ANGLE_table[5][9] ), .B(
        \u_cordic/mycordic/add_233/carry [9]), .Q(\u_cordic/mycordic/N543 ) );
  INV3 U3543 ( .A(\u_cordic/mycordic/n443 ), .Q(n1447) );
  AOI221 U3544 ( .A(\u_cordic/mycordic/N544 ), .B(n770), .C(
        \u_cordic/mycordic/N560 ), .D(n1903), .Q(\u_cordic/mycordic/n443 ) );
  XNR21 U3545 ( .A(\u_cordic/mycordic/present_ANGLE_table[5][10] ), .B(
        \u_cordic/mycordic/sub_236/carry [10]), .Q(\u_cordic/mycordic/N560 )
         );
  XOR21 U3546 ( .A(\u_cordic/mycordic/present_ANGLE_table[5][10] ), .B(
        \u_cordic/mycordic/add_233/carry [10]), .Q(\u_cordic/mycordic/N544 )
         );
  NAND22 U3547 ( .A(\u_decoder/fir_filter/I_data_mult_1_buff [6]), .B(n1160), 
        .Q(\u_decoder/fir_filter/n1124 ) );
  NAND22 U3548 ( .A(\u_decoder/fir_filter/I_data_mult_7_buff [6]), .B(n1156), 
        .Q(\u_decoder/fir_filter/n1026 ) );
  NAND22 U3549 ( .A(\u_decoder/fir_filter/Q_data_mult_1_buff [6]), .B(n1152), 
        .Q(\u_decoder/fir_filter/n827 ) );
  NAND22 U3550 ( .A(\u_decoder/fir_filter/Q_data_mult_7_buff [6]), .B(n1153), 
        .Q(\u_decoder/fir_filter/n729 ) );
  NAND22 U3551 ( .A(\u_decoder/fir_filter/I_data_mult_0_buff [5]), .B(n1157), 
        .Q(\u_decoder/fir_filter/n1139 ) );
  NAND22 U3552 ( .A(\u_decoder/fir_filter/Q_data_mult_0_buff [5]), .B(n1151), 
        .Q(\u_decoder/fir_filter/n842 ) );
  AOI221 U3553 ( .A(\u_inFIFO/N148 ), .B(\u_inFIFO/n533 ), .C(\u_inFIFO/N139 ), 
        .D(\u_inFIFO/n534 ), .Q(\u_inFIFO/n539 ) );
  AOI221 U3554 ( .A(\u_inFIFO/N146 ), .B(\u_inFIFO/n533 ), .C(\u_inFIFO/N137 ), 
        .D(\u_inFIFO/n534 ), .Q(\u_inFIFO/n537 ) );
  AOI221 U3555 ( .A(\u_inFIFO/N147 ), .B(\u_inFIFO/n533 ), .C(\u_inFIFO/N138 ), 
        .D(\u_inFIFO/n534 ), .Q(\u_inFIFO/n538 ) );
  INV3 U3556 ( .A(\u_outFIFO/n1118 ), .Q(n1804) );
  AOI221 U3557 ( .A(\u_outFIFO/N141 ), .B(\u_outFIFO/n1119 ), .C(
        \u_outFIFO/outReadCount[6] ), .D(\u_outFIFO/n1120 ), .Q(
        \u_outFIFO/n1118 ) );
  XOR21 U3558 ( .A(\u_outFIFO/add_260/carry [6]), .B(
        \u_outFIFO/outReadCount[6] ), .Q(\u_outFIFO/N141 ) );
  NAND22 U3559 ( .A(\u_decoder/fir_filter/I_data_mult_1_buff [2]), .B(n1159), 
        .Q(\u_decoder/fir_filter/n1120 ) );
  NAND22 U3560 ( .A(\u_decoder/fir_filter/I_data_mult_7_buff [2]), .B(n1155), 
        .Q(\u_decoder/fir_filter/n1022 ) );
  NAND22 U3561 ( .A(\u_decoder/fir_filter/Q_data_mult_1_buff [2]), .B(n1152), 
        .Q(\u_decoder/fir_filter/n823 ) );
  NAND22 U3562 ( .A(\u_decoder/fir_filter/Q_data_mult_7_buff [2]), .B(n1153), 
        .Q(\u_decoder/fir_filter/n725 ) );
  NAND31 U3563 ( .A(\u_coder/N1149 ), .B(\u_coder/n94 ), .C(\u_coder/n213 ), 
        .Q(\u_coder/n313 ) );
  NAND22 U3564 ( .A(\u_decoder/fir_filter/I_data_mult_0_buff [0]), .B(n1160), 
        .Q(\u_decoder/fir_filter/n1134 ) );
  NAND22 U3565 ( .A(\u_decoder/fir_filter/I_data_mult_1_buff [0]), .B(n1159), 
        .Q(\u_decoder/fir_filter/n1118 ) );
  NAND22 U3566 ( .A(\u_decoder/fir_filter/I_data_mult_2_buff [1]), .B(n1158), 
        .Q(\u_decoder/fir_filter/n1103 ) );
  NAND22 U3567 ( .A(\u_decoder/fir_filter/I_data_mult_3_buff [0]), .B(n1157), 
        .Q(\u_decoder/fir_filter/n1086 ) );
  NAND22 U3568 ( .A(\u_decoder/fir_filter/I_data_mult_5_buff [0]), .B(n1153), 
        .Q(\u_decoder/fir_filter/n1054 ) );
  NAND22 U3569 ( .A(\u_decoder/fir_filter/I_data_mult_6_buff [1]), .B(n1157), 
        .Q(\u_decoder/fir_filter/n1038 ) );
  NAND22 U3570 ( .A(\u_decoder/fir_filter/I_data_mult_7_buff [0]), .B(n1159), 
        .Q(\u_decoder/fir_filter/n1020 ) );
  NAND22 U3571 ( .A(\u_decoder/fir_filter/Q_data_mult_0_buff [0]), .B(n1152), 
        .Q(\u_decoder/fir_filter/n837 ) );
  NAND22 U3572 ( .A(\u_decoder/fir_filter/Q_data_mult_1_buff [0]), .B(n1151), 
        .Q(\u_decoder/fir_filter/n821 ) );
  NAND22 U3573 ( .A(\u_decoder/fir_filter/Q_data_mult_2_buff [1]), .B(n1155), 
        .Q(\u_decoder/fir_filter/n806 ) );
  NAND22 U3574 ( .A(\u_decoder/fir_filter/Q_data_mult_3_buff [0]), .B(n1153), 
        .Q(\u_decoder/fir_filter/n789 ) );
  NAND22 U3575 ( .A(\u_decoder/fir_filter/Q_data_mult_5_buff [0]), .B(n1155), 
        .Q(\u_decoder/fir_filter/n757 ) );
  NAND22 U3576 ( .A(\u_decoder/fir_filter/Q_data_mult_6_buff [1]), .B(n1153), 
        .Q(\u_decoder/fir_filter/n741 ) );
  NAND22 U3577 ( .A(\u_decoder/fir_filter/Q_data_mult_7_buff [0]), .B(n1153), 
        .Q(\u_decoder/fir_filter/n723 ) );
  BUF2 U3578 ( .A(\u_outFIFO/N39 ), .Q(n759) );
  INV3 U3579 ( .A(\u_outFIFO/n1111 ), .Q(n1793) );
  INV3 U3580 ( .A(\u_outFIFO/n1106 ), .Q(n1791) );
  INV3 U3581 ( .A(\u_outFIFO/n1099 ), .Q(n1788) );
  INV3 U3582 ( .A(\u_outFIFO/n1097 ), .Q(n1787) );
  INV3 U3583 ( .A(\u_outFIFO/n1091 ), .Q(n1784) );
  INV3 U3584 ( .A(\u_outFIFO/n1089 ), .Q(n1783) );
  INV3 U3585 ( .A(\u_outFIFO/n1080 ), .Q(n1779) );
  INV3 U3586 ( .A(\u_outFIFO/n1072 ), .Q(n1775) );
  INV3 U3587 ( .A(\u_outFIFO/n1064 ), .Q(n1771) );
  INV3 U3588 ( .A(\u_outFIFO/n1056 ), .Q(n1767) );
  INV3 U3589 ( .A(\u_outFIFO/n1049 ), .Q(n1764) );
  INV3 U3590 ( .A(\u_outFIFO/n1047 ), .Q(n1763) );
  INV3 U3591 ( .A(\u_outFIFO/n1045 ), .Q(n1762) );
  INV3 U3592 ( .A(\u_outFIFO/n1043 ), .Q(n1761) );
  INV3 U3593 ( .A(\u_outFIFO/n1041 ), .Q(n1760) );
  INV3 U3594 ( .A(\u_outFIFO/n1039 ), .Q(n1759) );
  INV3 U3595 ( .A(\u_outFIFO/n1037 ), .Q(n1758) );
  INV3 U3596 ( .A(\u_outFIFO/n1035 ), .Q(n1757) );
  INV3 U3597 ( .A(\u_outFIFO/n1033 ), .Q(n1756) );
  INV3 U3598 ( .A(\u_outFIFO/n1031 ), .Q(n1755) );
  INV3 U3599 ( .A(\u_outFIFO/n1029 ), .Q(n1754) );
  INV3 U3600 ( .A(\u_outFIFO/n1023 ), .Q(n1751) );
  INV3 U3601 ( .A(\u_outFIFO/n1021 ), .Q(n1750) );
  INV3 U3602 ( .A(\u_outFIFO/n1018 ), .Q(n1749) );
  INV3 U3603 ( .A(\u_outFIFO/n1016 ), .Q(n1748) );
  INV3 U3604 ( .A(\u_outFIFO/n1014 ), .Q(n1747) );
  INV3 U3605 ( .A(\u_outFIFO/n1009 ), .Q(n1745) );
  INV3 U3606 ( .A(\u_outFIFO/n1005 ), .Q(n1743) );
  INV3 U3607 ( .A(\u_outFIFO/n996 ), .Q(n1739) );
  INV3 U3608 ( .A(\u_outFIFO/n991 ), .Q(n1737) );
  INV3 U3609 ( .A(\u_outFIFO/n989 ), .Q(n1736) );
  INV3 U3610 ( .A(\u_outFIFO/n987 ), .Q(n1735) );
  INV3 U3611 ( .A(\u_outFIFO/n980 ), .Q(n1733) );
  INV3 U3612 ( .A(\u_outFIFO/n974 ), .Q(n1731) );
  INV3 U3613 ( .A(\u_outFIFO/n938 ), .Q(n1714) );
  INV3 U3614 ( .A(\u_outFIFO/n936 ), .Q(n1713) );
  INV3 U3615 ( .A(\u_outFIFO/n934 ), .Q(n1712) );
  INV3 U3616 ( .A(\u_outFIFO/n932 ), .Q(n1711) );
  INV3 U3617 ( .A(\u_outFIFO/n930 ), .Q(n1710) );
  INV3 U3618 ( .A(\u_outFIFO/n928 ), .Q(n1709) );
  INV3 U3619 ( .A(\u_outFIFO/n926 ), .Q(n1708) );
  INV3 U3620 ( .A(\u_outFIFO/n924 ), .Q(n1707) );
  INV3 U3621 ( .A(\u_outFIFO/n922 ), .Q(n1706) );
  INV3 U3622 ( .A(\u_outFIFO/n920 ), .Q(n1705) );
  INV3 U3623 ( .A(\u_outFIFO/n918 ), .Q(n1704) );
  INV3 U3624 ( .A(\u_outFIFO/n916 ), .Q(n1703) );
  INV3 U3625 ( .A(\u_outFIFO/n914 ), .Q(n1702) );
  INV3 U3626 ( .A(\u_outFIFO/n912 ), .Q(n1701) );
  INV3 U3627 ( .A(\u_outFIFO/n910 ), .Q(n1700) );
  INV3 U3628 ( .A(\u_outFIFO/n908 ), .Q(n1699) );
  INV3 U3629 ( .A(\u_outFIFO/n906 ), .Q(n1698) );
  INV3 U3630 ( .A(\u_outFIFO/n904 ), .Q(n1697) );
  INV3 U3631 ( .A(\u_outFIFO/n902 ), .Q(n1696) );
  INV3 U3632 ( .A(\u_outFIFO/n892 ), .Q(n1691) );
  INV3 U3633 ( .A(\u_outFIFO/n884 ), .Q(n1687) );
  INV3 U3634 ( .A(\u_outFIFO/n880 ), .Q(n1685) );
  INV3 U3635 ( .A(\u_outFIFO/n878 ), .Q(n1684) );
  INV3 U3636 ( .A(\u_outFIFO/n872 ), .Q(n1681) );
  INV3 U3637 ( .A(\u_outFIFO/n858 ), .Q(n1674) );
  INV3 U3638 ( .A(\u_outFIFO/n856 ), .Q(n1673) );
  INV3 U3639 ( .A(\u_outFIFO/n854 ), .Q(n1672) );
  INV3 U3640 ( .A(\u_outFIFO/n850 ), .Q(n1670) );
  INV3 U3641 ( .A(\u_outFIFO/n847 ), .Q(n1669) );
  INV3 U3642 ( .A(\u_outFIFO/n838 ), .Q(n1666) );
  INV3 U3643 ( .A(\u_outFIFO/n836 ), .Q(n1665) );
  INV3 U3644 ( .A(\u_outFIFO/n832 ), .Q(n1663) );
  INV3 U3645 ( .A(\u_outFIFO/n829 ), .Q(n1662) );
  INV3 U3646 ( .A(\u_outFIFO/n827 ), .Q(n1661) );
  INV3 U3647 ( .A(\u_outFIFO/n823 ), .Q(n1659) );
  INV3 U3648 ( .A(\u_outFIFO/n821 ), .Q(n1658) );
  INV3 U3649 ( .A(\u_outFIFO/n819 ), .Q(n1657) );
  INV3 U3650 ( .A(\u_outFIFO/n815 ), .Q(n1655) );
  INV3 U3651 ( .A(\u_outFIFO/n813 ), .Q(n1654) );
  INV3 U3652 ( .A(\u_outFIFO/n811 ), .Q(n1653) );
  INV3 U3653 ( .A(\u_outFIFO/n807 ), .Q(n1651) );
  INV3 U3654 ( .A(\u_outFIFO/n805 ), .Q(n1650) );
  INV3 U3655 ( .A(\u_outFIFO/n803 ), .Q(n1649) );
  INV3 U3656 ( .A(\u_outFIFO/n801 ), .Q(n1648) );
  INV3 U3657 ( .A(\u_outFIFO/n799 ), .Q(n1647) );
  INV3 U3658 ( .A(\u_outFIFO/n797 ), .Q(n1646) );
  INV3 U3659 ( .A(\u_outFIFO/n795 ), .Q(n1645) );
  INV3 U3660 ( .A(\u_outFIFO/n793 ), .Q(n1644) );
  INV3 U3661 ( .A(\u_outFIFO/n791 ), .Q(n1643) );
  INV3 U3662 ( .A(\u_outFIFO/n789 ), .Q(n1642) );
  INV3 U3663 ( .A(\u_outFIFO/n787 ), .Q(n1641) );
  INV3 U3664 ( .A(\u_outFIFO/n785 ), .Q(n1640) );
  INV3 U3665 ( .A(\u_outFIFO/n783 ), .Q(n1639) );
  INV3 U3666 ( .A(\u_outFIFO/n781 ), .Q(n1638) );
  INV3 U3667 ( .A(\u_outFIFO/n779 ), .Q(n1637) );
  INV3 U3668 ( .A(\u_outFIFO/n777 ), .Q(n1636) );
  INV3 U3669 ( .A(\u_outFIFO/n775 ), .Q(n1635) );
  INV3 U3670 ( .A(\u_outFIFO/n771 ), .Q(n1633) );
  INV3 U3671 ( .A(\u_outFIFO/n769 ), .Q(n1632) );
  INV3 U3672 ( .A(\u_outFIFO/n767 ), .Q(n1631) );
  INV3 U3673 ( .A(\u_outFIFO/n765 ), .Q(n1630) );
  INV3 U3674 ( .A(\u_outFIFO/n763 ), .Q(n1629) );
  INV3 U3675 ( .A(\u_outFIFO/n761 ), .Q(n1628) );
  INV3 U3676 ( .A(\u_outFIFO/n759 ), .Q(n1627) );
  INV3 U3677 ( .A(\u_outFIFO/n757 ), .Q(n1626) );
  INV3 U3678 ( .A(\u_outFIFO/n755 ), .Q(n1625) );
  INV3 U3679 ( .A(\u_outFIFO/n753 ), .Q(n1624) );
  INV3 U3680 ( .A(\u_outFIFO/n751 ), .Q(n1623) );
  INV3 U3681 ( .A(\u_outFIFO/n749 ), .Q(n1622) );
  INV3 U3682 ( .A(\u_outFIFO/n747 ), .Q(n1621) );
  INV3 U3683 ( .A(\u_outFIFO/n745 ), .Q(n1620) );
  INV3 U3684 ( .A(\u_outFIFO/n743 ), .Q(n1619) );
  INV3 U3685 ( .A(\u_outFIFO/n741 ), .Q(n1618) );
  INV3 U3686 ( .A(\u_outFIFO/n739 ), .Q(n1617) );
  INV3 U3687 ( .A(\u_outFIFO/n733 ), .Q(n1614) );
  INV3 U3688 ( .A(\u_outFIFO/n725 ), .Q(n1610) );
  INV3 U3689 ( .A(\u_outFIFO/n717 ), .Q(n1606) );
  INV3 U3690 ( .A(\u_outFIFO/n714 ), .Q(n1605) );
  INV3 U3691 ( .A(\u_outFIFO/n705 ), .Q(n1602) );
  INV3 U3692 ( .A(\u_outFIFO/n703 ), .Q(n1601) );
  INV3 U3693 ( .A(\u_outFIFO/n701 ), .Q(n1600) );
  INV3 U3694 ( .A(\u_outFIFO/n699 ), .Q(n1599) );
  INV3 U3695 ( .A(\u_outFIFO/n697 ), .Q(n1598) );
  INV3 U3696 ( .A(\u_outFIFO/n695 ), .Q(n1597) );
  INV3 U3697 ( .A(\u_outFIFO/n693 ), .Q(n1596) );
  INV3 U3698 ( .A(\u_outFIFO/n691 ), .Q(n1595) );
  INV3 U3699 ( .A(\u_outFIFO/n689 ), .Q(n1594) );
  INV3 U3700 ( .A(\u_outFIFO/n687 ), .Q(n1593) );
  INV3 U3701 ( .A(\u_outFIFO/n685 ), .Q(n1592) );
  INV3 U3702 ( .A(\u_outFIFO/n683 ), .Q(n1591) );
  NAND31 U3703 ( .A(\u_coder/N1143 ), .B(\u_coder/n91 ), .C(n2105), .Q(
        \u_coder/n306 ) );
  NAND22 U3704 ( .A(\u_decoder/fir_filter/I_data_mult_8_buff [14]), .B(n1158), 
        .Q(\u_decoder/fir_filter/n1011 ) );
  NAND22 U3705 ( .A(\u_decoder/fir_filter/I_data_mult_8_buff [13]), .B(n1154), 
        .Q(\u_decoder/fir_filter/n1010 ) );
  NAND22 U3706 ( .A(\u_decoder/fir_filter/I_data_mult_8_buff [12]), .B(n1156), 
        .Q(\u_decoder/fir_filter/n1009 ) );
  NAND22 U3707 ( .A(\u_decoder/fir_filter/Q_data_mult_8_buff [14]), .B(n1151), 
        .Q(\u_decoder/fir_filter/n713 ) );
  NAND22 U3708 ( .A(\u_decoder/fir_filter/Q_data_mult_8_buff [13]), .B(n1151), 
        .Q(\u_decoder/fir_filter/n712 ) );
  NAND22 U3709 ( .A(\u_decoder/fir_filter/Q_data_mult_8_buff [12]), .B(n1151), 
        .Q(\u_decoder/fir_filter/n711 ) );
  NAND22 U3710 ( .A(\u_decoder/fir_filter/I_data_mult_8_buff [11]), .B(n1153), 
        .Q(\u_decoder/fir_filter/n1008 ) );
  NAND22 U3711 ( .A(\u_decoder/fir_filter/I_data_mult_8_buff [10]), .B(n1152), 
        .Q(\u_decoder/fir_filter/n1007 ) );
  NAND22 U3712 ( .A(\u_decoder/fir_filter/I_data_mult_8_buff [9]), .B(n1152), 
        .Q(\u_decoder/fir_filter/n1006 ) );
  NAND22 U3713 ( .A(\u_decoder/fir_filter/I_data_mult_8_buff [8]), .B(n1151), 
        .Q(\u_decoder/fir_filter/n1005 ) );
  NAND22 U3714 ( .A(\u_decoder/fir_filter/I_data_mult_8_buff [7]), .B(n1160), 
        .Q(\u_decoder/fir_filter/n1004 ) );
  NAND22 U3715 ( .A(\u_decoder/fir_filter/I_data_mult_8_buff [6]), .B(n1158), 
        .Q(\u_decoder/fir_filter/n1003 ) );
  NAND22 U3716 ( .A(\u_decoder/fir_filter/I_data_mult_8_buff [5]), .B(n1150), 
        .Q(\u_decoder/fir_filter/n1002 ) );
  NAND22 U3717 ( .A(\u_decoder/fir_filter/I_data_mult_8_buff [4]), .B(n1150), 
        .Q(\u_decoder/fir_filter/n1001 ) );
  NAND22 U3718 ( .A(\u_decoder/fir_filter/I_data_mult_8_buff [3]), .B(n1150), 
        .Q(\u_decoder/fir_filter/n1000 ) );
  NAND22 U3719 ( .A(\u_decoder/fir_filter/I_data_mult_8_buff [2]), .B(n1150), 
        .Q(\u_decoder/fir_filter/n999 ) );
  NAND22 U3720 ( .A(\u_decoder/fir_filter/I_data_mult_8_buff [1]), .B(n1150), 
        .Q(\u_decoder/fir_filter/n998 ) );
  NAND22 U3721 ( .A(\u_decoder/fir_filter/I_data_mult_8_buff [0]), .B(n1150), 
        .Q(\u_decoder/fir_filter/n997 ) );
  NAND22 U3722 ( .A(\u_decoder/fir_filter/Q_data_mult_8_buff [11]), .B(n1151), 
        .Q(\u_decoder/fir_filter/n710 ) );
  NAND22 U3723 ( .A(\u_decoder/fir_filter/Q_data_mult_8_buff [10]), .B(n1151), 
        .Q(\u_decoder/fir_filter/n709 ) );
  NAND22 U3724 ( .A(\u_decoder/fir_filter/Q_data_mult_8_buff [9]), .B(n1151), 
        .Q(\u_decoder/fir_filter/n708 ) );
  NAND22 U3725 ( .A(\u_decoder/fir_filter/Q_data_mult_8_buff [8]), .B(n1151), 
        .Q(\u_decoder/fir_filter/n707 ) );
  NAND22 U3726 ( .A(\u_decoder/fir_filter/Q_data_mult_8_buff [7]), .B(n1151), 
        .Q(\u_decoder/fir_filter/n706 ) );
  NAND22 U3727 ( .A(\u_decoder/fir_filter/Q_data_mult_8_buff [6]), .B(n1151), 
        .Q(\u_decoder/fir_filter/n705 ) );
  NAND22 U3728 ( .A(\u_decoder/fir_filter/Q_data_mult_8_buff [5]), .B(n1151), 
        .Q(\u_decoder/fir_filter/n704 ) );
  NAND22 U3729 ( .A(\u_decoder/fir_filter/Q_data_mult_8_buff [4]), .B(n1150), 
        .Q(\u_decoder/fir_filter/n703 ) );
  NAND22 U3730 ( .A(\u_decoder/fir_filter/Q_data_mult_8_buff [3]), .B(n1150), 
        .Q(\u_decoder/fir_filter/n702 ) );
  NAND22 U3731 ( .A(\u_decoder/fir_filter/Q_data_mult_8_buff [2]), .B(n1150), 
        .Q(\u_decoder/fir_filter/n701 ) );
  NAND22 U3732 ( .A(\u_decoder/fir_filter/Q_data_mult_8_buff [1]), .B(n1150), 
        .Q(\u_decoder/fir_filter/n700 ) );
  NAND22 U3733 ( .A(\u_decoder/fir_filter/Q_data_mult_8_buff [0]), .B(n1150), 
        .Q(\u_decoder/fir_filter/n699 ) );
  NAND22 U3734 ( .A(\u_decoder/fir_filter/I_data_mult_2_buff [3]), .B(n1158), 
        .Q(\u_decoder/fir_filter/n1105 ) );
  NAND22 U3735 ( .A(\u_decoder/fir_filter/I_data_mult_6_buff [3]), .B(n1157), 
        .Q(\u_decoder/fir_filter/n1040 ) );
  NAND22 U3736 ( .A(\u_decoder/fir_filter/Q_data_mult_2_buff [3]), .B(n1160), 
        .Q(\u_decoder/fir_filter/n808 ) );
  NAND22 U3737 ( .A(\u_decoder/fir_filter/Q_data_mult_6_buff [3]), .B(n1155), 
        .Q(\u_decoder/fir_filter/n743 ) );
  NAND22 U3738 ( .A(\u_decoder/fir_filter/I_data_mult_1_buff [3]), .B(n1159), 
        .Q(\u_decoder/fir_filter/n1121 ) );
  NAND22 U3739 ( .A(\u_decoder/fir_filter/I_data_mult_7_buff [3]), .B(n1156), 
        .Q(\u_decoder/fir_filter/n1023 ) );
  NAND22 U3740 ( .A(\u_decoder/fir_filter/Q_data_mult_1_buff [3]), .B(n1152), 
        .Q(\u_decoder/fir_filter/n824 ) );
  NAND22 U3741 ( .A(\u_decoder/fir_filter/Q_data_mult_7_buff [3]), .B(n1153), 
        .Q(\u_decoder/fir_filter/n726 ) );
  NAND22 U3742 ( .A(\u_decoder/fir_filter/I_data_mult_3_buff [1]), .B(n1159), 
        .Q(\u_decoder/fir_filter/n1087 ) );
  NAND22 U3743 ( .A(\u_decoder/fir_filter/I_data_mult_5_buff [1]), .B(n1157), 
        .Q(\u_decoder/fir_filter/n1055 ) );
  NAND22 U3744 ( .A(\u_decoder/fir_filter/Q_data_mult_3_buff [1]), .B(n1153), 
        .Q(\u_decoder/fir_filter/n790 ) );
  NAND22 U3745 ( .A(\u_decoder/fir_filter/Q_data_mult_5_buff [1]), .B(n1155), 
        .Q(\u_decoder/fir_filter/n758 ) );
  NAND22 U3746 ( .A(\u_decoder/fir_filter/I_data_mult_0_buff [2]), .B(n1160), 
        .Q(\u_decoder/fir_filter/n1136 ) );
  NAND22 U3747 ( .A(\u_decoder/fir_filter/Q_data_mult_0_buff [2]), .B(n1161), 
        .Q(\u_decoder/fir_filter/n839 ) );
  NAND22 U3748 ( .A(\u_decoder/fir_filter/I_data_mult_1_buff [7]), .B(n1160), 
        .Q(\u_decoder/fir_filter/n1125 ) );
  NAND22 U3749 ( .A(\u_decoder/fir_filter/I_data_mult_7_buff [7]), .B(n1158), 
        .Q(\u_decoder/fir_filter/n1027 ) );
  NAND22 U3750 ( .A(\u_decoder/fir_filter/Q_data_mult_1_buff [7]), .B(n1152), 
        .Q(\u_decoder/fir_filter/n828 ) );
  NAND22 U3751 ( .A(\u_decoder/fir_filter/Q_data_mult_7_buff [7]), .B(n1154), 
        .Q(\u_decoder/fir_filter/n730 ) );
  NAND22 U3752 ( .A(\u_decoder/fir_filter/I_data_mult_0_buff [6]), .B(n1160), 
        .Q(\u_decoder/fir_filter/n1140 ) );
  NAND22 U3753 ( .A(\u_decoder/fir_filter/Q_data_mult_0_buff [6]), .B(n1151), 
        .Q(\u_decoder/fir_filter/n843 ) );
  NAND22 U3754 ( .A(\u_decoder/fir_filter/I_data_mult_1_buff [4]), .B(n1159), 
        .Q(\u_decoder/fir_filter/n1122 ) );
  NAND22 U3755 ( .A(\u_decoder/fir_filter/I_data_mult_2_buff [6]), .B(n1158), 
        .Q(\u_decoder/fir_filter/n1108 ) );
  NAND22 U3756 ( .A(\u_decoder/fir_filter/I_data_mult_2_buff [5]), .B(n1158), 
        .Q(\u_decoder/fir_filter/n1107 ) );
  NAND22 U3757 ( .A(\u_decoder/fir_filter/I_data_mult_2_buff [4]), .B(n1158), 
        .Q(\u_decoder/fir_filter/n1106 ) );
  NAND22 U3758 ( .A(\u_decoder/fir_filter/I_data_mult_3_buff [6]), .B(n1158), 
        .Q(\u_decoder/fir_filter/n1092 ) );
  NAND22 U3759 ( .A(\u_decoder/fir_filter/I_data_mult_3_buff [5]), .B(n1163), 
        .Q(\u_decoder/fir_filter/n1091 ) );
  NAND22 U3760 ( .A(\u_decoder/fir_filter/I_data_mult_3_buff [4]), .B(n1157), 
        .Q(\u_decoder/fir_filter/n1090 ) );
  NAND22 U3761 ( .A(\u_decoder/fir_filter/I_data_mult_3_buff [3]), .B(n1159), 
        .Q(\u_decoder/fir_filter/n1089 ) );
  NAND22 U3762 ( .A(\u_decoder/fir_filter/I_data_mult_3_buff [2]), .B(n1158), 
        .Q(\u_decoder/fir_filter/n1088 ) );
  NAND22 U3763 ( .A(\u_decoder/fir_filter/I_data_mult_5_buff [6]), .B(n1159), 
        .Q(\u_decoder/fir_filter/n1060 ) );
  NAND22 U3764 ( .A(\u_decoder/fir_filter/I_data_mult_5_buff [5]), .B(n1152), 
        .Q(\u_decoder/fir_filter/n1059 ) );
  NAND22 U3765 ( .A(\u_decoder/fir_filter/I_data_mult_5_buff [4]), .B(n1161), 
        .Q(\u_decoder/fir_filter/n1058 ) );
  NAND22 U3766 ( .A(\u_decoder/fir_filter/I_data_mult_5_buff [3]), .B(n1151), 
        .Q(\u_decoder/fir_filter/n1057 ) );
  NAND22 U3767 ( .A(\u_decoder/fir_filter/I_data_mult_5_buff [2]), .B(n1166), 
        .Q(\u_decoder/fir_filter/n1056 ) );
  NAND22 U3768 ( .A(\u_decoder/fir_filter/I_data_mult_6_buff [6]), .B(n1157), 
        .Q(\u_decoder/fir_filter/n1043 ) );
  NAND22 U3769 ( .A(\u_decoder/fir_filter/I_data_mult_6_buff [5]), .B(n1157), 
        .Q(\u_decoder/fir_filter/n1042 ) );
  NAND22 U3770 ( .A(\u_decoder/fir_filter/I_data_mult_6_buff [4]), .B(n1157), 
        .Q(\u_decoder/fir_filter/n1041 ) );
  NAND22 U3771 ( .A(\u_decoder/fir_filter/I_data_mult_7_buff [4]), .B(n1156), 
        .Q(\u_decoder/fir_filter/n1024 ) );
  NAND22 U3772 ( .A(\u_decoder/fir_filter/Q_data_mult_1_buff [4]), .B(n1152), 
        .Q(\u_decoder/fir_filter/n825 ) );
  NAND22 U3773 ( .A(\u_decoder/fir_filter/Q_data_mult_2_buff [6]), .B(n1157), 
        .Q(\u_decoder/fir_filter/n811 ) );
  NAND22 U3774 ( .A(\u_decoder/fir_filter/Q_data_mult_2_buff [5]), .B(n1164), 
        .Q(\u_decoder/fir_filter/n810 ) );
  NAND22 U3775 ( .A(\u_decoder/fir_filter/Q_data_mult_2_buff [4]), .B(n1165), 
        .Q(\u_decoder/fir_filter/n809 ) );
  NAND22 U3776 ( .A(\u_decoder/fir_filter/Q_data_mult_3_buff [6]), .B(n1154), 
        .Q(\u_decoder/fir_filter/n795 ) );
  NAND22 U3777 ( .A(\u_decoder/fir_filter/Q_data_mult_3_buff [5]), .B(n1153), 
        .Q(\u_decoder/fir_filter/n794 ) );
  NAND22 U3778 ( .A(\u_decoder/fir_filter/Q_data_mult_3_buff [4]), .B(n1153), 
        .Q(\u_decoder/fir_filter/n793 ) );
  NAND22 U3779 ( .A(\u_decoder/fir_filter/Q_data_mult_3_buff [3]), .B(n1153), 
        .Q(\u_decoder/fir_filter/n792 ) );
  NAND22 U3780 ( .A(\u_decoder/fir_filter/Q_data_mult_3_buff [2]), .B(n1153), 
        .Q(\u_decoder/fir_filter/n791 ) );
  NAND22 U3781 ( .A(\u_decoder/fir_filter/Q_data_mult_5_buff [6]), .B(n1155), 
        .Q(\u_decoder/fir_filter/n763 ) );
  NAND22 U3782 ( .A(\u_decoder/fir_filter/Q_data_mult_5_buff [5]), .B(n1155), 
        .Q(\u_decoder/fir_filter/n762 ) );
  NAND22 U3783 ( .A(\u_decoder/fir_filter/Q_data_mult_5_buff [4]), .B(n1155), 
        .Q(\u_decoder/fir_filter/n761 ) );
  NAND22 U3784 ( .A(\u_decoder/fir_filter/Q_data_mult_5_buff [3]), .B(n1155), 
        .Q(\u_decoder/fir_filter/n760 ) );
  NAND22 U3785 ( .A(\u_decoder/fir_filter/Q_data_mult_5_buff [2]), .B(n1155), 
        .Q(\u_decoder/fir_filter/n759 ) );
  NAND22 U3786 ( .A(\u_decoder/fir_filter/Q_data_mult_6_buff [6]), .B(n1154), 
        .Q(\u_decoder/fir_filter/n746 ) );
  NAND22 U3787 ( .A(\u_decoder/fir_filter/Q_data_mult_6_buff [5]), .B(n1156), 
        .Q(\u_decoder/fir_filter/n745 ) );
  NAND22 U3788 ( .A(\u_decoder/fir_filter/Q_data_mult_6_buff [4]), .B(n1154), 
        .Q(\u_decoder/fir_filter/n744 ) );
  NAND22 U3789 ( .A(\u_decoder/fir_filter/Q_data_mult_7_buff [4]), .B(n1153), 
        .Q(\u_decoder/fir_filter/n727 ) );
  NAND22 U3790 ( .A(\u_decoder/fir_filter/I_data_mult_0_buff [3]), .B(n1155), 
        .Q(\u_decoder/fir_filter/n1137 ) );
  NAND22 U3791 ( .A(\u_decoder/fir_filter/Q_data_mult_0_buff [3]), .B(n1153), 
        .Q(\u_decoder/fir_filter/n840 ) );
  IMUX40 U3792 ( .A(\u_inFIFO/N203 ), .B(\u_inFIFO/N201 ), .C(\u_inFIFO/N202 ), 
        .D(\u_inFIFO/N200 ), .S0(\u_inFIFO/N45 ), .S1(\u_inFIFO/N44 ), .Q(n379) );
  NOR21 U3793 ( .A(\u_outFIFO/n266 ), .B(\u_outFIFO/outReadCount[0] ), .Q(
        n2748) );
  INV3 U3794 ( .A(\u_cordic/mycordic/n404 ), .Q(n1873) );
  NAND22 U3795 ( .A(\u_cordic/mycordic/next_ANGLE_table[6][10] ), .B(n1215), 
        .Q(\u_cordic/mycordic/n404 ) );
  BUF2 U3796 ( .A(\u_outFIFO/N40 ), .Q(n760) );
  BUF2 U3797 ( .A(\u_inFIFO/N38 ), .Q(n764) );
  XOR21 U3798 ( .A(\u_cordic/mycordic/add_262/carry [9]), .B(
        \u_cordic/mycordic/present_ANGLE_table[6][9] ), .Q(
        \u_cordic/mycordic/N624 ) );
  XOR21 U3799 ( .A(\u_cordic/mycordic/add_262/carry [12]), .B(
        \u_cordic/mycordic/present_ANGLE_table[6][12] ), .Q(
        \u_cordic/mycordic/N627 ) );
  INV3 U3800 ( .A(\u_cordic/mycordic/n405 ), .Q(n1874) );
  NAND22 U3801 ( .A(\u_cordic/mycordic/next_ANGLE_table[6][9] ), .B(n1215), 
        .Q(\u_cordic/mycordic/n405 ) );
  INV3 U3802 ( .A(\u_cordic/mycordic/n403 ), .Q(n1872) );
  NAND22 U3803 ( .A(\u_cordic/mycordic/next_ANGLE_table[6][11] ), .B(n1215), 
        .Q(\u_cordic/mycordic/n403 ) );
  INV3 U3804 ( .A(\u_cordic/mycordic/n402 ), .Q(n1871) );
  NAND22 U3805 ( .A(\u_cordic/mycordic/next_ANGLE_table[6][12] ), .B(n1215), 
        .Q(\u_cordic/mycordic/n402 ) );
  NOR21 U3806 ( .A(\u_coder/i [6]), .B(\u_coder/i [5]), .Q(n2737) );
  INV3 U3807 ( .A(\u_outFIFO/n679 ), .Q(n1589) );
  INV3 U3808 ( .A(\u_outFIFO/n668 ), .Q(n1585) );
  INV3 U3809 ( .A(\u_outFIFO/n898 ), .Q(n1694) );
  INV3 U3810 ( .A(\u_outFIFO/n890 ), .Q(n1690) );
  INV3 U3811 ( .A(\u_outFIFO/n882 ), .Q(n1686) );
  INV3 U3812 ( .A(\u_outFIFO/n876 ), .Q(n1683) );
  INV3 U3813 ( .A(\u_outFIFO/n874 ), .Q(n1682) );
  INV3 U3814 ( .A(\u_outFIFO/n773 ), .Q(n1634) );
  INV3 U3815 ( .A(\u_outFIFO/n1076 ), .Q(n1777) );
  INV3 U3816 ( .A(\u_outFIFO/n1074 ), .Q(n1776) );
  INV3 U3817 ( .A(\u_outFIFO/n1070 ), .Q(n1774) );
  INV3 U3818 ( .A(\u_outFIFO/n1062 ), .Q(n1770) );
  INV3 U3819 ( .A(\u_outFIFO/n1054 ), .Q(n1766) );
  INV3 U3820 ( .A(\u_outFIFO/n1012 ), .Q(n1746) );
  INV3 U3821 ( .A(\u_outFIFO/n985 ), .Q(n1734) );
  INV3 U3822 ( .A(\u_outFIFO/n864 ), .Q(n1677) );
  INV3 U3823 ( .A(\u_outFIFO/n1103 ), .Q(n1790) );
  INV3 U3824 ( .A(\u_outFIFO/n1095 ), .Q(n1786) );
  INV3 U3825 ( .A(\u_outFIFO/n1087 ), .Q(n1782) );
  INV3 U3826 ( .A(\u_outFIFO/n1082 ), .Q(n1780) );
  INV3 U3827 ( .A(\u_outFIFO/n1003 ), .Q(n1742) );
  INV3 U3828 ( .A(\u_outFIFO/n866 ), .Q(n1678) );
  INV3 U3829 ( .A(\u_outFIFO/n969 ), .Q(n1729) );
  INV3 U3830 ( .A(\u_outFIFO/n965 ), .Q(n1727) );
  INV3 U3831 ( .A(\u_outFIFO/n962 ), .Q(n1726) );
  INV3 U3832 ( .A(\u_outFIFO/n960 ), .Q(n1725) );
  INV3 U3833 ( .A(\u_outFIFO/n956 ), .Q(n1723) );
  INV3 U3834 ( .A(\u_outFIFO/n954 ), .Q(n1722) );
  INV3 U3835 ( .A(\u_outFIFO/n952 ), .Q(n1721) );
  INV3 U3836 ( .A(\u_outFIFO/n948 ), .Q(n1719) );
  INV3 U3837 ( .A(\u_outFIFO/n946 ), .Q(n1718) );
  INV3 U3838 ( .A(\u_outFIFO/n994 ), .Q(n1738) );
  INV3 U3839 ( .A(\u_outFIFO/n862 ), .Q(n1676) );
  INV3 U3840 ( .A(\u_outFIFO/n860 ), .Q(n1675) );
  INV3 U3841 ( .A(\u_outFIFO/n729 ), .Q(n1612) );
  INV3 U3842 ( .A(\u_outFIFO/n727 ), .Q(n1611) );
  INV3 U3843 ( .A(\u_outFIFO/n1078 ), .Q(n1778) );
  INV3 U3844 ( .A(\u_outFIFO/n940 ), .Q(n1715) );
  INV3 U3845 ( .A(\u_outFIFO/n971 ), .Q(n1730) );
  INV3 U3846 ( .A(n2735), .Q(n2158) );
  NOR21 U3847 ( .A(\u_coder/i [18]), .B(\u_coder/i [17]), .Q(n2735) );
  INV3 U3848 ( .A(\u_inFIFO/n521 ), .Q(n1820) );
  AOI221 U3849 ( .A(n912), .B(\u_inFIFO/N43 ), .C(\u_inFIFO/n523 ), .D(
        \u_inFIFO/N131 ), .Q(\u_inFIFO/n521 ) );
  XOR21 U3850 ( .A(\u_inFIFO/add_253/carry [6]), .B(\u_inFIFO/N43 ), .Q(
        \u_inFIFO/N131 ) );
  INV3 U3851 ( .A(\u_cordic/mycordic/n406 ), .Q(n1875) );
  NAND22 U3852 ( .A(\u_cordic/mycordic/next_ANGLE_table[6][8] ), .B(n1215), 
        .Q(\u_cordic/mycordic/n406 ) );
  XNR21 U3853 ( .A(\u_cordic/mycordic/r173/carry [8]), .B(
        \u_cordic/mycordic/present_ANGLE_table[6][8] ), .Q(n380) );
  XNR21 U3854 ( .A(\u_cordic/mycordic/r173/carry [9]), .B(
        \u_cordic/mycordic/present_ANGLE_table[6][9] ), .Q(n381) );
  XNR21 U3855 ( .A(\u_cordic/mycordic/r173/carry [12]), .B(
        \u_cordic/mycordic/present_ANGLE_table[6][12] ), .Q(n382) );
  XNR21 U3856 ( .A(\u_outFIFO/add_360/carry [6]), .B(\u_outFIFO/N45 ), .Q(n383) );
  INV3 U3857 ( .A(\u_inFIFO/n518 ), .Q(n1960) );
  AOI221 U3858 ( .A(\u_inFIFO/N212 ), .B(\u_inFIFO/n513 ), .C(n1211), .D(
        \u_inFIFO/j_FIFO [1]), .Q(\u_inFIFO/n518 ) );
  INV3 U3859 ( .A(\u_inFIFO/n517 ), .Q(n1961) );
  AOI221 U3860 ( .A(\u_inFIFO/N213 ), .B(\u_inFIFO/n513 ), .C(n1211), .D(
        \u_inFIFO/j_FIFO [2]), .Q(\u_inFIFO/n517 ) );
  INV3 U3861 ( .A(\u_inFIFO/n516 ), .Q(n1962) );
  AOI221 U3862 ( .A(\u_inFIFO/N214 ), .B(\u_inFIFO/n513 ), .C(n1211), .D(
        \u_inFIFO/j_FIFO [3]), .Q(\u_inFIFO/n516 ) );
  INV3 U3863 ( .A(\u_inFIFO/n514 ), .Q(n1964) );
  AOI221 U3864 ( .A(\u_inFIFO/N216 ), .B(\u_inFIFO/n513 ), .C(n1211), .D(
        \u_inFIFO/j_FIFO [5]), .Q(\u_inFIFO/n514 ) );
  INV3 U3865 ( .A(\u_cordic/mycordic/n383 ), .Q(n1490) );
  AOI221 U3866 ( .A(n1905), .B(\u_cordic/mycordic/N291 ), .C(n773), .D(
        \u_cordic/mycordic/N259 ), .Q(\u_cordic/mycordic/n383 ) );
  INV3 U3867 ( .A(\u_decoder/fir_filter/n773 ), .Q(n2326) );
  AOI221 U3868 ( .A(\u_decoder/fir_filter/Q_data_mult_0 [0]), .B(n1084), .C(
        \u_decoder/fir_filter/Q_data_mult_4_buff [0]), .D(n1158), .Q(
        \u_decoder/fir_filter/n773 ) );
  INV3 U3869 ( .A(n2746), .Q(n2226) );
  AOI211 U3870 ( .A(n161), .B(n2748), .C(\u_outFIFO/outWriteCount[1] ), .Q(
        n2746) );
  INV3 U3871 ( .A(\u_decoder/fir_filter/n1072 ), .Q(n2300) );
  AOI221 U3872 ( .A(n4), .B(n1091), .C(
        \u_decoder/fir_filter/I_data_mult_4_buff [2]), .D(n1164), .Q(
        \u_decoder/fir_filter/n1072 ) );
  INV3 U3873 ( .A(\u_decoder/fir_filter/n775 ), .Q(n2371) );
  AOI221 U3874 ( .A(n3), .B(n1084), .C(
        \u_decoder/fir_filter/Q_data_mult_4_buff [2]), .D(n1157), .Q(
        \u_decoder/fir_filter/n775 ) );
  INV3 U3875 ( .A(\u_decoder/fir_filter/n1077 ), .Q(n2269) );
  AOI221 U3876 ( .A(\u_decoder/fir_filter/I_data_mult_4 [7]), .B(n1091), .C(
        \u_decoder/fir_filter/I_data_mult_4_buff [7]), .D(n1163), .Q(
        \u_decoder/fir_filter/n1077 ) );
  XOR21 U3877 ( .A(n1192), .B(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/SUMB[7][0] ), .Q(
        \u_decoder/fir_filter/I_data_mult_4 [7]) );
  INV3 U3878 ( .A(\u_decoder/fir_filter/n780 ), .Q(n2340) );
  AOI221 U3879 ( .A(\u_decoder/fir_filter/Q_data_mult_4 [7]), .B(n1083), .C(
        \u_decoder/fir_filter/Q_data_mult_4_buff [7]), .D(n1163), .Q(
        \u_decoder/fir_filter/n780 ) );
  XOR21 U3880 ( .A(n1194), .B(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/SUMB[7][0] ), .Q(
        \u_decoder/fir_filter/Q_data_mult_4 [7]) );
  INV3 U3881 ( .A(\u_cordic/mycordic/n511 ), .Q(n1461) );
  AOI221 U3882 ( .A(\u_cordic/mycordic/N340 ), .B(n772), .C(
        \u_cordic/mycordic/N372 ), .D(n1904), .Q(\u_cordic/mycordic/n511 ) );
  XNR21 U3883 ( .A(\u_cordic/mycordic/present_ANGLE_table[1][8] ), .B(
        \u_cordic/mycordic/sub_196/carry[8] ), .Q(\u_cordic/mycordic/N372 ) );
  XOR21 U3884 ( .A(\u_cordic/mycordic/present_ANGLE_table[1][8] ), .B(
        \u_cordic/mycordic/add_191/carry[8] ), .Q(\u_cordic/mycordic/N340 ) );
  INV3 U3885 ( .A(\u_cordic/mycordic/n510 ), .Q(n1462) );
  AOI221 U3886 ( .A(\u_cordic/mycordic/N341 ), .B(\u_cordic/mycordic/n336 ), 
        .C(\u_cordic/mycordic/N373 ), .D(n1904), .Q(\u_cordic/mycordic/n510 )
         );
  XNR21 U3887 ( .A(\u_cordic/mycordic/present_ANGLE_table[1][9] ), .B(
        \u_cordic/mycordic/sub_196/carry[9] ), .Q(\u_cordic/mycordic/N373 ) );
  XOR21 U3888 ( .A(\u_cordic/mycordic/present_ANGLE_table[1][9] ), .B(
        \u_cordic/mycordic/add_191/carry[9] ), .Q(\u_cordic/mycordic/N341 ) );
  INV3 U3889 ( .A(\u_cordic/mycordic/n509 ), .Q(n1463) );
  AOI221 U3890 ( .A(\u_cordic/mycordic/N342 ), .B(n772), .C(
        \u_cordic/mycordic/N374 ), .D(n1904), .Q(\u_cordic/mycordic/n509 ) );
  XNR21 U3891 ( .A(\u_cordic/mycordic/present_ANGLE_table[1][10] ), .B(
        \u_cordic/mycordic/sub_196/carry[10] ), .Q(\u_cordic/mycordic/N374 )
         );
  XOR21 U3892 ( .A(\u_cordic/mycordic/present_ANGLE_table[1][10] ), .B(
        \u_cordic/mycordic/add_191/carry[10] ), .Q(\u_cordic/mycordic/N342 )
         );
  INV3 U3893 ( .A(\u_cordic/mycordic/n494 ), .Q(n1555) );
  AOI221 U3894 ( .A(\u_cordic/mycordic/N405 ), .B(n778), .C(
        \u_cordic/mycordic/N437 ), .D(n1908), .Q(\u_cordic/mycordic/n494 ) );
  XNR21 U3895 ( .A(\u_cordic/mycordic/present_ANGLE_table[2][9] ), .B(
        \u_cordic/mycordic/sub_207/carry [9]), .Q(\u_cordic/mycordic/N437 ) );
  XOR21 U3896 ( .A(\u_cordic/mycordic/present_ANGLE_table[2][9] ), .B(
        \u_cordic/mycordic/add_202/carry [9]), .Q(\u_cordic/mycordic/N405 ) );
  INV3 U3897 ( .A(\u_cordic/mycordic/n493 ), .Q(n1556) );
  AOI221 U3898 ( .A(\u_cordic/mycordic/N406 ), .B(\u_cordic/mycordic/n332 ), 
        .C(\u_cordic/mycordic/N438 ), .D(n1908), .Q(\u_cordic/mycordic/n493 )
         );
  XNR21 U3899 ( .A(\u_cordic/mycordic/present_ANGLE_table[2][10] ), .B(
        \u_cordic/mycordic/sub_207/carry [10]), .Q(\u_cordic/mycordic/N438 )
         );
  XOR21 U3900 ( .A(\u_cordic/mycordic/present_ANGLE_table[2][10] ), .B(
        \u_cordic/mycordic/add_202/carry [10]), .Q(\u_cordic/mycordic/N406 )
         );
  INV3 U3901 ( .A(\u_cordic/mycordic/n492 ), .Q(n1557) );
  AOI221 U3902 ( .A(\u_cordic/mycordic/N407 ), .B(n778), .C(
        \u_cordic/mycordic/N439 ), .D(n1908), .Q(\u_cordic/mycordic/n492 ) );
  XNR21 U3903 ( .A(\u_cordic/mycordic/present_ANGLE_table[2][11] ), .B(
        \u_cordic/mycordic/sub_207/carry [11]), .Q(\u_cordic/mycordic/N439 )
         );
  XOR21 U3904 ( .A(\u_cordic/mycordic/present_ANGLE_table[2][11] ), .B(
        \u_cordic/mycordic/add_202/carry [11]), .Q(\u_cordic/mycordic/N407 )
         );
  INV3 U3905 ( .A(\u_cordic/mycordic/n491 ), .Q(n1558) );
  AOI221 U3906 ( .A(\u_cordic/mycordic/N408 ), .B(\u_cordic/mycordic/n332 ), 
        .C(\u_cordic/mycordic/N440 ), .D(n1908), .Q(\u_cordic/mycordic/n491 )
         );
  XNR21 U3907 ( .A(\u_cordic/mycordic/present_ANGLE_table[2][12] ), .B(
        \u_cordic/mycordic/sub_207/carry [12]), .Q(\u_cordic/mycordic/N440 )
         );
  XOR21 U3908 ( .A(\u_cordic/mycordic/present_ANGLE_table[2][12] ), .B(
        \u_cordic/mycordic/add_202/carry [12]), .Q(\u_cordic/mycordic/N408 )
         );
  INV3 U3909 ( .A(\u_cordic/mycordic/n463 ), .Q(n1505) );
  AOI221 U3910 ( .A(\u_cordic/mycordic/N509 ), .B(n776), .C(
        \u_cordic/mycordic/N526 ), .D(n1906), .Q(\u_cordic/mycordic/n463 ) );
  XNR21 U3911 ( .A(\u_cordic/mycordic/present_ANGLE_table[4][8] ), .B(
        \u_cordic/mycordic/sub_229/carry[8] ), .Q(\u_cordic/mycordic/N526 ) );
  XOR21 U3912 ( .A(\u_cordic/mycordic/present_ANGLE_table[4][8] ), .B(
        \u_cordic/mycordic/add_224/carry[8] ), .Q(\u_cordic/mycordic/N509 ) );
  INV3 U3913 ( .A(\u_cordic/mycordic/n462 ), .Q(n1506) );
  AOI221 U3914 ( .A(\u_cordic/mycordic/N510 ), .B(\u_cordic/mycordic/n456 ), 
        .C(\u_cordic/mycordic/N527 ), .D(n1906), .Q(\u_cordic/mycordic/n462 )
         );
  XNR21 U3915 ( .A(\u_cordic/mycordic/present_ANGLE_table[4][9] ), .B(
        \u_cordic/mycordic/sub_229/carry[9] ), .Q(\u_cordic/mycordic/N527 ) );
  XOR21 U3916 ( .A(\u_cordic/mycordic/present_ANGLE_table[4][9] ), .B(
        \u_cordic/mycordic/add_224/carry[9] ), .Q(\u_cordic/mycordic/N510 ) );
  INV3 U3917 ( .A(\u_cordic/mycordic/n461 ), .Q(n1507) );
  AOI221 U3918 ( .A(\u_cordic/mycordic/N511 ), .B(n776), .C(
        \u_cordic/mycordic/N528 ), .D(n1906), .Q(\u_cordic/mycordic/n461 ) );
  XNR21 U3919 ( .A(\u_cordic/mycordic/present_ANGLE_table[4][10] ), .B(
        \u_cordic/mycordic/sub_229/carry[10] ), .Q(\u_cordic/mycordic/N528 )
         );
  XOR21 U3920 ( .A(\u_cordic/mycordic/present_ANGLE_table[4][10] ), .B(
        \u_cordic/mycordic/add_224/carry[10] ), .Q(\u_cordic/mycordic/N511 )
         );
  INV3 U3921 ( .A(\u_cordic/mycordic/n460 ), .Q(n1508) );
  AOI221 U3922 ( .A(\u_cordic/mycordic/N512 ), .B(n776), .C(
        \u_cordic/mycordic/N529 ), .D(n1906), .Q(\u_cordic/mycordic/n460 ) );
  XNR21 U3923 ( .A(\u_cordic/mycordic/present_ANGLE_table[4][11] ), .B(
        \u_cordic/mycordic/sub_229/carry[11] ), .Q(\u_cordic/mycordic/N529 )
         );
  XOR21 U3924 ( .A(\u_cordic/mycordic/present_ANGLE_table[4][11] ), .B(
        \u_cordic/mycordic/add_224/carry[11] ), .Q(\u_cordic/mycordic/N512 )
         );
  INV3 U3925 ( .A(\u_cordic/mycordic/n442 ), .Q(n1448) );
  AOI221 U3926 ( .A(\u_cordic/mycordic/N545 ), .B(n771), .C(
        \u_cordic/mycordic/N561 ), .D(n1903), .Q(\u_cordic/mycordic/n442 ) );
  XNR21 U3927 ( .A(\u_cordic/mycordic/present_ANGLE_table[5][11] ), .B(
        \u_cordic/mycordic/sub_236/carry [11]), .Q(\u_cordic/mycordic/N561 )
         );
  XOR21 U3928 ( .A(\u_cordic/mycordic/present_ANGLE_table[5][11] ), .B(
        \u_cordic/mycordic/add_233/carry [11]), .Q(\u_cordic/mycordic/N545 )
         );
  INV3 U3929 ( .A(\u_decoder/fir_filter/n1075 ), .Q(n2271) );
  AOI221 U3930 ( .A(\u_decoder/fir_filter/I_data_mult_4 [5]), .B(n1091), .C(
        \u_decoder/fir_filter/I_data_mult_4_buff [5]), .D(n1164), .Q(
        \u_decoder/fir_filter/n1075 ) );
  INV3 U3931 ( .A(\u_decoder/fir_filter/n1074 ), .Q(n2272) );
  AOI221 U3932 ( .A(\u_decoder/fir_filter/I_data_mult_4 [4]), .B(n1091), .C(
        \u_decoder/fir_filter/I_data_mult_4_buff [4]), .D(n1164), .Q(
        \u_decoder/fir_filter/n1074 ) );
  INV3 U3933 ( .A(\u_decoder/fir_filter/n995 ), .Q(n2635) );
  AOI221 U3934 ( .A(\u_decoder/fir_filter/I_data_add_7 [1]), .B(n1091), .C(
        \u_decoder/fir_filter/I_data_add_7_buff [1]), .D(n1164), .Q(
        \u_decoder/fir_filter/n995 ) );
  INV3 U3935 ( .A(\u_decoder/fir_filter/n994 ), .Q(n2634) );
  AOI221 U3936 ( .A(\u_decoder/fir_filter/I_data_add_7 [2]), .B(n1091), .C(
        \u_decoder/fir_filter/I_data_add_7_buff [2]), .D(n1164), .Q(
        \u_decoder/fir_filter/n994 ) );
  INV3 U3937 ( .A(\u_decoder/fir_filter/n993 ), .Q(n2633) );
  AOI221 U3938 ( .A(\u_decoder/fir_filter/I_data_add_7 [3]), .B(n1091), .C(
        \u_decoder/fir_filter/I_data_add_7_buff [3]), .D(n1164), .Q(
        \u_decoder/fir_filter/n993 ) );
  INV3 U3939 ( .A(\u_decoder/fir_filter/n992 ), .Q(n2632) );
  AOI221 U3940 ( .A(\u_decoder/fir_filter/I_data_add_7 [4]), .B(n1091), .C(
        \u_decoder/fir_filter/I_data_add_7_buff [4]), .D(n1164), .Q(
        \u_decoder/fir_filter/n992 ) );
  INV3 U3941 ( .A(\u_decoder/fir_filter/n991 ), .Q(n2631) );
  AOI221 U3942 ( .A(\u_decoder/fir_filter/I_data_add_7 [5]), .B(n1091), .C(
        \u_decoder/fir_filter/I_data_add_7_buff [5]), .D(n1164), .Q(
        \u_decoder/fir_filter/n991 ) );
  INV3 U3943 ( .A(\u_decoder/fir_filter/n990 ), .Q(n2630) );
  AOI221 U3944 ( .A(\u_decoder/fir_filter/I_data_add_7 [6]), .B(n1091), .C(
        \u_decoder/fir_filter/I_data_add_7_buff [6]), .D(n1164), .Q(
        \u_decoder/fir_filter/n990 ) );
  INV3 U3945 ( .A(\u_decoder/fir_filter/n974 ), .Q(n2620) );
  AOI221 U3946 ( .A(\u_decoder/fir_filter/I_data_add_6 [1]), .B(n1092), .C(
        \u_decoder/fir_filter/I_data_add_6_buff [1]), .D(n1165), .Q(
        \u_decoder/fir_filter/n974 ) );
  INV3 U3947 ( .A(\u_decoder/fir_filter/n973 ), .Q(n2619) );
  AOI221 U3948 ( .A(\u_decoder/fir_filter/I_data_add_6 [2]), .B(n1092), .C(
        \u_decoder/fir_filter/I_data_add_6_buff [2]), .D(n1165), .Q(
        \u_decoder/fir_filter/n973 ) );
  INV3 U3949 ( .A(\u_decoder/fir_filter/n972 ), .Q(n2618) );
  AOI221 U3950 ( .A(\u_decoder/fir_filter/I_data_add_6 [3]), .B(n1092), .C(
        \u_decoder/fir_filter/I_data_add_6_buff [3]), .D(n1165), .Q(
        \u_decoder/fir_filter/n972 ) );
  INV3 U3951 ( .A(\u_decoder/fir_filter/n971 ), .Q(n2617) );
  AOI221 U3952 ( .A(\u_decoder/fir_filter/I_data_add_6 [4]), .B(n1092), .C(
        \u_decoder/fir_filter/I_data_add_6_buff [4]), .D(n1165), .Q(
        \u_decoder/fir_filter/n971 ) );
  INV3 U3953 ( .A(\u_decoder/fir_filter/n970 ), .Q(n2616) );
  AOI221 U3954 ( .A(\u_decoder/fir_filter/I_data_add_6 [5]), .B(n1092), .C(
        \u_decoder/fir_filter/I_data_add_6_buff [5]), .D(n1165), .Q(
        \u_decoder/fir_filter/n970 ) );
  INV3 U3955 ( .A(\u_decoder/fir_filter/n969 ), .Q(n2615) );
  AOI221 U3956 ( .A(\u_decoder/fir_filter/I_data_add_6 [6]), .B(n1092), .C(
        \u_decoder/fir_filter/I_data_add_6_buff [6]), .D(n1165), .Q(
        \u_decoder/fir_filter/n969 ) );
  INV3 U3957 ( .A(\u_decoder/fir_filter/n953 ), .Q(n2605) );
  AOI221 U3958 ( .A(\u_decoder/fir_filter/I_data_add_5 [1]), .B(n1093), .C(
        \u_decoder/fir_filter/I_data_add_5_buff [1]), .D(n1166), .Q(
        \u_decoder/fir_filter/n953 ) );
  INV3 U3959 ( .A(\u_decoder/fir_filter/n952 ), .Q(n2604) );
  AOI221 U3960 ( .A(\u_decoder/fir_filter/I_data_add_5 [2]), .B(n1093), .C(
        \u_decoder/fir_filter/I_data_add_5_buff [2]), .D(n1166), .Q(
        \u_decoder/fir_filter/n952 ) );
  INV3 U3961 ( .A(\u_decoder/fir_filter/n951 ), .Q(n2603) );
  AOI221 U3962 ( .A(\u_decoder/fir_filter/I_data_add_5 [3]), .B(n1093), .C(
        \u_decoder/fir_filter/I_data_add_5_buff [3]), .D(n1166), .Q(
        \u_decoder/fir_filter/n951 ) );
  INV3 U3963 ( .A(\u_decoder/fir_filter/n950 ), .Q(n2602) );
  AOI221 U3964 ( .A(\u_decoder/fir_filter/I_data_add_5 [4]), .B(n1093), .C(
        \u_decoder/fir_filter/I_data_add_5_buff [4]), .D(n1166), .Q(
        \u_decoder/fir_filter/n950 ) );
  INV3 U3965 ( .A(\u_decoder/fir_filter/n949 ), .Q(n2601) );
  AOI221 U3966 ( .A(\u_decoder/fir_filter/I_data_add_5 [5]), .B(n1093), .C(
        \u_decoder/fir_filter/I_data_add_5_buff [5]), .D(n1166), .Q(
        \u_decoder/fir_filter/n949 ) );
  INV3 U3967 ( .A(\u_decoder/fir_filter/n948 ), .Q(n2600) );
  AOI221 U3968 ( .A(\u_decoder/fir_filter/I_data_add_5 [6]), .B(n1093), .C(
        \u_decoder/fir_filter/I_data_add_5_buff [6]), .D(n1166), .Q(
        \u_decoder/fir_filter/n948 ) );
  INV3 U3969 ( .A(\u_decoder/fir_filter/n911 ), .Q(n2575) );
  AOI221 U3970 ( .A(\u_decoder/fir_filter/I_data_add_3 [1]), .B(n1095), .C(
        \u_decoder/fir_filter/I_data_add_3_buff [1]), .D(n1161), .Q(
        \u_decoder/fir_filter/n911 ) );
  INV3 U3971 ( .A(\u_decoder/fir_filter/n910 ), .Q(n2574) );
  AOI221 U3972 ( .A(\u_decoder/fir_filter/I_data_add_3 [2]), .B(n1095), .C(
        \u_decoder/fir_filter/I_data_add_3_buff [2]), .D(n1164), .Q(
        \u_decoder/fir_filter/n910 ) );
  INV3 U3973 ( .A(\u_decoder/fir_filter/n909 ), .Q(n2573) );
  AOI221 U3974 ( .A(\u_decoder/fir_filter/I_data_add_3 [3]), .B(n1095), .C(
        \u_decoder/fir_filter/I_data_add_3_buff [3]), .D(n1165), .Q(
        \u_decoder/fir_filter/n909 ) );
  INV3 U3975 ( .A(\u_decoder/fir_filter/n908 ), .Q(n2572) );
  AOI221 U3976 ( .A(\u_decoder/fir_filter/I_data_add_3 [4]), .B(n1095), .C(
        \u_decoder/fir_filter/I_data_add_3_buff [4]), .D(n1157), .Q(
        \u_decoder/fir_filter/n908 ) );
  INV3 U3977 ( .A(\u_decoder/fir_filter/n907 ), .Q(n2571) );
  AOI221 U3978 ( .A(\u_decoder/fir_filter/I_data_add_3 [5]), .B(n1095), .C(
        \u_decoder/fir_filter/I_data_add_3_buff [5]), .D(n1164), .Q(
        \u_decoder/fir_filter/n907 ) );
  INV3 U3979 ( .A(\u_decoder/fir_filter/n906 ), .Q(n2570) );
  AOI221 U3980 ( .A(\u_decoder/fir_filter/I_data_add_3 [6]), .B(n1095), .C(
        \u_decoder/fir_filter/I_data_add_3_buff [6]), .D(n1165), .Q(
        \u_decoder/fir_filter/n906 ) );
  INV3 U3981 ( .A(\u_decoder/fir_filter/n890 ), .Q(n2560) );
  AOI221 U3982 ( .A(\u_decoder/fir_filter/I_data_add_2 [1]), .B(n1096), .C(
        \u_decoder/fir_filter/I_data_add_2_buff [1]), .D(n1166), .Q(
        \u_decoder/fir_filter/n890 ) );
  INV3 U3983 ( .A(\u_decoder/fir_filter/n889 ), .Q(n2559) );
  AOI221 U3984 ( .A(\u_decoder/fir_filter/I_data_add_2 [2]), .B(n1096), .C(
        \u_decoder/fir_filter/I_data_add_2_buff [2]), .D(n1165), .Q(
        \u_decoder/fir_filter/n889 ) );
  INV3 U3985 ( .A(\u_decoder/fir_filter/n888 ), .Q(n2558) );
  AOI221 U3986 ( .A(\u_decoder/fir_filter/I_data_add_2 [3]), .B(n1096), .C(
        \u_decoder/fir_filter/I_data_add_2_buff [3]), .D(n1163), .Q(
        \u_decoder/fir_filter/n888 ) );
  INV3 U3987 ( .A(\u_decoder/fir_filter/n887 ), .Q(n2557) );
  AOI221 U3988 ( .A(\u_decoder/fir_filter/I_data_add_2 [4]), .B(n1096), .C(
        \u_decoder/fir_filter/I_data_add_2_buff [4]), .D(n1154), .Q(
        \u_decoder/fir_filter/n887 ) );
  INV3 U3989 ( .A(\u_decoder/fir_filter/n886 ), .Q(n2556) );
  AOI221 U3990 ( .A(\u_decoder/fir_filter/I_data_add_2 [5]), .B(n1096), .C(
        \u_decoder/fir_filter/I_data_add_2_buff [5]), .D(n1162), .Q(
        \u_decoder/fir_filter/n886 ) );
  INV3 U3991 ( .A(\u_decoder/fir_filter/n885 ), .Q(n2555) );
  AOI221 U3992 ( .A(\u_decoder/fir_filter/I_data_add_2 [6]), .B(n1096), .C(
        \u_decoder/fir_filter/I_data_add_2_buff [6]), .D(n1161), .Q(
        \u_decoder/fir_filter/n885 ) );
  INV3 U3993 ( .A(\u_decoder/fir_filter/n869 ), .Q(n2545) );
  AOI221 U3994 ( .A(\u_decoder/fir_filter/I_data_add_1 [1]), .B(n1097), .C(
        \u_decoder/fir_filter/I_data_add_1_buff [1]), .D(n1155), .Q(
        \u_decoder/fir_filter/n869 ) );
  INV3 U3995 ( .A(\u_decoder/fir_filter/n868 ), .Q(n2543) );
  AOI221 U3996 ( .A(\u_decoder/fir_filter/I_data_add_1 [2]), .B(n1097), .C(
        \u_decoder/fir_filter/I_data_add_1_buff [2]), .D(n1154), .Q(
        \u_decoder/fir_filter/n868 ) );
  INV3 U3997 ( .A(\u_decoder/fir_filter/n867 ), .Q(n2541) );
  AOI221 U3998 ( .A(\u_decoder/fir_filter/I_data_add_1 [3]), .B(n1097), .C(
        \u_decoder/fir_filter/I_data_add_1_buff [3]), .D(n1155), .Q(
        \u_decoder/fir_filter/n867 ) );
  INV3 U3999 ( .A(\u_decoder/fir_filter/n866 ), .Q(n2539) );
  AOI221 U4000 ( .A(\u_decoder/fir_filter/I_data_add_1 [4]), .B(n1097), .C(
        \u_decoder/fir_filter/I_data_add_1_buff [4]), .D(n1153), .Q(
        \u_decoder/fir_filter/n866 ) );
  INV3 U4001 ( .A(\u_decoder/fir_filter/n865 ), .Q(n2537) );
  AOI221 U4002 ( .A(\u_decoder/fir_filter/I_data_add_1 [5]), .B(n1097), .C(
        \u_decoder/fir_filter/I_data_add_1_buff [5]), .D(n1152), .Q(
        \u_decoder/fir_filter/n865 ) );
  INV3 U4003 ( .A(\u_decoder/fir_filter/n864 ), .Q(n2535) );
  AOI221 U4004 ( .A(\u_decoder/fir_filter/I_data_add_1 [6]), .B(n1097), .C(
        \u_decoder/fir_filter/I_data_add_1_buff [6]), .D(n1152), .Q(
        \u_decoder/fir_filter/n864 ) );
  INV3 U4005 ( .A(\u_decoder/fir_filter/n778 ), .Q(n2342) );
  AOI221 U4006 ( .A(\u_decoder/fir_filter/Q_data_mult_4 [5]), .B(n1084), .C(
        \u_decoder/fir_filter/Q_data_mult_4_buff [5]), .D(n1158), .Q(
        \u_decoder/fir_filter/n778 ) );
  INV3 U4007 ( .A(\u_decoder/fir_filter/n777 ), .Q(n2343) );
  AOI221 U4008 ( .A(\u_decoder/fir_filter/Q_data_mult_4 [4]), .B(n1084), .C(
        \u_decoder/fir_filter/Q_data_mult_4_buff [4]), .D(n1159), .Q(
        \u_decoder/fir_filter/n777 ) );
  INV3 U4009 ( .A(\u_decoder/fir_filter/n697 ), .Q(n2515) );
  AOI221 U4010 ( .A(\u_decoder/fir_filter/Q_data_add_7 [1]), .B(n1084), .C(
        \u_decoder/fir_filter/Q_data_add_7_buff [1]), .D(n1163), .Q(
        \u_decoder/fir_filter/n697 ) );
  INV3 U4011 ( .A(\u_decoder/fir_filter/n696 ), .Q(n2514) );
  AOI221 U4012 ( .A(\u_decoder/fir_filter/Q_data_add_7 [2]), .B(n1084), .C(
        \u_decoder/fir_filter/Q_data_add_7_buff [2]), .D(n1163), .Q(
        \u_decoder/fir_filter/n696 ) );
  INV3 U4013 ( .A(\u_decoder/fir_filter/n695 ), .Q(n2513) );
  AOI221 U4014 ( .A(\u_decoder/fir_filter/Q_data_add_7 [3]), .B(n1084), .C(
        \u_decoder/fir_filter/Q_data_add_7_buff [3]), .D(n1163), .Q(
        \u_decoder/fir_filter/n695 ) );
  INV3 U4015 ( .A(\u_decoder/fir_filter/n694 ), .Q(n2512) );
  AOI221 U4016 ( .A(\u_decoder/fir_filter/Q_data_add_7 [4]), .B(n1084), .C(
        \u_decoder/fir_filter/Q_data_add_7_buff [4]), .D(n1163), .Q(
        \u_decoder/fir_filter/n694 ) );
  INV3 U4017 ( .A(\u_decoder/fir_filter/n693 ), .Q(n2511) );
  AOI221 U4018 ( .A(\u_decoder/fir_filter/Q_data_add_7 [5]), .B(n1084), .C(
        \u_decoder/fir_filter/Q_data_add_7_buff [5]), .D(n1163), .Q(
        \u_decoder/fir_filter/n693 ) );
  INV3 U4019 ( .A(\u_decoder/fir_filter/n692 ), .Q(n2510) );
  AOI221 U4020 ( .A(\u_decoder/fir_filter/Q_data_add_7 [6]), .B(n1084), .C(
        \u_decoder/fir_filter/Q_data_add_7_buff [6]), .D(n1163), .Q(
        \u_decoder/fir_filter/n692 ) );
  INV3 U4021 ( .A(\u_decoder/fir_filter/n676 ), .Q(n2500) );
  AOI221 U4022 ( .A(\u_decoder/fir_filter/Q_data_add_6 [1]), .B(n1085), .C(
        \u_decoder/fir_filter/Q_data_add_6_buff [1]), .D(n1157), .Q(
        \u_decoder/fir_filter/n676 ) );
  INV3 U4023 ( .A(\u_decoder/fir_filter/n675 ), .Q(n2499) );
  AOI221 U4024 ( .A(\u_decoder/fir_filter/Q_data_add_6 [2]), .B(n1085), .C(
        \u_decoder/fir_filter/Q_data_add_6_buff [2]), .D(n1159), .Q(
        \u_decoder/fir_filter/n675 ) );
  INV3 U4025 ( .A(\u_decoder/fir_filter/n674 ), .Q(n2498) );
  AOI221 U4026 ( .A(\u_decoder/fir_filter/Q_data_add_6 [3]), .B(n1085), .C(
        \u_decoder/fir_filter/Q_data_add_6_buff [3]), .D(n1157), .Q(
        \u_decoder/fir_filter/n674 ) );
  INV3 U4027 ( .A(\u_decoder/fir_filter/n673 ), .Q(n2497) );
  AOI221 U4028 ( .A(\u_decoder/fir_filter/Q_data_add_6 [4]), .B(n1085), .C(
        \u_decoder/fir_filter/Q_data_add_6_buff [4]), .D(n1158), .Q(
        \u_decoder/fir_filter/n673 ) );
  INV3 U4029 ( .A(\u_decoder/fir_filter/n672 ), .Q(n2496) );
  AOI221 U4030 ( .A(\u_decoder/fir_filter/Q_data_add_6 [5]), .B(n1085), .C(
        \u_decoder/fir_filter/Q_data_add_6_buff [5]), .D(n1152), .Q(
        \u_decoder/fir_filter/n672 ) );
  INV3 U4031 ( .A(\u_decoder/fir_filter/n671 ), .Q(n2495) );
  AOI221 U4032 ( .A(\u_decoder/fir_filter/Q_data_add_6 [6]), .B(n1085), .C(
        \u_decoder/fir_filter/Q_data_add_6_buff [6]), .D(n1151), .Q(
        \u_decoder/fir_filter/n671 ) );
  INV3 U4033 ( .A(\u_decoder/fir_filter/n655 ), .Q(n2485) );
  AOI221 U4034 ( .A(\u_decoder/fir_filter/Q_data_add_5 [1]), .B(n1086), .C(
        \u_decoder/fir_filter/Q_data_add_5_buff [1]), .D(n1164), .Q(
        \u_decoder/fir_filter/n655 ) );
  INV3 U4035 ( .A(\u_decoder/fir_filter/n654 ), .Q(n2484) );
  AOI221 U4036 ( .A(\u_decoder/fir_filter/Q_data_add_5 [2]), .B(n1086), .C(
        \u_decoder/fir_filter/Q_data_add_5_buff [2]), .D(n1165), .Q(
        \u_decoder/fir_filter/n654 ) );
  INV3 U4037 ( .A(\u_decoder/fir_filter/n653 ), .Q(n2483) );
  AOI221 U4038 ( .A(\u_decoder/fir_filter/Q_data_add_5 [3]), .B(n1086), .C(
        \u_decoder/fir_filter/Q_data_add_5_buff [3]), .D(n1166), .Q(
        \u_decoder/fir_filter/n653 ) );
  INV3 U4039 ( .A(\u_decoder/fir_filter/n652 ), .Q(n2482) );
  AOI221 U4040 ( .A(\u_decoder/fir_filter/Q_data_add_5 [4]), .B(n1086), .C(
        \u_decoder/fir_filter/Q_data_add_5_buff [4]), .D(n1164), .Q(
        \u_decoder/fir_filter/n652 ) );
  INV3 U4041 ( .A(\u_decoder/fir_filter/n651 ), .Q(n2481) );
  AOI221 U4042 ( .A(\u_decoder/fir_filter/Q_data_add_5 [5]), .B(n1086), .C(
        \u_decoder/fir_filter/Q_data_add_5_buff [5]), .D(n1163), .Q(
        \u_decoder/fir_filter/n651 ) );
  INV3 U4043 ( .A(\u_decoder/fir_filter/n650 ), .Q(n2480) );
  AOI221 U4044 ( .A(\u_decoder/fir_filter/Q_data_add_5 [6]), .B(n1086), .C(
        \u_decoder/fir_filter/Q_data_add_5_buff [6]), .D(n1162), .Q(
        \u_decoder/fir_filter/n650 ) );
  INV3 U4045 ( .A(\u_decoder/fir_filter/n613 ), .Q(n2455) );
  AOI221 U4046 ( .A(\u_decoder/fir_filter/Q_data_add_3 [1]), .B(n1088), .C(
        \u_decoder/fir_filter/Q_data_add_3_buff [1]), .D(n1162), .Q(
        \u_decoder/fir_filter/n613 ) );
  INV3 U4047 ( .A(\u_decoder/fir_filter/n612 ), .Q(n2454) );
  AOI221 U4048 ( .A(\u_decoder/fir_filter/Q_data_add_3 [2]), .B(n1088), .C(
        \u_decoder/fir_filter/Q_data_add_3_buff [2]), .D(n1162), .Q(
        \u_decoder/fir_filter/n612 ) );
  INV3 U4049 ( .A(\u_decoder/fir_filter/n611 ), .Q(n2453) );
  AOI221 U4050 ( .A(\u_decoder/fir_filter/Q_data_add_3 [3]), .B(n1088), .C(
        \u_decoder/fir_filter/Q_data_add_3_buff [3]), .D(n1162), .Q(
        \u_decoder/fir_filter/n611 ) );
  INV3 U4051 ( .A(\u_decoder/fir_filter/n610 ), .Q(n2452) );
  AOI221 U4052 ( .A(\u_decoder/fir_filter/Q_data_add_3 [4]), .B(n1088), .C(
        \u_decoder/fir_filter/Q_data_add_3_buff [4]), .D(n1162), .Q(
        \u_decoder/fir_filter/n610 ) );
  INV3 U4053 ( .A(\u_decoder/fir_filter/n609 ), .Q(n2451) );
  AOI221 U4054 ( .A(\u_decoder/fir_filter/Q_data_add_3 [5]), .B(n1088), .C(
        \u_decoder/fir_filter/Q_data_add_3_buff [5]), .D(n1162), .Q(
        \u_decoder/fir_filter/n609 ) );
  INV3 U4055 ( .A(\u_decoder/fir_filter/n608 ), .Q(n2450) );
  AOI221 U4056 ( .A(\u_decoder/fir_filter/Q_data_add_3 [6]), .B(n1088), .C(
        \u_decoder/fir_filter/Q_data_add_3_buff [6]), .D(n1162), .Q(
        \u_decoder/fir_filter/n608 ) );
  INV3 U4057 ( .A(\u_decoder/fir_filter/n592 ), .Q(n2440) );
  AOI221 U4058 ( .A(\u_decoder/fir_filter/Q_data_add_2 [1]), .B(n1088), .C(
        \u_decoder/fir_filter/Q_data_add_2_buff [1]), .D(n1161), .Q(
        \u_decoder/fir_filter/n592 ) );
  INV3 U4059 ( .A(\u_decoder/fir_filter/n591 ), .Q(n2439) );
  AOI221 U4060 ( .A(\u_decoder/fir_filter/Q_data_add_2 [2]), .B(n1088), .C(
        \u_decoder/fir_filter/Q_data_add_2_buff [2]), .D(n1161), .Q(
        \u_decoder/fir_filter/n591 ) );
  INV3 U4061 ( .A(\u_decoder/fir_filter/n590 ), .Q(n2438) );
  AOI221 U4062 ( .A(\u_decoder/fir_filter/Q_data_add_2 [3]), .B(n1089), .C(
        \u_decoder/fir_filter/Q_data_add_2_buff [3]), .D(n1161), .Q(
        \u_decoder/fir_filter/n590 ) );
  INV3 U4063 ( .A(\u_decoder/fir_filter/n589 ), .Q(n2437) );
  AOI221 U4064 ( .A(\u_decoder/fir_filter/Q_data_add_2 [4]), .B(n1089), .C(
        \u_decoder/fir_filter/Q_data_add_2_buff [4]), .D(n1161), .Q(
        \u_decoder/fir_filter/n589 ) );
  INV3 U4065 ( .A(\u_decoder/fir_filter/n588 ), .Q(n2436) );
  AOI221 U4066 ( .A(\u_decoder/fir_filter/Q_data_add_2 [5]), .B(n1089), .C(
        \u_decoder/fir_filter/Q_data_add_2_buff [5]), .D(n1161), .Q(
        \u_decoder/fir_filter/n588 ) );
  INV3 U4067 ( .A(\u_decoder/fir_filter/n587 ), .Q(n2435) );
  AOI221 U4068 ( .A(\u_decoder/fir_filter/Q_data_add_2 [6]), .B(n1089), .C(
        \u_decoder/fir_filter/Q_data_add_2_buff [6]), .D(n1161), .Q(
        \u_decoder/fir_filter/n587 ) );
  INV3 U4069 ( .A(\u_decoder/fir_filter/n571 ), .Q(n2425) );
  AOI221 U4070 ( .A(\u_decoder/fir_filter/Q_data_add_1 [1]), .B(n1089), .C(
        \u_decoder/fir_filter/Q_data_add_1_buff [1]), .D(n1162), .Q(
        \u_decoder/fir_filter/n571 ) );
  INV3 U4071 ( .A(\u_decoder/fir_filter/n570 ), .Q(n2423) );
  AOI221 U4072 ( .A(\u_decoder/fir_filter/Q_data_add_1 [2]), .B(n1089), .C(
        \u_decoder/fir_filter/Q_data_add_1_buff [2]), .D(n1161), .Q(
        \u_decoder/fir_filter/n570 ) );
  INV3 U4073 ( .A(\u_decoder/fir_filter/n569 ), .Q(n2421) );
  AOI221 U4074 ( .A(\u_decoder/fir_filter/Q_data_add_1 [3]), .B(n1089), .C(
        \u_decoder/fir_filter/Q_data_add_1_buff [3]), .D(n1152), .Q(
        \u_decoder/fir_filter/n569 ) );
  INV3 U4075 ( .A(\u_decoder/fir_filter/n568 ), .Q(n2419) );
  AOI221 U4076 ( .A(\u_decoder/fir_filter/Q_data_add_1 [4]), .B(n1089), .C(
        \u_decoder/fir_filter/Q_data_add_1_buff [4]), .D(n1161), .Q(
        \u_decoder/fir_filter/n568 ) );
  INV3 U4077 ( .A(\u_decoder/fir_filter/n567 ), .Q(n2417) );
  AOI221 U4078 ( .A(\u_decoder/fir_filter/Q_data_add_1 [5]), .B(n1090), .C(
        \u_decoder/fir_filter/Q_data_add_1_buff [5]), .D(n1162), .Q(
        \u_decoder/fir_filter/n567 ) );
  INV3 U4079 ( .A(\u_decoder/fir_filter/n566 ), .Q(n2415) );
  AOI221 U4080 ( .A(\u_decoder/fir_filter/Q_data_add_1 [6]), .B(n1090), .C(
        \u_decoder/fir_filter/Q_data_add_1_buff [6]), .D(n1159), .Q(
        \u_decoder/fir_filter/n566 ) );
  OAI311 U4081 ( .A(\u_inFIFO/n551 ), .B(\u_inFIFO/sigEnableCounter ), .C(
        n2146), .D(\u_inFIFO/n552 ), .Q(\u_inFIFO/n542 ) );
  NOR31 U4082 ( .A(\u_outFIFO/i_FIFO [4]), .B(\u_outFIFO/i_FIFO [5]), .C(
        \u_outFIFO/n267 ), .Q(\u_outFIFO/n659 ) );
  XNR21 U4083 ( .A(\u_coder/n123 ), .B(\u_coder/n238 ), .Q(\u_coder/n148 ) );
  AOI211 U4084 ( .A(\u_outFIFO/currentState [1]), .B(n2217), .C(n1237), .Q(
        \u_outFIFO/n311 ) );
  OAI2111 U4085 ( .A(\u_coder/i [2]), .B(n763), .C(\u_coder/i [1]), .D(
        \u_coder/n177 ), .Q(\u_coder/n174 ) );
  AOI211 U4086 ( .A(n763), .B(\u_coder/i [2]), .C(\u_coder/i [3]), .Q(
        \u_coder/n177 ) );
  NAND41 U4087 ( .A(\u_cdr/cnt_in [0]), .B(\u_cdr/cnt_in [2]), .C(n20), .D(n50), .Q(\u_cdr/N100 ) );
  NAND41 U4088 ( .A(\u_coder/n316 ), .B(\u_coder/n317 ), .C(\u_coder/n318 ), 
        .D(\u_coder/n319 ), .Q(\u_coder/n314 ) );
  NOR21 U4089 ( .A(\u_coder/c [14]), .B(\u_coder/c [13]), .Q(\u_coder/n316 )
         );
  NOR31 U4090 ( .A(\u_coder/c [15]), .B(\u_coder/c [17]), .C(\u_coder/c [16]), 
        .Q(\u_coder/n317 ) );
  NOR40 U4091 ( .A(\u_coder/n324 ), .B(\u_coder/c [10]), .C(\u_coder/c [12]), 
        .D(\u_coder/c [11]), .Q(\u_coder/n318 ) );
  NOR21 U4092 ( .A(\u_outFIFO/k_FIFO [1]), .B(\u_outFIFO/k_FIFO [0]), .Q(
        \u_outFIFO/n661 ) );
  NOR21 U4093 ( .A(\u_outFIFO/n279 ), .B(\u_outFIFO/n280 ), .Q(
        \u_outFIFO/n1010 ) );
  NOR31 U4094 ( .A(\u_outFIFO/n276 ), .B(\u_outFIFO/i_FIFO [6]), .C(
        \u_outFIFO/n275 ), .Q(\u_outFIFO/n607 ) );
  NOR31 U4095 ( .A(\u_outFIFO/i_FIFO [4]), .B(\u_outFIFO/i_FIFO [6]), .C(
        \u_outFIFO/n275 ), .Q(\u_outFIFO/n538 ) );
  NOR31 U4096 ( .A(\u_outFIFO/i_FIFO [5]), .B(\u_outFIFO/i_FIFO [6]), .C(
        \u_outFIFO/n276 ), .Q(\u_outFIFO/n469 ) );
  NOR31 U4097 ( .A(\u_outFIFO/n276 ), .B(\u_outFIFO/i_FIFO [5]), .C(
        \u_outFIFO/n267 ), .Q(\u_outFIFO/n830 ) );
  NOR31 U4098 ( .A(\u_outFIFO/n275 ), .B(\u_outFIFO/i_FIFO [4]), .C(
        \u_outFIFO/n267 ), .Q(\u_outFIFO/n963 ) );
  NOR31 U4099 ( .A(\u_outFIFO/n275 ), .B(\u_outFIFO/n276 ), .C(
        \u_outFIFO/n267 ), .Q(\u_outFIFO/n1104 ) );
  NOR21 U4100 ( .A(\u_outFIFO/i_FIFO [1]), .B(\u_outFIFO/i_FIFO [0]), .Q(
        \u_outFIFO/n982 ) );
  AOI221 U4101 ( .A(\sig_MUX_inMUX11[0] ), .B(n2136), .C(in_MUX_inSEL11), .D(
        sig_DEMUX_outDEMUX1[3]), .Q(n3114) );
  NOR31 U4102 ( .A(n2126), .B(in_DEMUX_inSEL1[2]), .C(\u_demux1/n4 ), .Q(
        sig_DEMUX_outDEMUX1[3]) );
  NOR21 U4103 ( .A(\u_outFIFO/n279 ), .B(\u_outFIFO/i_FIFO [0]), .Q(
        \u_outFIFO/n1001 ) );
  NOR21 U4104 ( .A(\u_outFIFO/n280 ), .B(\u_outFIFO/i_FIFO [1]), .Q(
        \u_outFIFO/n992 ) );
  XNR21 U4105 ( .A(\u_coder/n238 ), .B(\u_coder/sin_was_positiveQ ), .Q(
        \u_coder/n195 ) );
  NOR31 U4106 ( .A(\u_outFIFO/i_FIFO [5]), .B(\u_outFIFO/i_FIFO [6]), .C(
        \u_outFIFO/i_FIFO [4]), .Q(\u_outFIFO/n397 ) );
  OAI2111 U4107 ( .A(n763), .B(\u_coder/n101 ), .C(\u_coder/n160 ), .D(
        \u_coder/n161 ), .Q(\u_coder/n157 ) );
  AOI311 U4108 ( .A(n763), .B(\u_coder/n103 ), .C(\u_coder/i [1]), .D(
        \u_coder/n162 ), .Q(\u_coder/n161 ) );
  NOR31 U4109 ( .A(\u_coder/n105 ), .B(\u_coder/i [3]), .C(\u_coder/i [1]), 
        .Q(\u_coder/n162 ) );
  OAI2111 U4110 ( .A(\u_coder/n105 ), .B(\u_coder/n101 ), .C(\u_coder/n159 ), 
        .D(\u_coder/n104 ), .Q(\u_coder/n155 ) );
  NAND22 U4111 ( .A(\u_coder/my_clk_10M ), .B(\u_coder/stateI[0] ), .Q(
        \u_coder/n144 ) );
  MUX22 U4112 ( .A(\u_cordic/mycordic/present_C_table[7][1] ), .B(n757), .S(
        n766), .Q(n384) );
  NOR21 U4113 ( .A(\u_outFIFO/n278 ), .B(\u_outFIFO/i_FIFO [3]), .Q(
        \u_outFIFO/n1019 ) );
  NOR21 U4114 ( .A(\u_outFIFO/n277 ), .B(\u_outFIFO/i_FIFO [2]), .Q(
        \u_outFIFO/n1052 ) );
  NOR21 U4115 ( .A(\u_outFIFO/n277 ), .B(\u_outFIFO/n278 ), .Q(
        \u_outFIFO/n1085 ) );
  OAI2111 U4116 ( .A(\u_outFIFO/n1140 ), .B(\u_outFIFO/n1141 ), .C(
        \u_outFIFO/n1115 ), .D(\u_outFIFO/n1142 ), .Q(\u_outFIFO/n1128 ) );
  NAND41 U4117 ( .A(\u_outFIFO/n263 ), .B(\u_outFIFO/n262 ), .C(
        \u_outFIFO/n261 ), .D(\u_outFIFO/n260 ), .Q(\u_outFIFO/n1140 ) );
  NAND41 U4118 ( .A(\u_outFIFO/outWriteCount[7] ), .B(\u_outFIFO/n266 ), .C(
        \u_outFIFO/n265 ), .D(\u_outFIFO/n264 ), .Q(\u_outFIFO/n1141 ) );
  NAND22 U4119 ( .A(\u_coder/stateQ[0] ), .B(\u_coder/my_clk_10M ), .Q(
        \u_coder/n183 ) );
  XNR21 U4120 ( .A(\u_decoder/iq_demod/cossin_dig/n19 ), .B(
        \u_decoder/iq_demod/cossin_dig/n21 ), .Q(
        \u_decoder/iq_demod/cossin_dig/n54 ) );
  NAND22 U4121 ( .A(\u_coder/isPositiveQ ), .B(\u_coder/is9 ), .Q(
        \u_coder/n191 ) );
  XNR21 U4122 ( .A(n385), .B(n3112), .Q(\u_coder/n238 ) );
  NOR21 U4123 ( .A(\u_inFIFO/j_FIFO [3]), .B(\u_inFIFO/j_FIFO [2]), .Q(
        \u_inFIFO/n475 ) );
  INV3 U4124 ( .A(\u_cdr/n33 ), .Q(n1806) );
  AOI2111 U4125 ( .A(\u_coder/n120 ), .B(\u_coder/j [3]), .C(\u_coder/n203 ), 
        .D(n2183), .Q(\u_coder/n201 ) );
  AOI211 U4126 ( .A(\u_coder/j [0]), .B(n762), .C(\u_coder/n118 ), .Q(
        \u_coder/n203 ) );
  INV3 U4127 ( .A(\u_coder/n204 ), .Q(n2183) );
  AOI311 U4128 ( .A(\u_coder/j [0]), .B(\u_coder/n118 ), .C(n762), .D(
        \u_coder/n205 ), .Q(\u_coder/n204 ) );
  AOI221 U4129 ( .A(\sig_MUX_inMUX4[0] ), .B(n2131), .C(in_MUX_inSEL3), .D(
        sig_DEMUX_outDEMUX1[1]), .Q(n3112) );
  NOR31 U4130 ( .A(\u_demux1/n4 ), .B(in_DEMUX_inSEL1[2]), .C(
        in_DEMUX_inSEL1[1]), .Q(sig_DEMUX_outDEMUX1[1]) );
  NOR21 U4131 ( .A(\u_inFIFO/n206 ), .B(\u_inFIFO/j_FIFO [0]), .Q(
        \u_inFIFO/n481 ) );
  NOR21 U4132 ( .A(\u_inFIFO/j_FIFO [1]), .B(\u_inFIFO/j_FIFO [0]), .Q(
        \u_inFIFO/n474 ) );
  NOR21 U4133 ( .A(\u_inFIFO/n207 ), .B(\u_inFIFO/j_FIFO [1]), .Q(
        \u_inFIFO/n478 ) );
  NOR21 U4134 ( .A(\u_coder/n126 ), .B(\u_coder/n128 ), .Q(\u_coder/n149 ) );
  INV3 U4135 ( .A(n2725), .Q(n2157) );
  NAND41 U4136 ( .A(n2724), .B(n2723), .C(n2722), .D(n2721), .Q(n2725) );
  NOR40 U4137 ( .A(\u_coder/i [4]), .B(\u_coder/i [19]), .C(\u_coder/i [18]), 
        .D(\u_coder/i [17]), .Q(n2722) );
  NOR40 U4138 ( .A(\u_coder/i [16]), .B(\u_coder/i [15]), .C(\u_coder/i [14]), 
        .D(\u_coder/i [13]), .Q(n2723) );
  NAND22 U4139 ( .A(\u_coder/n103 ), .B(\u_coder/n104 ), .Q(\u_coder/n150 ) );
  NOR21 U4140 ( .A(\u_inFIFO/n206 ), .B(\u_inFIFO/n207 ), .Q(\u_inFIFO/n484 )
         );
  NAND31 U4141 ( .A(\u_cdr/cnt_d [1]), .B(\u_cdr/cnt_d [0]), .C(\u_cdr/flag ), 
        .Q(\u_cdr/n38 ) );
  NOR40 U4142 ( .A(\u_coder/i [12]), .B(\u_coder/i [11]), .C(\u_coder/i [10]), 
        .D(n2166), .Q(n2724) );
  INV3 U4143 ( .A(n2719), .Q(n2166) );
  OAI311 U4144 ( .A(n763), .B(\u_coder/i [2]), .C(\u_coder/i [1]), .D(
        \u_coder/i [3]), .Q(n2719) );
  NAND22 U4145 ( .A(\u_inFIFO/n555 ), .B(\u_inFIFO/n556 ), .Q(\u_inFIFO/n550 )
         );
  NOR40 U4146 ( .A(\u_inFIFO/outWriteCount[2] ), .B(
        \u_inFIFO/outWriteCount[1] ), .C(\u_inFIFO/outWriteCount[0] ), .D(
        \u_inFIFO/n179 ), .Q(\u_inFIFO/n555 ) );
  NOR40 U4147 ( .A(\u_inFIFO/outWriteCount[6] ), .B(
        \u_inFIFO/outWriteCount[5] ), .C(\u_inFIFO/outWriteCount[4] ), .D(
        \u_inFIFO/outWriteCount[3] ), .Q(\u_inFIFO/n556 ) );
  AOI221 U4148 ( .A(\u_coder/isPositiveQ ), .B(n2173), .C(n2185), .D(
        \u_coder/n228 ), .Q(\u_coder/n229 ) );
  NOR21 U4149 ( .A(\u_coder/j [2]), .B(n762), .Q(\u_coder/n190 ) );
  AOI221 U4150 ( .A(n2168), .B(\u_coder/n247 ), .C(\u_coder/isPositiveI ), .D(
        n2161), .Q(\u_coder/n248 ) );
  NAND22 U4151 ( .A(\u_coder/is9 ), .B(\u_coder/n191 ), .Q(\u_coder/n181 ) );
  NOR21 U4152 ( .A(\u_coder/n128 ), .B(\u_coder/n149 ), .Q(\u_coder/n137 ) );
  NAND31 U4153 ( .A(\u_coder/n105 ), .B(\u_coder/n101 ), .C(n2167), .Q(
        \u_coder/n159 ) );
  NOR40 U4154 ( .A(\u_coder/j [17]), .B(\u_coder/j [16]), .C(\u_coder/j [15]), 
        .D(\u_coder/j [14]), .Q(\u_coder/n328 ) );
  NOR40 U4155 ( .A(\u_coder/j [12]), .B(\u_coder/j [11]), .C(\u_coder/j [10]), 
        .D(n2180), .Q(n2717) );
  INV3 U4156 ( .A(n2712), .Q(n2180) );
  OAI311 U4157 ( .A(\u_coder/j [0]), .B(\u_coder/j [2]), .C(n762), .D(
        \u_coder/j [3]), .Q(n2712) );
  XNR21 U4158 ( .A(\u_outFIFO/outWriteCount[0] ), .B(n130), .Q(
        \u_outFIFO/N143 ) );
  XNR21 U4159 ( .A(\u_inFIFO/outWriteCount[0] ), .B(n129), .Q(\u_inFIFO/N133 )
         );
  NOR40 U4160 ( .A(\u_coder/j [7]), .B(n2178), .C(\u_coder/j [6]), .D(
        \u_coder/j [5]), .Q(n2714) );
  INV3 U4161 ( .A(n2713), .Q(n2178) );
  NOR21 U4162 ( .A(\u_coder/j [9]), .B(\u_coder/j [8]), .Q(n2713) );
  NOR40 U4163 ( .A(\u_coder/i [7]), .B(n2163), .C(\u_coder/i [6]), .D(
        \u_coder/i [5]), .Q(n2721) );
  INV3 U4164 ( .A(n2720), .Q(n2163) );
  NOR21 U4165 ( .A(\u_coder/i [9]), .B(\u_coder/i [8]), .Q(n2720) );
  NOR21 U4166 ( .A(\u_inFIFO/n205 ), .B(\u_inFIFO/j_FIFO [3]), .Q(
        \u_inFIFO/n487 ) );
  NOR21 U4167 ( .A(\u_inFIFO/n204 ), .B(\u_inFIFO/j_FIFO [2]), .Q(
        \u_inFIFO/n496 ) );
  OAI2111 U4168 ( .A(\u_coder/n94 ), .B(\u_coder/n223 ), .C(\u_coder/n224 ), 
        .D(\u_coder/n225 ), .Q(\u_coder/n340 ) );
  NAND41 U4169 ( .A(n1212), .B(\u_coder/is9 ), .C(\u_coder/stateQ[0] ), .D(
        \u_coder/stateI[0] ), .Q(\u_coder/n225 ) );
  OAI2111 U4170 ( .A(\u_coder/n209 ), .B(\u_coder/n223 ), .C(\u_coder/n224 ), 
        .D(\u_coder/n240 ), .Q(\u_coder/n346 ) );
  NAND31 U4171 ( .A(\u_coder/n236 ), .B(\u_coder/n167 ), .C(
        \sig_MUX_inMUX3[0] ), .Q(\u_coder/n240 ) );
  NOR40 U4172 ( .A(\u_coder/n320 ), .B(n2202), .C(\u_coder/c [19]), .D(
        \u_coder/c [18]), .Q(\u_coder/n319 ) );
  INV3 U4173 ( .A(\u_coder/n321 ), .Q(n2202) );
  NAND22 U4174 ( .A(\u_coder/n322 ), .B(\u_coder/n323 ), .Q(\u_coder/n320 ) );
  NOR31 U4175 ( .A(\u_coder/c [1]), .B(\u_coder/c [4]), .C(\u_coder/c [3]), 
        .Q(\u_coder/n321 ) );
  INV3 U4176 ( .A(\u_inFIFO/n547 ), .Q(n1822) );
  AOI221 U4177 ( .A(n129), .B(n2094), .C(\u_inFIFO/outReadCount[0] ), .D(
        \u_inFIFO/n542 ), .Q(\u_inFIFO/n547 ) );
  INV3 U4178 ( .A(\u_inFIFO/n546 ), .Q(n1823) );
  AOI221 U4179 ( .A(\u_inFIFO/N119 ), .B(n2094), .C(\u_inFIFO/outReadCount[1] ), .D(\u_inFIFO/n542 ), .Q(\u_inFIFO/n546 ) );
  INV3 U4180 ( .A(\u_inFIFO/n545 ), .Q(n1824) );
  AOI221 U4181 ( .A(\u_inFIFO/N120 ), .B(n2094), .C(\u_inFIFO/outReadCount[2] ), .D(\u_inFIFO/n542 ), .Q(\u_inFIFO/n545 ) );
  INV3 U4182 ( .A(\u_inFIFO/n544 ), .Q(n1825) );
  AOI221 U4183 ( .A(\u_inFIFO/N121 ), .B(n2094), .C(\u_inFIFO/outReadCount[3] ), .D(\u_inFIFO/n542 ), .Q(\u_inFIFO/n544 ) );
  INV3 U4184 ( .A(\u_inFIFO/n543 ), .Q(n1826) );
  AOI221 U4185 ( .A(\u_inFIFO/N122 ), .B(n2094), .C(\u_inFIFO/outReadCount[4] ), .D(\u_inFIFO/n542 ), .Q(\u_inFIFO/n543 ) );
  NOR21 U4186 ( .A(\u_inFIFO/n204 ), .B(\u_inFIFO/n205 ), .Q(\u_inFIFO/n505 )
         );
  NAND31 U4187 ( .A(\u_inFIFO/j_FIFO [5]), .B(\u_inFIFO/j_FIFO [4]), .C(
        \u_inFIFO/j_FIFO [6]), .Q(\u_inFIFO/n473 ) );
  NAND31 U4188 ( .A(\u_inFIFO/j_FIFO [5]), .B(\u_inFIFO/n203 ), .C(
        \u_inFIFO/j_FIFO [6]), .Q(\u_inFIFO/n440 ) );
  NAND31 U4189 ( .A(\u_inFIFO/j_FIFO [4]), .B(\u_inFIFO/n202 ), .C(
        \u_inFIFO/j_FIFO [6]), .Q(\u_inFIFO/n407 ) );
  NAND31 U4190 ( .A(\u_inFIFO/n203 ), .B(\u_inFIFO/n202 ), .C(
        \u_inFIFO/j_FIFO [6]), .Q(\u_inFIFO/n374 ) );
  NOR21 U4191 ( .A(n1236), .B(\u_outFIFO/sigEnableCounter ), .Q(
        \u_outFIFO/n1142 ) );
  NAND31 U4192 ( .A(\u_inFIFO/j_FIFO [4]), .B(\u_inFIFO/n201 ), .C(
        \u_inFIFO/j_FIFO [5]), .Q(\u_inFIFO/n341 ) );
  NAND31 U4193 ( .A(\u_inFIFO/n203 ), .B(\u_inFIFO/n201 ), .C(
        \u_inFIFO/j_FIFO [5]), .Q(\u_inFIFO/n308 ) );
  NAND31 U4194 ( .A(\u_inFIFO/n202 ), .B(\u_inFIFO/n201 ), .C(
        \u_inFIFO/j_FIFO [4]), .Q(\u_inFIFO/n275 ) );
  NAND22 U4195 ( .A(n2218), .B(\u_outFIFO/n257 ), .Q(\u_outFIFO/n1115 ) );
  XNR21 U4196 ( .A(\u_cordic/mycordic/present_Q_table[0][7] ), .B(
        \u_cordic/mycordic/sub_add_151_b0/carry [7]), .Q(
        \u_cordic/mycordic/N247 ) );
  INV3 U4197 ( .A(\u_cordic/mycordic/n514 ), .Q(n1458) );
  AOI221 U4198 ( .A(\u_cordic/mycordic/N337 ), .B(\u_cordic/mycordic/n336 ), 
        .C(\u_cordic/mycordic/N369 ), .D(n1904), .Q(\u_cordic/mycordic/n514 )
         );
  XNR21 U4199 ( .A(\u_cordic/mycordic/present_ANGLE_table[1][5] ), .B(
        \u_cordic/mycordic/sub_196/carry[5] ), .Q(\u_cordic/mycordic/N369 ) );
  XOR21 U4200 ( .A(\u_cordic/mycordic/present_ANGLE_table[1][5] ), .B(
        \u_cordic/mycordic/add_191/carry[5] ), .Q(\u_cordic/mycordic/N337 ) );
  NAND31 U4201 ( .A(\u_inFIFO/n202 ), .B(\u_inFIFO/n201 ), .C(\u_inFIFO/n203 ), 
        .Q(\u_inFIFO/n227 ) );
  NOR31 U4202 ( .A(\u_coder/n256 ), .B(\u_coder/n150 ), .C(\u_coder/n105 ), 
        .Q(\u_coder/n261 ) );
  INV3 U4203 ( .A(\u_cordic/mycordic/n448 ), .Q(n1442) );
  AOI221 U4204 ( .A(\u_cordic/mycordic/N539 ), .B(n771), .C(
        \u_cordic/mycordic/N555 ), .D(n1903), .Q(\u_cordic/mycordic/n448 ) );
  XNR21 U4205 ( .A(\u_cordic/mycordic/present_ANGLE_table[5][5] ), .B(
        \u_cordic/mycordic/sub_236/carry [5]), .Q(\u_cordic/mycordic/N555 ) );
  XOR21 U4206 ( .A(\u_cordic/mycordic/present_ANGLE_table[5][5] ), .B(
        \u_cordic/mycordic/add_233/carry [5]), .Q(\u_cordic/mycordic/N539 ) );
  INV3 U4207 ( .A(\u_cordic/mycordic/n447 ), .Q(n1443) );
  AOI221 U4208 ( .A(\u_cordic/mycordic/N540 ), .B(n770), .C(
        \u_cordic/mycordic/N556 ), .D(n1903), .Q(\u_cordic/mycordic/n447 ) );
  XNR21 U4209 ( .A(\u_cordic/mycordic/present_ANGLE_table[5][6] ), .B(
        \u_cordic/mycordic/sub_236/carry [6]), .Q(\u_cordic/mycordic/N556 ) );
  XOR21 U4210 ( .A(\u_cordic/mycordic/present_ANGLE_table[5][6] ), .B(
        \u_cordic/mycordic/add_233/carry [6]), .Q(\u_cordic/mycordic/N540 ) );
  INV3 U4211 ( .A(\u_cordic/mycordic/n446 ), .Q(n1444) );
  AOI221 U4212 ( .A(\u_cordic/mycordic/N541 ), .B(n771), .C(
        \u_cordic/mycordic/N557 ), .D(n1903), .Q(\u_cordic/mycordic/n446 ) );
  XNR21 U4213 ( .A(\u_cordic/mycordic/present_ANGLE_table[5][7] ), .B(
        \u_cordic/mycordic/sub_236/carry [7]), .Q(\u_cordic/mycordic/N557 ) );
  XOR21 U4214 ( .A(\u_cordic/mycordic/present_ANGLE_table[5][7] ), .B(
        \u_cordic/mycordic/add_233/carry [7]), .Q(\u_cordic/mycordic/N541 ) );
  INV3 U4215 ( .A(\u_cordic/mycordic/n445 ), .Q(n1445) );
  AOI221 U4216 ( .A(\u_cordic/mycordic/N542 ), .B(n770), .C(
        \u_cordic/mycordic/N558 ), .D(n1903), .Q(\u_cordic/mycordic/n445 ) );
  XNR21 U4217 ( .A(\u_cordic/mycordic/present_ANGLE_table[5][8] ), .B(
        \u_cordic/mycordic/sub_236/carry [8]), .Q(\u_cordic/mycordic/N558 ) );
  XOR21 U4218 ( .A(\u_cordic/mycordic/present_ANGLE_table[5][8] ), .B(
        \u_cordic/mycordic/add_233/carry [8]), .Q(\u_cordic/mycordic/N542 ) );
  NAND22 U4219 ( .A(n2108), .B(n1217), .Q(\u_outFIFO/n315 ) );
  INV3 U4220 ( .A(n3116), .Q(n2108) );
  AOI221 U4221 ( .A(\sig_MUX_inMUX13[0] ), .B(n2137), .C(in_MUX_inSEL12), .D(
        sig_DEMUX_outDEMUX2[4]), .Q(n3116) );
  NOR31 U4222 ( .A(n3118), .B(in_DEMUX_inSEL2[1]), .C(n2128), .Q(
        sig_DEMUX_outDEMUX2[4]) );
  NAND31 U4223 ( .A(n1219), .B(\u_cdr/n38 ), .C(\u_cdr/flag ), .Q(\u_cdr/n35 )
         );
  BUF2 U4224 ( .A(\u_inFIFO/N40 ), .Q(n1202) );
  INV3 U4225 ( .A(\u_outFIFO/N216 ), .Q(n2216) );
  INV3 U4226 ( .A(\u_outFIFO/N217 ), .Q(n2215) );
  INV3 U4227 ( .A(\u_outFIFO/N218 ), .Q(n2214) );
  INV3 U4228 ( .A(\u_outFIFO/N130 ), .Q(n2234) );
  NOR31 U4229 ( .A(\u_cordic/n11 ), .B(\u_cordic/present_state [1]), .C(
        \u_cordic/n9 ), .Q(\sig_MUX_inMUX11[0] ) );
  AOI211 U4230 ( .A(\u_cdr/cnt_d [1]), .B(n1219), .C(\u_cdr/n27 ), .Q(
        \u_cdr/n42 ) );
  INV3 U4231 ( .A(\u_decoder/iq_demod/cossin_dig/n35 ), .Q(n2683) );
  AOI211 U4232 ( .A(\u_decoder/iq_demod/sin_out [2]), .B(n756), .C(
        \u_decoder/iq_demod/cossin_dig/n34 ), .Q(
        \u_decoder/iq_demod/cossin_dig/n35 ) );
  INV3 U4233 ( .A(\u_decoder/iq_demod/cossin_dig/n33 ), .Q(n2682) );
  AOI211 U4234 ( .A(\u_decoder/iq_demod/sin_out [1]), .B(n756), .C(
        \u_decoder/iq_demod/cossin_dig/n34 ), .Q(
        \u_decoder/iq_demod/cossin_dig/n33 ) );
  NOR21 U4235 ( .A(\u_outFIFO/n664 ), .B(\u_outFIFO/n666 ), .Q(
        \u_outFIFO/n1116 ) );
  INV3 U4236 ( .A(\u_coder/n148 ), .Q(n2095) );
  BUF2 U4237 ( .A(\u_outFIFO/N42 ), .Q(n1183) );
  OAI311 U4238 ( .A(n20), .B(\u_cdr/cnt_in [0]), .C(\u_cdr/n30 ), .D(n1225), 
        .Q(\u_cdr/n28 ) );
  NAND22 U4239 ( .A(n1218), .B(\u_coder/old_i_data ), .Q(\u_coder/n258 ) );
  INV3 U4240 ( .A(\u_coder/n257 ), .Q(n2160) );
  NAND22 U4241 ( .A(\u_cdr/cnt_in [2]), .B(\u_cdr/N100 ), .Q(
        \u_cdr/dp_cluster_0/mult_add_59_aco/PROD_not[2] ) );
  OAI311 U4242 ( .A(n289), .B(\u_cdr/cnt_in [1]), .C(\u_cdr/n30 ), .D(n1225), 
        .Q(\u_cdr/n31 ) );
  NAND22 U4243 ( .A(\u_cdr/cnt_in [0]), .B(\u_cdr/N100 ), .Q(
        \u_cdr/dp_cluster_0/mult_add_59_aco/PROD_not[0] ) );
  NAND41 U4244 ( .A(\u_cdr/cnt [1]), .B(\u_cdr/cnt [0]), .C(\u_cdr/n33 ), .D(
        \u_cdr/n16 ), .Q(\u_cdr/n37 ) );
  AOI211 U4245 ( .A(\u_cdr/n33 ), .B(\u_cdr/n17 ), .C(\u_cdr/n34 ), .Q(
        \u_cdr/n36 ) );
  BUF2 U4246 ( .A(\u_cordic/mycordic/n108 ), .Q(n757) );
  OAI311 U4247 ( .A(\u_decoder/fir_filter/n1150 ), .B(
        \u_decoder/fir_filter/n1149 ), .C(\u_decoder/fir_filter/n1151 ), .D(
        \u_decoder/fir_filter/n1152 ), .Q(\u_decoder/fir_filter/n1451 ) );
  NAND22 U4248 ( .A(\sig_MUX_inMUX8[0] ), .B(\u_decoder/fir_filter/n1150 ), 
        .Q(\u_decoder/fir_filter/n1152 ) );
  NOR21 U4249 ( .A(n1167), .B(\u_decoder/fir_filter/n1151 ), .Q(
        \u_decoder/fir_filter/n1150 ) );
  NAND22 U4250 ( .A(\u_coder/n261 ), .B(\u_coder/i [3]), .Q(\u_coder/n242 ) );
  OAI311 U4251 ( .A(n290), .B(\u_cdr/n23 ), .C(\u_cdr/n24 ), .D(\u_cdr/n25 ), 
        .Q(\u_cdr/n50 ) );
  MAJ31 U4252 ( .A(\u_cdr/n20 ), .B(\u_cdr/n19 ), .C(\u_cdr/n3 ), .Q(
        \u_cdr/n23 ) );
  NOR21 U4253 ( .A(\u_cdr/cnt_in [2]), .B(n1238), .Q(\u_cdr/n26 ) );
  NAND22 U4254 ( .A(\u_outFIFO/outReadCount[0] ), .B(\u_outFIFO/n266 ), .Q(
        n2761) );
  XNR21 U4255 ( .A(\u_cordic/mycordic/r173/carry [4]), .B(n387), .Q(n386) );
  XNR21 U4256 ( .A(\u_cordic/mycordic/r173/carry [7]), .B(n389), .Q(n388) );
  NAND22 U4257 ( .A(\u_outFIFO/outReadCount[6] ), .B(\u_outFIFO/n260 ), .Q(
        n2759) );
  NAND31 U4258 ( .A(n2185), .B(\u_coder/n117 ), .C(n2176), .Q(\u_coder/n260 )
         );
  NAND22 U4259 ( .A(\u_outFIFO/outReadCount[5] ), .B(\u_outFIFO/n261 ), .Q(
        n2757) );
  NOR31 U4260 ( .A(\u_coder/c [7]), .B(\u_coder/c [9]), .C(\u_coder/c [8]), 
        .Q(\u_coder/n323 ) );
  AOI221 U4261 ( .A(\u_outFIFO/n266 ), .B(n1912), .C(\u_outFIFO/N143 ), .D(
        \u_outFIFO/n1131 ), .Q(\u_outFIFO/n1137 ) );
  AOI221 U4262 ( .A(\u_outFIFO/N120 ), .B(n1912), .C(\u_outFIFO/N144 ), .D(
        \u_outFIFO/n1131 ), .Q(\u_outFIFO/n1136 ) );
  AOI221 U4263 ( .A(\u_outFIFO/N121 ), .B(n1912), .C(\u_outFIFO/N145 ), .D(
        \u_outFIFO/n1131 ), .Q(\u_outFIFO/n1135 ) );
  AOI221 U4264 ( .A(\u_outFIFO/N122 ), .B(n1912), .C(\u_outFIFO/N146 ), .D(
        \u_outFIFO/n1131 ), .Q(\u_outFIFO/n1134 ) );
  INV3 U4265 ( .A(\u_cordic/mycordic/n498 ), .Q(n1551) );
  AOI221 U4266 ( .A(\u_cordic/mycordic/N401 ), .B(n778), .C(
        \u_cordic/mycordic/N433 ), .D(n1908), .Q(\u_cordic/mycordic/n498 ) );
  XNR21 U4267 ( .A(\u_cordic/mycordic/present_ANGLE_table[2][5] ), .B(
        \u_cordic/mycordic/sub_207/carry [5]), .Q(\u_cordic/mycordic/N433 ) );
  XOR21 U4268 ( .A(\u_cordic/mycordic/present_ANGLE_table[2][5] ), .B(
        \u_cordic/mycordic/add_202/carry [5]), .Q(\u_cordic/mycordic/N401 ) );
  INV3 U4269 ( .A(\u_cordic/mycordic/n483 ), .Q(n1525) );
  AOI221 U4270 ( .A(\u_cordic/mycordic/N460 ), .B(n777), .C(
        \u_cordic/mycordic/N488 ), .D(n1907), .Q(\u_cordic/mycordic/n483 ) );
  XNR21 U4271 ( .A(\u_cordic/mycordic/present_ANGLE_table[3][4] ), .B(
        \u_cordic/mycordic/sub_218/carry[4] ), .Q(\u_cordic/mycordic/N488 ) );
  XOR21 U4272 ( .A(\u_cordic/mycordic/present_ANGLE_table[3][4] ), .B(
        \u_cordic/mycordic/add_213/carry[4] ), .Q(\u_cordic/mycordic/N460 ) );
  AOI221 U4273 ( .A(\u_inFIFO/n188 ), .B(\u_inFIFO/n533 ), .C(\u_inFIFO/N133 ), 
        .D(\u_inFIFO/n534 ), .Q(\u_inFIFO/n540 ) );
  AOI221 U4274 ( .A(\u_inFIFO/N143 ), .B(\u_inFIFO/n533 ), .C(\u_inFIFO/N134 ), 
        .D(\u_inFIFO/n534 ), .Q(\u_inFIFO/n532 ) );
  AOI221 U4275 ( .A(\u_inFIFO/N144 ), .B(\u_inFIFO/n533 ), .C(\u_inFIFO/N135 ), 
        .D(\u_inFIFO/n534 ), .Q(\u_inFIFO/n535 ) );
  AOI221 U4276 ( .A(\u_inFIFO/N145 ), .B(\u_inFIFO/n533 ), .C(\u_inFIFO/N136 ), 
        .D(\u_inFIFO/n534 ), .Q(\u_inFIFO/n536 ) );
  NAND41 U4277 ( .A(n1212), .B(\u_coder/IorQ ), .C(\u_coder/n235 ), .D(
        \u_coder/n309 ), .Q(\u_coder/n308 ) );
  NOR21 U4278 ( .A(n2161), .B(n2173), .Q(\u_coder/n307 ) );
  NAND22 U4279 ( .A(\u_outFIFO/outReadCount[3] ), .B(\u_outFIFO/n263 ), .Q(
        n2750) );
  AOI2111 U4280 ( .A(\u_cdr/n39 ), .B(\u_cdr/n40 ), .C(n1240), .D(\u_cdr/n41 ), 
        .Q(\u_cdr/n53 ) );
  NOR31 U4281 ( .A(\u_cdr/n16 ), .B(\u_cdr/cnt [1]), .C(\u_cdr/cnt [0]), .Q(
        \u_cdr/n41 ) );
  NAND22 U4282 ( .A(\u_cdr/flag ), .B(n3114), .Q(\u_cdr/n40 ) );
  NAND22 U4283 ( .A(\u_outFIFO/outReadCount[2] ), .B(\u_outFIFO/n264 ), .Q(
        n2747) );
  NOR21 U4284 ( .A(\u_decoder/iq_demod/cossin_dig/n56 ), .B(
        \u_decoder/iq_demod/cossin_dig/n31 ), .Q(
        \u_decoder/iq_demod/cossin_dig/n34 ) );
  NAND22 U4285 ( .A(\u_outFIFO/outReadCount[4] ), .B(\u_outFIFO/n262 ), .Q(
        n2751) );
  INV3 U4286 ( .A(n2718), .Q(n2170) );
  NAND41 U4287 ( .A(n2717), .B(n2716), .C(n2715), .D(n2714), .Q(n2718) );
  NOR40 U4288 ( .A(\u_coder/j [4]), .B(\u_coder/j [19]), .C(\u_coder/j [18]), 
        .D(\u_coder/j [17]), .Q(n2715) );
  NOR40 U4289 ( .A(\u_coder/j [16]), .B(\u_coder/j [15]), .C(\u_coder/j [14]), 
        .D(\u_coder/j [13]), .Q(n2716) );
  INV3 U4290 ( .A(\u_coder/n220 ), .Q(n2181) );
  OAI2111 U4291 ( .A(\u_coder/j [2]), .B(\u_coder/j [0]), .C(n762), .D(
        \u_coder/n221 ), .Q(\u_coder/n220 ) );
  AOI211 U4292 ( .A(\u_coder/j [0]), .B(\u_coder/j [2]), .C(\u_coder/j [3]), 
        .Q(\u_coder/n221 ) );
  NOR31 U4293 ( .A(\u_coder/n120 ), .B(\u_coder/j [3]), .C(n762), .Q(
        \u_coder/n205 ) );
  BUF2 U4294 ( .A(\u_inFIFO/n522 ), .Q(n912) );
  NOR21 U4295 ( .A(n1235), .B(\u_inFIFO/sigEnableCounter ), .Q(\u_inFIFO/n522 ) );
  NOR21 U4296 ( .A(n895), .B(\u_coder/c [0]), .Q(\u_coder/N503 ) );
  BUF2 U4297 ( .A(\u_inFIFO/N41 ), .Q(n765) );
  NAND22 U4298 ( .A(\u_cdr/N100 ), .B(\u_cdr/cnt_in [3]), .Q(
        \u_cdr/dp_cluster_0/mult_add_59_aco/PROD_not[3] ) );
  INV3 U4299 ( .A(\u_cdr/dp_cluster_0/mult_add_59_aco/PROD_not[1] ), .Q(n2211)
         );
  NAND22 U4300 ( .A(\u_cdr/cnt_in [1]), .B(\u_cdr/N100 ), .Q(
        \u_cdr/dp_cluster_0/mult_add_59_aco/PROD_not[1] ) );
  XNR21 U4301 ( .A(\u_cordic/mycordic/add_262/carry [5]), .B(
        \u_cordic/mycordic/present_ANGLE_table[6][5] ), .Q(
        \u_cordic/mycordic/N620 ) );
  XOR21 U4302 ( .A(\u_cordic/mycordic/add_262/carry [7]), .B(
        \u_cordic/mycordic/present_ANGLE_table[6][7] ), .Q(
        \u_cordic/mycordic/N622 ) );
  XNR21 U4303 ( .A(\u_cordic/mycordic/add_262/carry [6]), .B(
        \u_cordic/mycordic/present_ANGLE_table[6][6] ), .Q(
        \u_cordic/mycordic/N621 ) );
  XNR21 U4304 ( .A(\u_cordic/mycordic/add_262/carry [8]), .B(
        \u_cordic/mycordic/present_ANGLE_table[6][8] ), .Q(
        \u_cordic/mycordic/N623 ) );
  INV3 U4305 ( .A(\u_decoder/fir_filter/n1102 ), .Q(n2638) );
  NAND22 U4306 ( .A(\u_decoder/fir_filter/I_data_mult_2_buff [0]), .B(n1158), 
        .Q(\u_decoder/fir_filter/n1102 ) );
  INV3 U4307 ( .A(\u_cordic/mycordic/n436 ), .Q(n1902) );
  NAND22 U4308 ( .A(\u_cordic/mycordic/next_ANGLE_table[6][0] ), .B(n1213), 
        .Q(\u_cordic/mycordic/n436 ) );
  INV3 U4309 ( .A(\u_cordic/mycordic/n424 ), .Q(n1893) );
  NAND22 U4310 ( .A(\u_cordic/mycordic/next_ANGLE_table[6][1] ), .B(n1213), 
        .Q(\u_cordic/mycordic/n424 ) );
  NAND22 U4311 ( .A(\u_coder/c [2]), .B(\u_coder/n33 ), .Q(\u_coder/n324 ) );
  INV3 U4312 ( .A(\u_coder/n310 ), .Q(n2174) );
  NAND31 U4313 ( .A(\u_coder/j [2]), .B(n2177), .C(\u_coder/n311 ), .Q(
        \u_coder/n310 ) );
  NOR31 U4314 ( .A(\u_coder/j [0]), .B(\u_coder/j [3]), .C(n762), .Q(
        \u_coder/n311 ) );
  NAND22 U4315 ( .A(\u_coder/n261 ), .B(\u_coder/n101 ), .Q(\u_coder/n259 ) );
  NOR31 U4316 ( .A(\u_outFIFO/n284 ), .B(\u_outFIFO/n285 ), .C(
        \u_outFIFO/n1153 ), .Q(\u_outFIFO/N198 ) );
  INV3 U4317 ( .A(n2726), .Q(n2171) );
  NOR21 U4318 ( .A(\u_coder/j [18]), .B(\u_coder/j [17]), .Q(n2726) );
  XNR21 U4319 ( .A(\u_cordic/mycordic/r173/carry [5]), .B(n391), .Q(n390) );
  INV3 U4320 ( .A(\u_cordic/mycordic/n407 ), .Q(n1876) );
  NAND22 U4321 ( .A(\u_cordic/mycordic/next_ANGLE_table[6][7] ), .B(n1215), 
        .Q(\u_cordic/mycordic/n407 ) );
  INV3 U4322 ( .A(\u_cordic/mycordic/n413 ), .Q(n1882) );
  NAND22 U4323 ( .A(\u_cordic/mycordic/next_ANGLE_table[6][2] ), .B(n1214), 
        .Q(\u_cordic/mycordic/n413 ) );
  XNR21 U4324 ( .A(\u_cordic/mycordic/r173/carry [6]), .B(
        \u_cordic/mycordic/present_ANGLE_table[6][6] ), .Q(n392) );
  INV3 U4325 ( .A(\u_outFIFO/N131 ), .Q(n2233) );
  INV3 U4326 ( .A(\u_outFIFO/n1126 ), .Q(n1798) );
  AOI221 U4327 ( .A(n130), .B(\u_outFIFO/n1119 ), .C(
        \u_outFIFO/outReadCount[0] ), .D(\u_outFIFO/n1120 ), .Q(
        \u_outFIFO/n1126 ) );
  INV3 U4328 ( .A(\u_outFIFO/n1125 ), .Q(n1799) );
  AOI221 U4329 ( .A(\u_outFIFO/N136 ), .B(\u_outFIFO/n1119 ), .C(
        \u_outFIFO/outReadCount[1] ), .D(\u_outFIFO/n1120 ), .Q(
        \u_outFIFO/n1125 ) );
  INV3 U4330 ( .A(\u_outFIFO/n1124 ), .Q(n1800) );
  AOI221 U4331 ( .A(\u_outFIFO/N137 ), .B(\u_outFIFO/n1119 ), .C(
        \u_outFIFO/outReadCount[2] ), .D(\u_outFIFO/n1120 ), .Q(
        \u_outFIFO/n1124 ) );
  INV3 U4332 ( .A(\u_outFIFO/n1123 ), .Q(n1801) );
  AOI221 U4333 ( .A(\u_outFIFO/N138 ), .B(\u_outFIFO/n1119 ), .C(
        \u_outFIFO/outReadCount[3] ), .D(\u_outFIFO/n1120 ), .Q(
        \u_outFIFO/n1123 ) );
  INV3 U4334 ( .A(\u_outFIFO/n1122 ), .Q(n1802) );
  AOI221 U4335 ( .A(\u_outFIFO/N139 ), .B(\u_outFIFO/n1119 ), .C(
        \u_outFIFO/outReadCount[4] ), .D(\u_outFIFO/n1120 ), .Q(
        \u_outFIFO/n1122 ) );
  INV3 U4336 ( .A(\u_coder/n237 ), .Q(n1812) );
  AOI221 U4337 ( .A(\u_coder/isPositiveQ ), .B(\u_coder/n236 ), .C(n2097), .D(
        \u_coder/n209 ), .Q(\u_coder/n237 ) );
  INV3 U4338 ( .A(\u_outFIFO/n309 ), .Q(n1584) );
  AOI221 U4339 ( .A(\u_outFIFO/N202 ), .B(\u_outFIFO/n310 ), .C(
        sig_outFIFO_outData[3]), .D(\u_outFIFO/n311 ), .Q(\u_outFIFO/n309 ) );
  INV3 U4340 ( .A(\u_outFIFO/n312 ), .Q(n1583) );
  AOI221 U4341 ( .A(\u_outFIFO/N203 ), .B(\u_outFIFO/n310 ), .C(
        sig_outFIFO_outData[2]), .D(\u_outFIFO/n311 ), .Q(\u_outFIFO/n312 ) );
  INV3 U4342 ( .A(\u_outFIFO/n313 ), .Q(n1582) );
  AOI221 U4343 ( .A(\u_outFIFO/N204 ), .B(\u_outFIFO/n310 ), .C(
        sig_outFIFO_outData[1]), .D(\u_outFIFO/n311 ), .Q(\u_outFIFO/n313 ) );
  INV3 U4344 ( .A(\u_outFIFO/n314 ), .Q(n1581) );
  AOI221 U4345 ( .A(\u_outFIFO/N205 ), .B(\u_outFIFO/n310 ), .C(
        sig_outFIFO_outData[0]), .D(\u_outFIFO/n311 ), .Q(\u_outFIFO/n314 ) );
  INV3 U4346 ( .A(\u_cordic/mycordic/n513 ), .Q(n1459) );
  AOI221 U4347 ( .A(\u_cordic/mycordic/N338 ), .B(n772), .C(
        \u_cordic/mycordic/N370 ), .D(n1904), .Q(\u_cordic/mycordic/n513 ) );
  XNR21 U4348 ( .A(\u_cordic/mycordic/present_ANGLE_table[1][6] ), .B(
        \u_cordic/mycordic/sub_196/carry[6] ), .Q(\u_cordic/mycordic/N370 ) );
  XOR21 U4349 ( .A(\u_cordic/mycordic/present_ANGLE_table[1][6] ), .B(
        \u_cordic/mycordic/add_191/carry[6] ), .Q(\u_cordic/mycordic/N338 ) );
  INV3 U4350 ( .A(\u_cordic/mycordic/n512 ), .Q(n1460) );
  AOI221 U4351 ( .A(\u_cordic/mycordic/N339 ), .B(\u_cordic/mycordic/n336 ), 
        .C(\u_cordic/mycordic/N371 ), .D(n1904), .Q(\u_cordic/mycordic/n512 )
         );
  XNR21 U4352 ( .A(\u_cordic/mycordic/present_ANGLE_table[1][7] ), .B(
        \u_cordic/mycordic/sub_196/carry[7] ), .Q(\u_cordic/mycordic/N371 ) );
  XOR21 U4353 ( .A(\u_cordic/mycordic/present_ANGLE_table[1][7] ), .B(
        \u_cordic/mycordic/add_191/carry[7] ), .Q(\u_cordic/mycordic/N339 ) );
  INV3 U4354 ( .A(\u_cordic/mycordic/n497 ), .Q(n1552) );
  AOI221 U4355 ( .A(\u_cordic/mycordic/N402 ), .B(\u_cordic/mycordic/n332 ), 
        .C(\u_cordic/mycordic/N434 ), .D(n1908), .Q(\u_cordic/mycordic/n497 )
         );
  XNR21 U4356 ( .A(\u_cordic/mycordic/present_ANGLE_table[2][6] ), .B(
        \u_cordic/mycordic/sub_207/carry [6]), .Q(\u_cordic/mycordic/N434 ) );
  XOR21 U4357 ( .A(\u_cordic/mycordic/present_ANGLE_table[2][6] ), .B(
        \u_cordic/mycordic/add_202/carry [6]), .Q(\u_cordic/mycordic/N402 ) );
  INV3 U4358 ( .A(\u_cordic/mycordic/n496 ), .Q(n1553) );
  AOI221 U4359 ( .A(\u_cordic/mycordic/N403 ), .B(n778), .C(
        \u_cordic/mycordic/N435 ), .D(n1908), .Q(\u_cordic/mycordic/n496 ) );
  XNR21 U4360 ( .A(\u_cordic/mycordic/present_ANGLE_table[2][7] ), .B(
        \u_cordic/mycordic/sub_207/carry [7]), .Q(\u_cordic/mycordic/N435 ) );
  XOR21 U4361 ( .A(\u_cordic/mycordic/present_ANGLE_table[2][7] ), .B(
        \u_cordic/mycordic/add_202/carry [7]), .Q(\u_cordic/mycordic/N403 ) );
  INV3 U4362 ( .A(\u_cordic/mycordic/n495 ), .Q(n1554) );
  AOI221 U4363 ( .A(\u_cordic/mycordic/N404 ), .B(\u_cordic/mycordic/n332 ), 
        .C(\u_cordic/mycordic/N436 ), .D(n1908), .Q(\u_cordic/mycordic/n495 )
         );
  XNR21 U4364 ( .A(\u_cordic/mycordic/present_ANGLE_table[2][8] ), .B(
        \u_cordic/mycordic/sub_207/carry [8]), .Q(\u_cordic/mycordic/N436 ) );
  XOR21 U4365 ( .A(\u_cordic/mycordic/present_ANGLE_table[2][8] ), .B(
        \u_cordic/mycordic/add_202/carry [8]), .Q(\u_cordic/mycordic/N404 ) );
  INV3 U4366 ( .A(\u_cordic/mycordic/n482 ), .Q(n1526) );
  AOI221 U4367 ( .A(\u_cordic/mycordic/N461 ), .B(\u_cordic/mycordic/n363 ), 
        .C(\u_cordic/mycordic/N489 ), .D(n1907), .Q(\u_cordic/mycordic/n482 )
         );
  XNR21 U4368 ( .A(\u_cordic/mycordic/present_ANGLE_table[3][5] ), .B(
        \u_cordic/mycordic/sub_218/carry[5] ), .Q(\u_cordic/mycordic/N489 ) );
  XOR21 U4369 ( .A(\u_cordic/mycordic/present_ANGLE_table[3][5] ), .B(
        \u_cordic/mycordic/add_213/carry[5] ), .Q(\u_cordic/mycordic/N461 ) );
  INV3 U4370 ( .A(\u_cordic/mycordic/n481 ), .Q(n1527) );
  AOI221 U4371 ( .A(\u_cordic/mycordic/N462 ), .B(n777), .C(
        \u_cordic/mycordic/N490 ), .D(n1907), .Q(\u_cordic/mycordic/n481 ) );
  XNR21 U4372 ( .A(\u_cordic/mycordic/present_ANGLE_table[3][6] ), .B(
        \u_cordic/mycordic/sub_218/carry[6] ), .Q(\u_cordic/mycordic/N490 ) );
  XOR21 U4373 ( .A(\u_cordic/mycordic/present_ANGLE_table[3][6] ), .B(
        \u_cordic/mycordic/add_213/carry[6] ), .Q(\u_cordic/mycordic/N462 ) );
  INV3 U4374 ( .A(\u_cordic/mycordic/n480 ), .Q(n1528) );
  AOI221 U4375 ( .A(\u_cordic/mycordic/N463 ), .B(\u_cordic/mycordic/n363 ), 
        .C(\u_cordic/mycordic/N491 ), .D(n1907), .Q(\u_cordic/mycordic/n480 )
         );
  XNR21 U4376 ( .A(\u_cordic/mycordic/present_ANGLE_table[3][7] ), .B(
        \u_cordic/mycordic/sub_218/carry[7] ), .Q(\u_cordic/mycordic/N491 ) );
  XOR21 U4377 ( .A(\u_cordic/mycordic/present_ANGLE_table[3][7] ), .B(
        \u_cordic/mycordic/add_213/carry[7] ), .Q(\u_cordic/mycordic/N463 ) );
  INV3 U4378 ( .A(\u_cordic/mycordic/n467 ), .Q(n1501) );
  AOI221 U4379 ( .A(\u_cordic/mycordic/N505 ), .B(n776), .C(
        \u_cordic/mycordic/N522 ), .D(n1906), .Q(\u_cordic/mycordic/n467 ) );
  XNR21 U4380 ( .A(\u_cordic/mycordic/present_ANGLE_table[4][4] ), .B(
        \u_cordic/mycordic/sub_229/carry[4] ), .Q(\u_cordic/mycordic/N522 ) );
  XOR21 U4381 ( .A(\u_cordic/mycordic/present_ANGLE_table[4][4] ), .B(
        \u_cordic/mycordic/add_224/carry[4] ), .Q(\u_cordic/mycordic/N505 ) );
  INV3 U4382 ( .A(\u_cordic/mycordic/n466 ), .Q(n1502) );
  AOI221 U4383 ( .A(\u_cordic/mycordic/N506 ), .B(n776), .C(
        \u_cordic/mycordic/N523 ), .D(n1906), .Q(\u_cordic/mycordic/n466 ) );
  XNR21 U4384 ( .A(\u_cordic/mycordic/present_ANGLE_table[4][5] ), .B(
        \u_cordic/mycordic/sub_229/carry[5] ), .Q(\u_cordic/mycordic/N523 ) );
  XOR21 U4385 ( .A(\u_cordic/mycordic/present_ANGLE_table[4][5] ), .B(
        \u_cordic/mycordic/add_224/carry[5] ), .Q(\u_cordic/mycordic/N506 ) );
  INV3 U4386 ( .A(\u_cordic/mycordic/n465 ), .Q(n1503) );
  AOI221 U4387 ( .A(\u_cordic/mycordic/N507 ), .B(\u_cordic/mycordic/n456 ), 
        .C(\u_cordic/mycordic/N524 ), .D(n1906), .Q(\u_cordic/mycordic/n465 )
         );
  XNR21 U4388 ( .A(\u_cordic/mycordic/present_ANGLE_table[4][6] ), .B(
        \u_cordic/mycordic/sub_229/carry[6] ), .Q(\u_cordic/mycordic/N524 ) );
  XOR21 U4389 ( .A(\u_cordic/mycordic/present_ANGLE_table[4][6] ), .B(
        \u_cordic/mycordic/add_224/carry[6] ), .Q(\u_cordic/mycordic/N507 ) );
  INV3 U4390 ( .A(\u_cordic/mycordic/n464 ), .Q(n1504) );
  AOI221 U4391 ( .A(\u_cordic/mycordic/N508 ), .B(n776), .C(
        \u_cordic/mycordic/N525 ), .D(n1906), .Q(\u_cordic/mycordic/n464 ) );
  XNR21 U4392 ( .A(\u_cordic/mycordic/present_ANGLE_table[4][7] ), .B(
        \u_cordic/mycordic/sub_229/carry[7] ), .Q(\u_cordic/mycordic/N525 ) );
  XOR21 U4393 ( .A(\u_cordic/mycordic/present_ANGLE_table[4][7] ), .B(
        \u_cordic/mycordic/add_224/carry[7] ), .Q(\u_cordic/mycordic/N508 ) );
  INV3 U4394 ( .A(\u_cordic/mycordic/n515 ), .Q(n1457) );
  AOI221 U4395 ( .A(\u_cordic/mycordic/N336 ), .B(n772), .C(
        \u_cordic/mycordic/N368 ), .D(n1904), .Q(\u_cordic/mycordic/n515 ) );
  XOR21 U4396 ( .A(\u_cordic/mycordic/present_ANGLE_table[1][4] ), .B(
        \u_cordic/mycordic/sub_196/carry[4] ), .Q(\u_cordic/mycordic/N368 ) );
  XNR21 U4397 ( .A(\u_cordic/mycordic/present_ANGLE_table[1][4] ), .B(
        \u_cordic/mycordic/add_191/carry[4] ), .Q(\u_cordic/mycordic/N336 ) );
  INV3 U4398 ( .A(\u_decoder/fir_filter/n1037 ), .Q(n2637) );
  NAND22 U4399 ( .A(\u_decoder/fir_filter/I_data_mult_6_buff [0]), .B(n1156), 
        .Q(\u_decoder/fir_filter/n1037 ) );
  INV3 U4400 ( .A(\u_decoder/fir_filter/n805 ), .Q(n2518) );
  NAND22 U4401 ( .A(\u_decoder/fir_filter/Q_data_mult_2_buff [0]), .B(n1154), 
        .Q(\u_decoder/fir_filter/n805 ) );
  INV3 U4402 ( .A(\u_decoder/fir_filter/n740 ), .Q(n2517) );
  NAND22 U4403 ( .A(\u_decoder/fir_filter/Q_data_mult_6_buff [0]), .B(n1156), 
        .Q(\u_decoder/fir_filter/n740 ) );
  INV3 U4404 ( .A(\u_cordic/mycordic/n411 ), .Q(n1880) );
  NAND22 U4405 ( .A(\u_cordic/mycordic/next_ANGLE_table[6][3] ), .B(n1214), 
        .Q(\u_cordic/mycordic/n411 ) );
  INV3 U4406 ( .A(\u_cordic/mycordic/n410 ), .Q(n1879) );
  NAND22 U4407 ( .A(\u_cordic/mycordic/next_ANGLE_table[6][4] ), .B(n1214), 
        .Q(\u_cordic/mycordic/n410 ) );
  INV3 U4408 ( .A(\u_cordic/mycordic/n409 ), .Q(n1878) );
  NAND22 U4409 ( .A(\u_cordic/mycordic/next_ANGLE_table[6][5] ), .B(n1215), 
        .Q(\u_cordic/mycordic/n409 ) );
  INV3 U4410 ( .A(\u_cordic/mycordic/n408 ), .Q(n1877) );
  NAND22 U4411 ( .A(\u_cordic/mycordic/next_ANGLE_table[6][6] ), .B(n1214), 
        .Q(\u_cordic/mycordic/n408 ) );
  NAND31 U4412 ( .A(n756), .B(\u_decoder/iq_demod/cossin_dig/n23 ), .C(n1217), 
        .Q(\u_decoder/iq_demod/cossin_dig/n44 ) );
  INV3 U4413 ( .A(\u_cordic/mycordic/n554 ), .Q(n1908) );
  NAND22 U4414 ( .A(\u_cordic/mycordic/present_Q_table[3][7] ), .B(n1212), .Q(
        \u_cordic/mycordic/n554 ) );
  NAND22 U4415 ( .A(\u_cordic/mycordic/present_Q_table[2][7] ), .B(n1213), .Q(
        \u_cordic/mycordic/n520 ) );
  NOR40 U4416 ( .A(\u_cordic/mycordic/present_Q_table[0][3] ), .B(
        \u_cordic/mycordic/present_Q_table[0][4] ), .C(n2658), .D(n769), .Q(
        \u_cordic/mycordic/N212 ) );
  INV3 U4417 ( .A(\u_cordic/mycordic/n435 ), .Q(n2658) );
  NOR31 U4418 ( .A(\u_cordic/mycordic/present_Q_table[0][5] ), .B(
        \u_cordic/mycordic/present_Q_table[0][7] ), .C(
        \u_cordic/mycordic/present_Q_table[0][6] ), .Q(
        \u_cordic/mycordic/n435 ) );
  NAND22 U4419 ( .A(sig_DEMUX_outDEMUX2[2]), .B(n2133), .Q(\u_mux8/n3 ) );
  AOI221 U4420 ( .A(\sig_MUX_inMUX8[0] ), .B(n2133), .C(in_MUX_inSEL6[0]), .D(
        sig_DEMUX_outDEMUX2[2]), .Q(\u_mux8/n4 ) );
  NOR31 U4421 ( .A(n3118), .B(in_DEMUX_inSEL2[2]), .C(n2129), .Q(
        sig_DEMUX_outDEMUX2[2]) );
  AOI211 U4422 ( .A(\u_decoder/iq_demod/cossin_dig/val_counter [1]), .B(
        \u_decoder/iq_demod/cossin_dig/N55 ), .C(
        \u_decoder/iq_demod/cossin_dig/val_counter [2]), .Q(
        \u_decoder/iq_demod/cossin_dig/n37 ) );
  NAND22 U4423 ( .A(\u_outFIFO/n253 ), .B(\u_outFIFO/n254 ), .Q(
        \u_outFIFO/n1155 ) );
  NAND22 U4424 ( .A(\u_cordic/mycordic/present_I_table[0][7] ), .B(n1213), .Q(
        \u_cordic/mycordic/n391 ) );
  NAND22 U4425 ( .A(\u_cordic/n11 ), .B(\u_cordic/n9 ), .Q(\u_cordic/n19 ) );
  NOR21 U4426 ( .A(\u_decoder/iq_demod/cossin_dig/n23 ), .B(n756), .Q(
        \u_decoder/iq_demod/cossin_dig/n26 ) );
  INV3 U4427 ( .A(\u_cordic/mycordic/n537 ), .Q(n1905) );
  NAND22 U4428 ( .A(\u_cordic/mycordic/present_Q_table[1][7] ), .B(n1212), .Q(
        \u_cordic/mycordic/n537 ) );
  INV3 U4429 ( .A(\u_cordic/mycordic/n454 ), .Q(n1903) );
  NAND22 U4430 ( .A(\u_cordic/mycordic/present_Q_table[6][7] ), .B(n1212), .Q(
        \u_cordic/mycordic/n454 ) );
  NOR31 U4431 ( .A(\u_outFIFO/n256 ), .B(\u_outFIFO/currentState [0]), .C(
        \u_outFIFO/n1155 ), .Q(\u_outFIFO/n1148 ) );
  NOR31 U4432 ( .A(\u_inFIFO/n177 ), .B(\u_inFIFO/n176 ), .C(\u_inFIFO/n568 ), 
        .Q(\u_inFIFO/n560 ) );
  NAND31 U4433 ( .A(\u_inFIFO/currentState [0]), .B(\u_inFIFO/n176 ), .C(n2142), .Q(\u_inFIFO/n563 ) );
  NOR21 U4434 ( .A(\u_cordic/present_state [1]), .B(
        \u_cordic/present_state [0]), .Q(\u_cordic/n15 ) );
  NOR40 U4435 ( .A(n2690), .B(n3055), .C(\u_cdr/phd1/cnt_phd/cnt [1]), .D(
        n1239), .Q(\u_cdr/phd1/cnt_phd/N84 ) );
  INV3 U4436 ( .A(n3068), .Q(n2690) );
  NOR40 U4437 ( .A(\u_cdr/phd1/cnt_phd/cnt [2]), .B(
        \u_cdr/phd1/cnt_phd/cnt [3]), .C(\u_cdr/phd1/cnt_phd/cnt [4]), .D(
        \u_cdr/phd1/cnt_phd/cnt [5]), .Q(n3068) );
  INV3 U4438 ( .A(\u_cordic/mycordic/n539 ), .Q(n1906) );
  NAND22 U4439 ( .A(\u_cordic/mycordic/present_Q_table[5][7] ), .B(n1212), .Q(
        \u_cordic/mycordic/n539 ) );
  OAI2111 U4440 ( .A(\u_cordic/mycordic/present_Q_table[0][7] ), .B(
        \u_cordic/mycordic/n391 ), .C(\u_cordic/mycordic/n432 ), .D(n1426), 
        .Q(\u_cordic/mycordic/N211 ) );
  NAND22 U4441 ( .A(\u_cordic/mycordic/present_Q_table[0][7] ), .B(
        \u_cordic/mycordic/n354 ), .Q(\u_cordic/mycordic/n432 ) );
  INV3 U4442 ( .A(\u_cordic/mycordic/N212 ), .Q(n1426) );
  NAND22 U4443 ( .A(\u_decoder/iq_demod/cossin_dig/counter [1]), .B(
        \u_decoder/iq_demod/cossin_dig/counter [0]), .Q(
        \u_decoder/iq_demod/cossin_dig/n43 ) );
  NOR31 U4444 ( .A(\u_cdr/cnt_in [1]), .B(\u_cdr/cnt_in [3]), .C(
        \u_cdr/cnt_in [0]), .Q(\u_cdr/n43 ) );
  NOR31 U4445 ( .A(\u_outFIFO/n257 ), .B(\u_outFIFO/n256 ), .C(
        \u_outFIFO/n1155 ), .Q(\u_outFIFO/n1147 ) );
  NOR21 U4446 ( .A(\u_decoder/fir_filter/n410 ), .B(
        \u_decoder/fir_filter/state [1]), .Q(\u_decoder/fir_filter/n1151 ) );
  INV3 U4447 ( .A(\u_cordic/n26 ), .Q(n2117) );
  AOI221 U4448 ( .A(sig_MUX_outMUX7[3]), .B(\u_cordic/n18 ), .C(
        \u_cordic/Q [3]), .D(\u_cordic/n19 ), .Q(\u_cordic/n26 ) );
  NAND22 U4449 ( .A(sig_DEMUX_outDEMUX18[7]), .B(n2133), .Q(n3110) );
  INV3 U4450 ( .A(\u_cordic/n25 ), .Q(n2119) );
  AOI221 U4451 ( .A(sig_MUX_outMUX7[2]), .B(\u_cordic/n18 ), .C(
        \u_cordic/Q [2]), .D(\u_cordic/n19 ), .Q(\u_cordic/n25 ) );
  NAND22 U4452 ( .A(sig_DEMUX_outDEMUX18[6]), .B(n2133), .Q(n3108) );
  INV3 U4453 ( .A(\u_cordic/n24 ), .Q(n2121) );
  AOI221 U4454 ( .A(sig_MUX_outMUX7[1]), .B(\u_cordic/n18 ), .C(
        \u_cordic/Q [1]), .D(\u_cordic/n19 ), .Q(\u_cordic/n24 ) );
  NAND22 U4455 ( .A(sig_DEMUX_outDEMUX18[5]), .B(n2133), .Q(n3106) );
  INV3 U4456 ( .A(\u_cordic/n23 ), .Q(n2123) );
  AOI221 U4457 ( .A(sig_MUX_outMUX7[0]), .B(\u_cordic/n18 ), .C(
        \u_cordic/Q [0]), .D(\u_cordic/n19 ), .Q(\u_cordic/n23 ) );
  NAND22 U4458 ( .A(sig_DEMUX_outDEMUX18[4]), .B(n2133), .Q(n3104) );
  INV3 U4459 ( .A(\u_cordic/n22 ), .Q(n2109) );
  AOI221 U4460 ( .A(sig_MUX_outMUX6[3]), .B(\u_cordic/n18 ), .C(
        \u_cordic/I [3]), .D(\u_cordic/n19 ), .Q(\u_cordic/n22 ) );
  NAND22 U4461 ( .A(sig_DEMUX_outDEMUX17[7]), .B(n2133), .Q(n3102) );
  INV3 U4462 ( .A(\u_cordic/n21 ), .Q(n2111) );
  AOI221 U4463 ( .A(sig_MUX_outMUX6[2]), .B(\u_cordic/n18 ), .C(
        \u_cordic/I [2]), .D(\u_cordic/n19 ), .Q(\u_cordic/n21 ) );
  NAND22 U4464 ( .A(sig_DEMUX_outDEMUX17[6]), .B(n2133), .Q(n3100) );
  INV3 U4465 ( .A(\u_cordic/n20 ), .Q(n2113) );
  AOI221 U4466 ( .A(sig_MUX_outMUX6[1]), .B(\u_cordic/n18 ), .C(
        \u_cordic/I [1]), .D(\u_cordic/n19 ), .Q(\u_cordic/n20 ) );
  NAND22 U4467 ( .A(sig_DEMUX_outDEMUX17[5]), .B(n2133), .Q(n3098) );
  INV3 U4468 ( .A(\u_cordic/n17 ), .Q(n2115) );
  AOI221 U4469 ( .A(sig_MUX_outMUX6[0]), .B(\u_cordic/n18 ), .C(
        \u_cordic/I [0]), .D(\u_cordic/n19 ), .Q(\u_cordic/n17 ) );
  NAND22 U4470 ( .A(sig_DEMUX_outDEMUX17[4]), .B(n2133), .Q(n3096) );
  INV3 U4471 ( .A(\u_cordic/mycordic/n547 ), .Q(n1513) );
  AOI221 U4472 ( .A(\u_cordic/mycordic/N448 ), .B(n777), .C(
        \u_cordic/mycordic/N476 ), .D(n1907), .Q(\u_cordic/mycordic/n547 ) );
  XOR21 U4473 ( .A(\u_cordic/mycordic/present_Q_table[4][0] ), .B(
        \u_cordic/mycordic/present_I_table[4][3] ), .Q(
        \u_cordic/mycordic/N476 ) );
  XNR21 U4474 ( .A(\u_cordic/mycordic/present_Q_table[4][0] ), .B(n163), .Q(
        \u_cordic/mycordic/N448 ) );
  INV3 U4475 ( .A(\u_cordic/mycordic/n487 ), .Q(n1521) );
  AOI221 U4476 ( .A(n295), .B(n777), .C(n295), .D(n1907), .Q(
        \u_cordic/mycordic/n487 ) );
  INV3 U4477 ( .A(\u_cordic/mycordic/n486 ), .Q(n1522) );
  AOI221 U4478 ( .A(\u_cordic/mycordic/N457 ), .B(\u_cordic/mycordic/n363 ), 
        .C(\u_cordic/mycordic/N485 ), .D(n1907), .Q(\u_cordic/mycordic/n486 )
         );
  XOR21 U4479 ( .A(\u_cordic/mycordic/present_ANGLE_table[3][1] ), .B(
        \u_cordic/mycordic/present_ANGLE_table[3][0] ), .Q(
        \u_cordic/mycordic/N485 ) );
  XNR21 U4480 ( .A(\u_cordic/mycordic/present_ANGLE_table[3][1] ), .B(
        \u_cordic/mycordic/present_ANGLE_table[3][0] ), .Q(
        \u_cordic/mycordic/N457 ) );
  INV3 U4481 ( .A(\u_cordic/mycordic/n453 ), .Q(n1437) );
  AOI221 U4482 ( .A(\u_cordic/mycordic/N550 ), .B(n770), .C(
        \u_cordic/mycordic/N550 ), .D(n1903), .Q(\u_cordic/mycordic/n453 ) );
  INV3 U4483 ( .A(\u_cordic/mycordic/n452 ), .Q(n1438) );
  AOI221 U4484 ( .A(n296), .B(n771), .C(n296), .D(n1903), .Q(
        \u_cordic/mycordic/n452 ) );
  INV3 U4485 ( .A(\u_cordic/mycordic/n451 ), .Q(n1439) );
  AOI221 U4486 ( .A(\u_cordic/mycordic/N536 ), .B(n770), .C(
        \u_cordic/mycordic/N552 ), .D(n1903), .Q(\u_cordic/mycordic/n451 ) );
  XNR21 U4487 ( .A(\u_cordic/mycordic/present_ANGLE_table[5][2] ), .B(
        \u_cordic/mycordic/present_ANGLE_table[5][1] ), .Q(
        \u_cordic/mycordic/N552 ) );
  XOR21 U4488 ( .A(\u_cordic/mycordic/present_ANGLE_table[5][2] ), .B(
        \u_cordic/mycordic/present_ANGLE_table[5][1] ), .Q(
        \u_cordic/mycordic/N536 ) );
  INV3 U4489 ( .A(\u_cordic/mycordic/n450 ), .Q(n1440) );
  AOI221 U4490 ( .A(\u_cordic/mycordic/N537 ), .B(n771), .C(
        \u_cordic/mycordic/N553 ), .D(n1903), .Q(\u_cordic/mycordic/n450 ) );
  XNR21 U4491 ( .A(\u_cordic/mycordic/present_ANGLE_table[5][3] ), .B(
        \u_cordic/mycordic/sub_236/carry [3]), .Q(\u_cordic/mycordic/N553 ) );
  XOR21 U4492 ( .A(\u_cordic/mycordic/present_ANGLE_table[5][3] ), .B(
        \u_cordic/mycordic/add_233/carry [3]), .Q(\u_cordic/mycordic/N537 ) );
  INV3 U4493 ( .A(\u_cordic/mycordic/n355 ), .Q(n1435) );
  AOI221 U4494 ( .A(n1901), .B(\u_cordic/mycordic/N246 ), .C(
        \u_cordic/mycordic/n354 ), .D(
        \u_cordic/mycordic/present_Q_table[0][6] ), .Q(
        \u_cordic/mycordic/n355 ) );
  XOR21 U4495 ( .A(\u_cordic/mycordic/sub_add_151_b0/carry [6]), .B(n53), .Q(
        \u_cordic/mycordic/N246 ) );
  INV3 U4496 ( .A(\u_inFIFO/os1/dff1/n2 ), .Q(n1848) );
  NAND22 U4497 ( .A(n1218), .B(n2100), .Q(\u_inFIFO/os1/dff1/n2 ) );
  INV3 U4498 ( .A(\u_mux3/n3 ), .Q(n2100) );
  AOI221 U4499 ( .A(\sig_MUX_inMUX3[0] ), .B(n2131), .C(in_MUX_inSEL3), .D(
        sig_DEMUX_outDEMUX1[2]), .Q(\u_mux3/n3 ) );
  INV3 U4500 ( .A(\u_cordic/mycordic/n393 ), .Q(n1430) );
  AOI221 U4501 ( .A(\u_cordic/mycordic/present_I_table[0][5] ), .B(
        \u_cordic/mycordic/n354 ), .C(\u_cordic/mycordic/N237 ), .D(n1901), 
        .Q(\u_cordic/mycordic/n393 ) );
  XOR21 U4502 ( .A(\u_cordic/mycordic/sub_add_150_b0/carry [5]), .B(n56), .Q(
        \u_cordic/mycordic/N237 ) );
  INV3 U4503 ( .A(\u_cordic/mycordic/n392 ), .Q(n1431) );
  AOI221 U4504 ( .A(\u_cordic/mycordic/present_I_table[0][6] ), .B(
        \u_cordic/mycordic/n354 ), .C(\u_cordic/mycordic/N238 ), .D(n1901), 
        .Q(\u_cordic/mycordic/n392 ) );
  XOR21 U4505 ( .A(\u_cordic/mycordic/sub_add_150_b0/carry [6]), .B(n57), .Q(
        \u_cordic/mycordic/N238 ) );
  INV3 U4506 ( .A(\u_decoder/iq_demod/cossin_dig/n39 ), .Q(n1845) );
  NAND22 U4507 ( .A(\u_cdr/cnt_d [1]), .B(\u_cdr/cnt_d [0]), .Q(
        \u_cdr/dec1/cnt_dec/n24 ) );
  NAND22 U4508 ( .A(\u_cdr/cnt_d [1]), .B(\u_cdr/cnt_d [0]), .Q(n3064) );
  NAND22 U4509 ( .A(\u_cdr/cnt_d [1]), .B(\u_cdr/cnt_d [0]), .Q(
        \u_cdr/div1/cnt_div/n41 ) );
  XNR21 U4510 ( .A(\u_inFIFO/n197 ), .B(\u_inFIFO/n198 ), .Q(\u_inFIFO/n530 )
         );
  NOR40 U4511 ( .A(n1239), .B(\u_inFIFO/n197 ), .C(\u_inFIFO/n198 ), .D(
        \u_inFIFO/n531 ), .Q(\u_inFIFO/N196 ) );
  AOI221 U4512 ( .A(sig_decod_outQ[3]), .B(n2133), .C(in_MUX_inSEL6[0]), .D(
        sig_coder_outSinQMasked[3]), .Q(n3111) );
  AOI221 U4513 ( .A(sig_decod_outQ[2]), .B(n2133), .C(in_MUX_inSEL6[0]), .D(
        sig_coder_outSinQMasked[2]), .Q(n3109) );
  AOI221 U4514 ( .A(sig_decod_outQ[1]), .B(n2133), .C(in_MUX_inSEL6[0]), .D(
        sig_coder_outSinQMasked[1]), .Q(n3107) );
  AOI221 U4515 ( .A(sig_decod_outQ[0]), .B(n2133), .C(in_MUX_inSEL6[0]), .D(
        sig_coder_outSinQMasked[0]), .Q(n3105) );
  AOI221 U4516 ( .A(sig_decod_outI[3]), .B(n2133), .C(in_MUX_inSEL6[0]), .D(
        sig_coder_outSinIMasked[3]), .Q(n3103) );
  AOI221 U4517 ( .A(sig_decod_outI[2]), .B(n2133), .C(in_MUX_inSEL6[0]), .D(
        sig_coder_outSinIMasked[2]), .Q(n3101) );
  AOI221 U4518 ( .A(sig_decod_outI[1]), .B(n2133), .C(in_MUX_inSEL6[0]), .D(
        sig_coder_outSinIMasked[1]), .Q(n3099) );
  AOI221 U4519 ( .A(sig_decod_outI[0]), .B(n2133), .C(in_MUX_inSEL6[0]), .D(
        sig_coder_outSinIMasked[0]), .Q(n3097) );
  NOR21 U4520 ( .A(\u_inFIFO/n176 ), .B(\u_inFIFO/currentState [0]), .Q(
        \u_inFIFO/n212 ) );
  BUF2 U4521 ( .A(\u_outFIFO/N44 ), .Q(n761) );
  NAND22 U4522 ( .A(\u_outFIFO/sigEnableCounter ), .B(n1212), .Q(
        \u_outFIFO/n1129 ) );
  NAND22 U4523 ( .A(\u_inFIFO/sigEnableCounter ), .B(n1217), .Q(
        \u_inFIFO/n553 ) );
  NOR21 U4524 ( .A(n1236), .B(\u_cordic/mycordic/present_Q_table[3][7] ), .Q(
        \u_cordic/mycordic/n332 ) );
  NAND22 U4525 ( .A(\u_inFIFO/n154 ), .B(\u_inFIFO/n173 ), .Q(\u_inFIFO/n568 )
         );
  OAI311 U4526 ( .A(\u_decoder/iq_demod/cossin_dig/n43 ), .B(
        \u_decoder/iq_demod/cossin_dig/counter [2]), .C(
        \u_decoder/iq_demod/cossin_dig/n44 ), .D(
        \u_decoder/iq_demod/cossin_dig/n46 ), .Q(
        \u_decoder/iq_demod/cossin_dig/N22 ) );
  NOR21 U4527 ( .A(\u_decoder/iq_demod/cossin_dig/counter [1]), .B(
        \u_decoder/iq_demod/cossin_dig/n44 ), .Q(
        \u_decoder/iq_demod/cossin_dig/n47 ) );
  NAND22 U4528 ( .A(\u_outFIFO/n257 ), .B(\u_outFIFO/n256 ), .Q(
        \u_outFIFO/n1144 ) );
  NOR21 U4529 ( .A(n1239), .B(\u_cordic/mycordic/present_Q_table[2][7] ), .Q(
        \u_cordic/mycordic/n336 ) );
  NAND22 U4530 ( .A(\u_decoder/iq_demod/sin_out [0]), .B(n756), .Q(
        \u_decoder/iq_demod/cossin_dig/n32 ) );
  BUF2 U4531 ( .A(\u_decoder/iq_demod/cossin_dig/state[0] ), .Q(n756) );
  INV3 U4532 ( .A(\u_cordic/mycordic/n449 ), .Q(n1441) );
  AOI221 U4533 ( .A(\u_cordic/mycordic/N538 ), .B(n770), .C(
        \u_cordic/mycordic/N554 ), .D(n1903), .Q(\u_cordic/mycordic/n449 ) );
  XNR21 U4534 ( .A(\u_cordic/mycordic/present_ANGLE_table[5][4] ), .B(
        \u_cordic/mycordic/sub_236/carry [4]), .Q(\u_cordic/mycordic/N554 ) );
  XOR21 U4535 ( .A(\u_cordic/mycordic/present_ANGLE_table[5][4] ), .B(
        \u_cordic/mycordic/add_233/carry [4]), .Q(\u_cordic/mycordic/N538 ) );
  BUF2 U4536 ( .A(\u_cordic/mycordic/n108 ), .Q(n758) );
  NAND31 U4537 ( .A(\u_cordic/dir ), .B(\u_cordic/n15 ), .C(
        \u_cordic/present_state [2]), .Q(\u_cordic/n16 ) );
  NOR21 U4538 ( .A(\u_cdr/phd1/w_en_f ), .B(\u_cdr/phd1/w_en_d ), .Q(
        \u_cdr/phd1/n15 ) );
  NOR21 U4539 ( .A(n1232), .B(\u_cordic/mycordic/present_Q_table[1][7] ), .Q(
        \u_cordic/mycordic/n345 ) );
  NAND22 U4540 ( .A(\u_coder/n150 ), .B(\u_coder/n101 ), .Q(\u_coder/n145 ) );
  NOR21 U4541 ( .A(\u_decoder/iq_demod/cossin_dig/n44 ), .B(
        \u_decoder/iq_demod/cossin_dig/counter [0]), .Q(
        \u_decoder/iq_demod/cossin_dig/N20 ) );
  AOI311 U4542 ( .A(n2221), .B(\u_outFIFO/n253 ), .C(
        \u_outFIFO/sig_fsm_start_R ), .D(\u_outFIFO/n1148 ), .Q(
        \u_outFIFO/n1157 ) );
  INV3 U4543 ( .A(\u_outFIFO/n1144 ), .Q(n2221) );
  AOI2111 U4544 ( .A(\u_cordic/n29 ), .B(\u_cordic/n30 ), .C(n1240), .D(
        \u_cordic/present_state [2]), .Q(\u_cordic/N15 ) );
  NAND22 U4545 ( .A(\u_cordic/present_state [1]), .B(\u_cordic/n11 ), .Q(
        \u_cordic/n29 ) );
  NAND31 U4546 ( .A(\u_cordic/present_state [0]), .B(\u_cordic/n10 ), .C(
        sig_MUX_outMUX8), .Q(\u_cordic/n30 ) );
  AOI311 U4547 ( .A(\u_inFIFO/n567 ), .B(\u_inFIFO/n154 ), .C(\u_inFIFO/n557 ), 
        .D(\u_inFIFO/n560 ), .Q(\u_inFIFO/n565 ) );
  XOR21 U4548 ( .A(\u_inFIFO/sig_fsm_start_R ), .B(\u_inFIFO/sig_fsm_start_W ), 
        .Q(\u_inFIFO/n567 ) );
  NOR21 U4549 ( .A(\u_inFIFO/os2/sigQout2 ), .B(n317), .Q(
        \u_inFIFO/sig_fsm_start_W ) );
  NOR21 U4550 ( .A(\u_outFIFO/os1/sigQout2 ), .B(n284), .Q(
        \u_outFIFO/sig_fsm_start_R ) );
  NOR21 U4551 ( .A(\u_inFIFO/os1/sigQout2 ), .B(n318), .Q(
        \u_inFIFO/sig_fsm_start_R ) );
  NAND22 U4552 ( .A(\u_decoder/iq_demod/state [1]), .B(
        \u_decoder/iq_demod/n30 ), .Q(\u_decoder/iq_demod/n59 ) );
  NAND22 U4553 ( .A(\u_decoder/iq_demod/cossin_dig/n26 ), .B(n2686), .Q(
        \u_decoder/iq_demod/cossin_dig/n27 ) );
  INV3 U4554 ( .A(\u_decoder/iq_demod/cossin_dig/n55 ), .Q(n2686) );
  NOR21 U4555 ( .A(\u_inFIFO/currentState [0]), .B(\u_inFIFO/currentState [1]), 
        .Q(\u_inFIFO/n557 ) );
  NOR21 U4556 ( .A(n1237), .B(\u_cordic/mycordic/present_Q_table[6][7] ), .Q(
        \u_cordic/mycordic/n438 ) );
  AOI211 U4557 ( .A(\u_decoder/iq_demod/cossin_dig/n10 ), .B(
        \u_decoder/iq_demod/cossin_dig/n43 ), .C(
        \u_decoder/iq_demod/cossin_dig/n44 ), .Q(
        \u_decoder/iq_demod/cossin_dig/N42 ) );
  AOI211 U4558 ( .A(\u_cordic/n19 ), .B(\u_cordic/n31 ), .C(n1241), .Q(
        \u_cordic/N14 ) );
  INV3 U4559 ( .A(sig_MUX_outMUX8), .Q(n2107) );
  AOI211 U4560 ( .A(\u_cordic/n27 ), .B(\u_cordic/n28 ), .C(n1241), .Q(
        \u_cordic/N16 ) );
  NAND31 U4561 ( .A(\u_cordic/present_state [0]), .B(\u_cordic/n9 ), .C(
        \u_cordic/present_state [1]), .Q(\u_cordic/n28 ) );
  NAND22 U4562 ( .A(\u_cordic/present_state [2]), .B(\u_cordic/n15 ), .Q(
        \u_cordic/n27 ) );
  AOI211 U4563 ( .A(\u_decoder/iq_demod/cossin_dig/state[0] ), .B(
        \u_decoder/iq_demod/cossin_dig/n45 ), .C(n1241), .Q(
        \u_decoder/iq_demod/cossin_dig/N41 ) );
  NAND31 U4564 ( .A(\u_decoder/iq_demod/cossin_dig/n10 ), .B(
        \u_decoder/iq_demod/cossin_dig/n23 ), .C(
        \u_decoder/iq_demod/cossin_dig/n43 ), .Q(
        \u_decoder/iq_demod/cossin_dig/n45 ) );
  AOI211 U4565 ( .A(n320), .B(n1336), .C(n1235), .Q(n1833) );
  INV3 U4566 ( .A(\u_cordic/mycordic/n456 ), .Q(n775) );
  NOR21 U4567 ( .A(n1236), .B(\u_cordic/mycordic/present_Q_table[5][7] ), .Q(
        \u_cordic/mycordic/n456 ) );
  NOR31 U4568 ( .A(n294), .B(\u_decoder/fir_filter/state [1]), .C(n1239), .Q(
        \u_decoder/fir_filter/N12 ) );
  XOR21 U4569 ( .A(\u_cordic/mycordic/present_ANGLE_table[6][3] ), .B(
        \u_cordic/mycordic/present_ANGLE_table[6][4] ), .Q(
        \u_cordic/mycordic/N619 ) );
  INV3 U4570 ( .A(n3052), .Q(n1830) );
  NAND22 U4571 ( .A(n1218), .B(n2687), .Q(n3052) );
  INV3 U4572 ( .A(\u_cdr/phd1/n13 ), .Q(n2687) );
  AOI221 U4573 ( .A(\u_cdr/phd1/w_en_f ), .B(\u_cdr/phd1/w_s1 ), .C(n300), .D(
        \u_cdr/phd1/w_s2 ), .Q(\u_cdr/phd1/n13 ) );
  NOR21 U4574 ( .A(\u_outFIFO/os2/sigQout2 ), .B(n285), .Q(
        \u_outFIFO/sig_fsm_start_W ) );
  BUF2 U4575 ( .A(\u_decoder/iq_demod/n42 ), .Q(n779) );
  NOR21 U4576 ( .A(\u_decoder/iq_demod/n30 ), .B(\u_decoder/iq_demod/state [1]), .Q(\u_decoder/iq_demod/n42 ) );
  INV3 U4577 ( .A(\u_cordic/mycordic/n354 ), .Q(n769) );
  NOR21 U4578 ( .A(n1238), .B(\u_cordic/mycordic/present_I_table[0][7] ), .Q(
        \u_cordic/mycordic/n354 ) );
  NOR21 U4579 ( .A(\u_coder/c [6]), .B(\u_coder/c [5]), .Q(\u_coder/n322 ) );
  NOR21 U4580 ( .A(\u_decoder/iq_demod/cossin_dig/n48 ), .B(
        \u_decoder/iq_demod/cossin_dig/n44 ), .Q(
        \u_decoder/iq_demod/cossin_dig/N21 ) );
  XNR21 U4581 ( .A(\u_decoder/iq_demod/cossin_dig/counter [1]), .B(
        \u_decoder/iq_demod/cossin_dig/counter [0]), .Q(
        \u_decoder/iq_demod/cossin_dig/n48 ) );
  NOR21 U4582 ( .A(\u_cordic/mycordic/n391 ), .B(n51), .Q(
        \u_cordic/mycordic/N44 ) );
  NAND22 U4583 ( .A(\u_decoder/iq_demod/cossin_dig/n27 ), .B(
        \u_decoder/iq_demod/cossin_dig/n29 ), .Q(
        \u_decoder/iq_demod/cossin_dig/n50 ) );
  NAND22 U4584 ( .A(\u_decoder/iq_demod/cos_out [2]), .B(n756), .Q(
        \u_decoder/iq_demod/cossin_dig/n29 ) );
  NAND22 U4585 ( .A(\u_decoder/iq_demod/cossin_dig/n27 ), .B(
        \u_decoder/iq_demod/cossin_dig/n28 ), .Q(
        \u_decoder/iq_demod/cossin_dig/n49 ) );
  NAND22 U4586 ( .A(\u_decoder/iq_demod/cos_out [1]), .B(n756), .Q(
        \u_decoder/iq_demod/cossin_dig/n28 ) );
  INV3 U4587 ( .A(n3054), .Q(n1832) );
  NAND22 U4588 ( .A(n1219), .B(n2688), .Q(n3054) );
  INV3 U4589 ( .A(\u_cdr/phd1/n11 ), .Q(n2688) );
  AOI221 U4590 ( .A(\u_cdr/phd1/w_en_f ), .B(\u_cdr/phd1/w_s3 ), .C(n300), .D(
        \u_cdr/phd1/w_s4 ), .Q(\u_cdr/phd1/n11 ) );
  INV3 U4591 ( .A(\u_inFIFO/n566 ), .Q(n1829) );
  INV3 U4592 ( .A(\u_outFIFO/n1158 ), .Q(n1913) );
  NAND22 U4593 ( .A(\u_cdr/n33 ), .B(\u_cdr/n17 ), .Q(\u_cdr/n32 ) );
  INV3 U4594 ( .A(\u_cdr/n34 ), .Q(n1805) );
  INV3 U4595 ( .A(\u_cdr/n29 ), .Q(n1914) );
  NAND22 U4596 ( .A(n2106), .B(n1212), .Q(\u_cdr/n29 ) );
  INV3 U4597 ( .A(n3115), .Q(n2106) );
  AOI221 U4598 ( .A(\sig_MUX_inMUX14[0] ), .B(n2136), .C(in_MUX_inSEL11), .D(
        sig_DEMUX_outDEMUX2[3]), .Q(n3115) );
  XNR21 U4599 ( .A(\u_cordic/mycordic/present_ANGLE_table[6][2] ), .B(
        \u_cordic/mycordic/present_ANGLE_table[6][3] ), .Q(n393) );
  INV3 U4600 ( .A(\u_cdr/dec1/n24 ), .Q(n1849) );
  OAI2111 U4601 ( .A(\u_cdr/cnt_d [0]), .B(\u_cdr/cnt_d [1]), .C(n1220), .D(
        \u_cdr/dec1/n25 ), .Q(\u_cdr/dec1/n24 ) );
  INV3 U4602 ( .A(\u_decoder/iq_demod/cossin_dig/n25 ), .Q(n2680) );
  AOI221 U4603 ( .A(\u_decoder/iq_demod/cossin_dig/n26 ), .B(
        \u_decoder/iq_demod/cossin_dig/N55 ), .C(n756), .D(
        \u_decoder/iq_demod/cos_out [0]), .Q(
        \u_decoder/iq_demod/cossin_dig/n25 ) );
  INV3 U4604 ( .A(\u_outFIFO/N128 ), .Q(n2236) );
  INV3 U4605 ( .A(\u_outFIFO/N129 ), .Q(n2235) );
  INV3 U4606 ( .A(\u_cordic/mycordic/n433 ), .Q(n1427) );
  AOI211 U4607 ( .A(n1220), .B(\u_cordic/mycordic/present_Q_table[0][7] ), .C(
        \u_cordic/mycordic/N212 ), .Q(\u_cordic/mycordic/n433 ) );
  INV3 U4608 ( .A(\u_cordic/mycordic/n358 ), .Q(n1432) );
  AOI221 U4609 ( .A(n1901), .B(\u_cordic/mycordic/present_Q_table[0][3] ), .C(
        \u_cordic/mycordic/n354 ), .D(
        \u_cordic/mycordic/present_Q_table[0][3] ), .Q(
        \u_cordic/mycordic/n358 ) );
  INV3 U4610 ( .A(\u_decoder/iq_demod/cossin_dig/n30 ), .Q(n2681) );
  AOI221 U4611 ( .A(\u_decoder/iq_demod/cossin_dig/N52 ), .B(
        \u_decoder/iq_demod/cossin_dig/n26 ), .C(
        \u_decoder/iq_demod/cos_out [3]), .D(n756), .Q(
        \u_decoder/iq_demod/cossin_dig/n30 ) );
  INV3 U4612 ( .A(\u_cordic/mycordic/n395 ), .Q(n1428) );
  AOI221 U4613 ( .A(\u_cordic/mycordic/present_I_table[0][3] ), .B(
        \u_cordic/mycordic/n354 ), .C(
        \u_cordic/mycordic/present_I_table[0][3] ), .D(n1901), .Q(
        \u_cordic/mycordic/n395 ) );
  INV3 U4614 ( .A(\u_cordic/mycordic/n382 ), .Q(n1469) );
  AOI221 U4615 ( .A(\u_cordic/mycordic/N316 ), .B(n772), .C(
        \u_cordic/mycordic/N348 ), .D(n1904), .Q(\u_cordic/mycordic/n382 ) );
  XOR21 U4616 ( .A(\u_cordic/mycordic/present_I_table[2][0] ), .B(
        \u_cordic/mycordic/present_Q_table[2][1] ), .Q(
        \u_cordic/mycordic/N316 ) );
  XNR21 U4617 ( .A(\u_cordic/mycordic/present_I_table[2][0] ), .B(n173), .Q(
        \u_cordic/mycordic/N348 ) );
  INV3 U4618 ( .A(\u_cordic/mycordic/n374 ), .Q(n1562) );
  AOI221 U4619 ( .A(\u_cordic/mycordic/N380 ), .B(\u_cordic/mycordic/n332 ), 
        .C(\u_cordic/mycordic/N412 ), .D(n1908), .Q(\u_cordic/mycordic/n374 )
         );
  XOR21 U4620 ( .A(\u_cordic/mycordic/present_I_table[3][0] ), .B(
        \u_cordic/mycordic/present_Q_table[3][2] ), .Q(
        \u_cordic/mycordic/N380 ) );
  XNR21 U4621 ( .A(\u_cordic/mycordic/present_I_table[3][0] ), .B(n174), .Q(
        \u_cordic/mycordic/N412 ) );
  INV3 U4622 ( .A(\u_cordic/mycordic/n517 ), .Q(n1455) );
  AOI221 U4623 ( .A(\u_cordic/mycordic/N334 ), .B(n772), .C(
        \u_cordic/mycordic/N366 ), .D(n1904), .Q(\u_cordic/mycordic/n517 ) );
  XNR21 U4624 ( .A(\u_cordic/mycordic/present_ANGLE_table[1][2] ), .B(
        \u_cordic/mycordic/sub_196/carry[2] ), .Q(\u_cordic/mycordic/N366 ) );
  XOR21 U4625 ( .A(\u_cordic/mycordic/present_ANGLE_table[1][2] ), .B(
        \u_cordic/mycordic/add_191/carry[2] ), .Q(\u_cordic/mycordic/N334 ) );
  INV3 U4626 ( .A(\u_cordic/mycordic/n499 ), .Q(n1550) );
  AOI221 U4627 ( .A(\u_cordic/mycordic/N400 ), .B(\u_cordic/mycordic/n332 ), 
        .C(\u_cordic/mycordic/N432 ), .D(n1908), .Q(\u_cordic/mycordic/n499 )
         );
  XNR21 U4628 ( .A(\u_cordic/mycordic/present_ANGLE_table[2][4] ), .B(
        \u_cordic/mycordic/sub_207/carry [4]), .Q(\u_cordic/mycordic/N432 ) );
  XOR21 U4629 ( .A(\u_cordic/mycordic/present_ANGLE_table[2][4] ), .B(
        \u_cordic/mycordic/add_202/carry [4]), .Q(\u_cordic/mycordic/N400 ) );
  INV3 U4630 ( .A(\u_cordic/mycordic/n484 ), .Q(n1524) );
  AOI221 U4631 ( .A(\u_cordic/mycordic/N459 ), .B(\u_cordic/mycordic/n363 ), 
        .C(\u_cordic/mycordic/N487 ), .D(n1907), .Q(\u_cordic/mycordic/n484 )
         );
  XNR21 U4632 ( .A(\u_cordic/mycordic/present_ANGLE_table[3][3] ), .B(
        \u_cordic/mycordic/sub_218/carry[3] ), .Q(\u_cordic/mycordic/N487 ) );
  XOR21 U4633 ( .A(\u_cordic/mycordic/present_ANGLE_table[3][3] ), .B(
        \u_cordic/mycordic/add_213/carry[3] ), .Q(\u_cordic/mycordic/N459 ) );
  INV3 U4634 ( .A(\u_cordic/mycordic/n469 ), .Q(n1499) );
  AOI221 U4635 ( .A(\u_cordic/mycordic/N503 ), .B(n776), .C(
        \u_cordic/mycordic/N520 ), .D(n1906), .Q(\u_cordic/mycordic/n469 ) );
  XNR21 U4636 ( .A(\u_cordic/mycordic/present_ANGLE_table[4][2] ), .B(
        \u_cordic/mycordic/sub_229/carry[2] ), .Q(\u_cordic/mycordic/N520 ) );
  XOR21 U4637 ( .A(\u_cordic/mycordic/present_ANGLE_table[4][2] ), .B(
        \u_cordic/mycordic/add_224/carry[2] ), .Q(\u_cordic/mycordic/N503 ) );
  INV3 U4638 ( .A(\u_cordic/mycordic/n468 ), .Q(n1500) );
  AOI221 U4639 ( .A(\u_cordic/mycordic/N504 ), .B(\u_cordic/mycordic/n456 ), 
        .C(\u_cordic/mycordic/N521 ), .D(n1906), .Q(\u_cordic/mycordic/n468 )
         );
  XNR21 U4640 ( .A(\u_cordic/mycordic/present_ANGLE_table[4][3] ), .B(
        \u_cordic/mycordic/sub_229/carry[3] ), .Q(\u_cordic/mycordic/N521 ) );
  XOR21 U4641 ( .A(\u_cordic/mycordic/present_ANGLE_table[4][3] ), .B(
        \u_cordic/mycordic/add_224/carry[3] ), .Q(\u_cordic/mycordic/N504 ) );
  INV3 U4642 ( .A(\u_cordic/mycordic/n394 ), .Q(n1429) );
  AOI221 U4643 ( .A(\u_cordic/mycordic/present_I_table[0][4] ), .B(
        \u_cordic/mycordic/n354 ), .C(\u_cordic/mycordic/N236 ), .D(n1901), 
        .Q(\u_cordic/mycordic/n394 ) );
  XOR21 U4644 ( .A(n261), .B(n58), .Q(\u_cordic/mycordic/N236 ) );
  INV3 U4645 ( .A(\u_cordic/mycordic/n518 ), .Q(n1454) );
  AOI221 U4646 ( .A(\u_cordic/mycordic/N333 ), .B(\u_cordic/mycordic/n336 ), 
        .C(\u_cordic/mycordic/N365 ), .D(n1904), .Q(\u_cordic/mycordic/n518 )
         );
  XOR21 U4647 ( .A(\u_cordic/mycordic/present_ANGLE_table[1][1] ), .B(
        \u_cordic/mycordic/present_ANGLE_table[1][0] ), .Q(
        \u_cordic/mycordic/N365 ) );
  XNR21 U4648 ( .A(\u_cordic/mycordic/present_ANGLE_table[1][1] ), .B(
        \u_cordic/mycordic/present_ANGLE_table[1][0] ), .Q(
        \u_cordic/mycordic/N333 ) );
  INV3 U4649 ( .A(\u_cordic/mycordic/n501 ), .Q(n1548) );
  AOI221 U4650 ( .A(\u_cordic/mycordic/N398 ), .B(\u_cordic/mycordic/n332 ), 
        .C(\u_cordic/mycordic/N430 ), .D(n1908), .Q(\u_cordic/mycordic/n501 )
         );
  XOR21 U4651 ( .A(\u_cordic/mycordic/present_ANGLE_table[2][2] ), .B(
        \u_cordic/mycordic/present_ANGLE_table[2][1] ), .Q(
        \u_cordic/mycordic/N430 ) );
  XNR21 U4652 ( .A(\u_cordic/mycordic/present_ANGLE_table[2][2] ), .B(
        \u_cordic/mycordic/present_ANGLE_table[2][1] ), .Q(
        \u_cordic/mycordic/N398 ) );
  INV3 U4653 ( .A(\u_cordic/mycordic/n470 ), .Q(n1498) );
  AOI221 U4654 ( .A(\u_cordic/mycordic/N502 ), .B(\u_cordic/mycordic/n456 ), 
        .C(\u_cordic/mycordic/N519 ), .D(n1906), .Q(\u_cordic/mycordic/n470 )
         );
  XOR21 U4655 ( .A(\u_cordic/mycordic/present_ANGLE_table[4][1] ), .B(
        \u_cordic/mycordic/present_ANGLE_table[4][0] ), .Q(
        \u_cordic/mycordic/N519 ) );
  XNR21 U4656 ( .A(\u_cordic/mycordic/present_ANGLE_table[4][1] ), .B(
        \u_cordic/mycordic/present_ANGLE_table[4][0] ), .Q(
        \u_cordic/mycordic/N502 ) );
  INV3 U4657 ( .A(\u_cordic/mycordic/n357 ), .Q(n1433) );
  AOI221 U4658 ( .A(n1901), .B(\u_cordic/mycordic/N244 ), .C(
        \u_cordic/mycordic/n354 ), .D(
        \u_cordic/mycordic/present_Q_table[0][4] ), .Q(
        \u_cordic/mycordic/n357 ) );
  XOR21 U4659 ( .A(n260), .B(n55), .Q(\u_cordic/mycordic/N244 ) );
  INV3 U4660 ( .A(\u_cordic/mycordic/n356 ), .Q(n1434) );
  AOI221 U4661 ( .A(n1901), .B(\u_cordic/mycordic/N245 ), .C(
        \u_cordic/mycordic/n354 ), .D(
        \u_cordic/mycordic/present_Q_table[0][5] ), .Q(
        \u_cordic/mycordic/n356 ) );
  XOR21 U4662 ( .A(\u_cordic/mycordic/sub_add_151_b0/carry [5]), .B(n54), .Q(
        \u_cordic/mycordic/N245 ) );
  INV3 U4663 ( .A(\u_cordic/mycordic/n516 ), .Q(n1456) );
  AOI221 U4664 ( .A(\u_cordic/mycordic/N335 ), .B(\u_cordic/mycordic/n336 ), 
        .C(\u_cordic/mycordic/N367 ), .D(n1904), .Q(\u_cordic/mycordic/n516 )
         );
  XOR21 U4665 ( .A(\u_cordic/mycordic/present_ANGLE_table[1][3] ), .B(
        \u_cordic/mycordic/sub_196/carry[3] ), .Q(\u_cordic/mycordic/N367 ) );
  XNR21 U4666 ( .A(\u_cordic/mycordic/present_ANGLE_table[1][3] ), .B(
        \u_cordic/mycordic/add_191/carry[3] ), .Q(\u_cordic/mycordic/N335 ) );
  INV3 U4667 ( .A(\u_cordic/mycordic/n503 ), .Q(n1546) );
  AOI221 U4668 ( .A(\u_cordic/mycordic/N428 ), .B(\u_cordic/mycordic/n332 ), 
        .C(\u_cordic/mycordic/N428 ), .D(n1908), .Q(\u_cordic/mycordic/n503 )
         );
  INV3 U4669 ( .A(\u_cordic/mycordic/n343 ), .Q(n1477) );
  AOI221 U4670 ( .A(\u_cordic/mycordic/N324 ), .B(n772), .C(
        \u_cordic/mycordic/N356 ), .D(n1904), .Q(\u_cordic/mycordic/n343 ) );
  XOR21 U4671 ( .A(\u_cordic/mycordic/present_Q_table[2][0] ), .B(
        \u_cordic/mycordic/present_I_table[2][1] ), .Q(
        \u_cordic/mycordic/N356 ) );
  XNR21 U4672 ( .A(\u_cordic/mycordic/present_Q_table[2][0] ), .B(n175), .Q(
        \u_cordic/mycordic/N324 ) );
  INV3 U4673 ( .A(\u_cordic/mycordic/n334 ), .Q(n1570) );
  AOI221 U4674 ( .A(\u_cordic/mycordic/N388 ), .B(\u_cordic/mycordic/n332 ), 
        .C(\u_cordic/mycordic/N420 ), .D(n1908), .Q(\u_cordic/mycordic/n334 )
         );
  XOR21 U4675 ( .A(\u_cordic/mycordic/present_Q_table[3][0] ), .B(
        \u_cordic/mycordic/present_I_table[3][2] ), .Q(
        \u_cordic/mycordic/N420 ) );
  XNR21 U4676 ( .A(\u_cordic/mycordic/present_Q_table[3][0] ), .B(n176), .Q(
        \u_cordic/mycordic/N388 ) );
  INV3 U4677 ( .A(\u_cordic/mycordic/n500 ), .Q(n1549) );
  AOI221 U4678 ( .A(\u_cordic/mycordic/N399 ), .B(n778), .C(
        \u_cordic/mycordic/N431 ), .D(n1908), .Q(\u_cordic/mycordic/n500 ) );
  XOR21 U4679 ( .A(\u_cordic/mycordic/present_ANGLE_table[2][3] ), .B(
        \u_cordic/mycordic/sub_207/carry [3]), .Q(\u_cordic/mycordic/N431 ) );
  XNR21 U4680 ( .A(\u_cordic/mycordic/present_ANGLE_table[2][3] ), .B(
        \u_cordic/mycordic/add_202/carry [3]), .Q(\u_cordic/mycordic/N399 ) );
  INV3 U4681 ( .A(\u_cordic/mycordic/n485 ), .Q(n1523) );
  AOI221 U4682 ( .A(\u_cordic/mycordic/N458 ), .B(n777), .C(
        \u_cordic/mycordic/N486 ), .D(n1907), .Q(\u_cordic/mycordic/n485 ) );
  XOR21 U4683 ( .A(\u_cordic/mycordic/present_ANGLE_table[3][2] ), .B(
        \u_cordic/mycordic/sub_218/carry[2] ), .Q(\u_cordic/mycordic/N486 ) );
  XNR21 U4684 ( .A(\u_cordic/mycordic/present_ANGLE_table[3][2] ), .B(
        \u_cordic/mycordic/add_213/carry[2] ), .Q(\u_cordic/mycordic/N458 ) );
  INV3 U4685 ( .A(\u_decoder/iq_demod/n58 ), .Q(n2379) );
  AOI311 U4686 ( .A(\u_decoder/iq_demod/state [1]), .B(
        \u_decoder/iq_demod/n59 ), .C(\u_decoder/sample_ready ), .D(n779), .Q(
        \u_decoder/iq_demod/n58 ) );
  INV3 U4687 ( .A(\u_decoder/iq_demod/cossin_dig/n36 ), .Q(n2684) );
  AOI221 U4688 ( .A(\u_decoder/iq_demod/cossin_dig/N60 ), .B(n2685), .C(
        \u_decoder/iq_demod/sin_out [3]), .D(n756), .Q(
        \u_decoder/iq_demod/cossin_dig/n36 ) );
  INV3 U4689 ( .A(\u_decoder/iq_demod/cossin_dig/n31 ), .Q(n2685) );
  INV3 U4690 ( .A(\u_cordic/mycordic/n519 ), .Q(n1453) );
  AOI221 U4691 ( .A(n297), .B(n772), .C(n297), .D(n1904), .Q(
        \u_cordic/mycordic/n519 ) );
  INV3 U4692 ( .A(\u_cordic/mycordic/n502 ), .Q(n1547) );
  AOI221 U4693 ( .A(n298), .B(n778), .C(n298), .D(n1908), .Q(
        \u_cordic/mycordic/n502 ) );
  INV3 U4694 ( .A(\u_cordic/mycordic/n471 ), .Q(n1497) );
  AOI221 U4695 ( .A(n299), .B(\u_cordic/mycordic/n456 ), .C(n299), .D(n1906), 
        .Q(\u_cordic/mycordic/n471 ) );
  INV3 U4696 ( .A(\u_decoder/iq_demod/n67 ), .Q(n1574) );
  AOI221 U4697 ( .A(sig_DEMUX_outDEMUX18[2]), .B(n1910), .C(
        \u_decoder/iq_demod/I_if_signed [2]), .D(\u_decoder/iq_demod/n61 ), 
        .Q(\u_decoder/iq_demod/n67 ) );
  NOR21 U4698 ( .A(in_DEMUX_inSEL17), .B(n2120), .Q(sig_DEMUX_outDEMUX18[2])
         );
  INV3 U4699 ( .A(\u_decoder/iq_demod/n66 ), .Q(n1575) );
  AOI221 U4700 ( .A(sig_DEMUX_outDEMUX18[1]), .B(n1910), .C(
        \u_decoder/iq_demod/I_if_signed [1]), .D(\u_decoder/iq_demod/n61 ), 
        .Q(\u_decoder/iq_demod/n66 ) );
  NOR21 U4701 ( .A(in_DEMUX_inSEL17), .B(n2122), .Q(sig_DEMUX_outDEMUX18[1])
         );
  INV3 U4702 ( .A(\u_decoder/iq_demod/n65 ), .Q(n1576) );
  AOI221 U4703 ( .A(sig_DEMUX_outDEMUX18[0]), .B(n1910), .C(
        \u_decoder/iq_demod/I_if_signed [0]), .D(\u_decoder/iq_demod/n61 ), 
        .Q(\u_decoder/iq_demod/n65 ) );
  NOR21 U4704 ( .A(in_DEMUX_inSEL17), .B(n2124), .Q(sig_DEMUX_outDEMUX18[0])
         );
  INV3 U4705 ( .A(\u_decoder/iq_demod/n63 ), .Q(n1578) );
  AOI221 U4706 ( .A(sig_DEMUX_outDEMUX17[2]), .B(n1910), .C(
        \u_decoder/iq_demod/Q_if_signed [2]), .D(\u_decoder/iq_demod/n61 ), 
        .Q(\u_decoder/iq_demod/n63 ) );
  NOR21 U4707 ( .A(in_DEMUX_inSEL17), .B(n2112), .Q(sig_DEMUX_outDEMUX17[2])
         );
  INV3 U4708 ( .A(\u_decoder/iq_demod/n62 ), .Q(n1579) );
  AOI221 U4709 ( .A(sig_DEMUX_outDEMUX17[1]), .B(n1910), .C(
        \u_decoder/iq_demod/Q_if_signed [1]), .D(\u_decoder/iq_demod/n61 ), 
        .Q(\u_decoder/iq_demod/n62 ) );
  NOR21 U4710 ( .A(in_DEMUX_inSEL17), .B(n2114), .Q(sig_DEMUX_outDEMUX17[1])
         );
  INV3 U4711 ( .A(\u_decoder/iq_demod/n60 ), .Q(n1580) );
  AOI221 U4712 ( .A(sig_DEMUX_outDEMUX17[0]), .B(n1910), .C(
        \u_decoder/iq_demod/Q_if_signed [0]), .D(\u_decoder/iq_demod/n61 ), 
        .Q(\u_decoder/iq_demod/n60 ) );
  NOR21 U4713 ( .A(in_DEMUX_inSEL17), .B(n2116), .Q(sig_DEMUX_outDEMUX17[0])
         );
  INV3 U4714 ( .A(n3053), .Q(n1831) );
  NAND22 U4715 ( .A(n1218), .B(n2206), .Q(n3053) );
  INV3 U4716 ( .A(\u_cdr/phd1/n12 ), .Q(n2206) );
  AOI221 U4717 ( .A(n319), .B(\u_cdr/phd1/w_s3 ), .C(\u_cdr/dir ), .D(
        \u_cdr/phd1/w_en_m ), .Q(\u_cdr/phd1/n12 ) );
  INV3 U4718 ( .A(\u_cdr/phd1/f1/n2 ), .Q(n1844) );
  NAND22 U4719 ( .A(n1218), .B(n2207), .Q(\u_cdr/phd1/f1/n2 ) );
  INV3 U4720 ( .A(\u_cdr/phd1/n14 ), .Q(n2207) );
  AOI221 U4721 ( .A(n2689), .B(\u_cdr/dir ), .C(\u_cdr/phd1/w_s1 ), .D(
        \u_cdr/phd1/n15 ), .Q(\u_cdr/phd1/n14 ) );
  INV3 U4722 ( .A(\u_decoder/iq_demod/cossin_dig/n38 ), .Q(n1846) );
  NAND22 U4723 ( .A(\u_decoder/iq_demod/cossin_dig/n39 ), .B(
        \u_decoder/iq_demod/cossin_dig/val_counter [2]), .Q(
        \u_decoder/iq_demod/cossin_dig/n38 ) );
  INV3 U4724 ( .A(\u_cordic/my_rotation/n74 ), .Q(n1856) );
  NAND22 U4725 ( .A(\u_cordic/cordic_to_rotation [15]), .B(n1216), .Q(
        \u_cordic/my_rotation/n74 ) );
  INV3 U4726 ( .A(\u_cordic/my_rotation/n75 ), .Q(n1857) );
  NAND22 U4727 ( .A(\u_cordic/cordic_to_rotation [14]), .B(n1216), .Q(
        \u_cordic/my_rotation/n75 ) );
  INV3 U4728 ( .A(\u_cordic/my_rotation/n76 ), .Q(n1858) );
  NAND22 U4729 ( .A(\u_cordic/cordic_to_rotation [13]), .B(n1216), .Q(
        \u_cordic/my_rotation/n76 ) );
  INV3 U4730 ( .A(\u_cordic/my_rotation/n77 ), .Q(n1859) );
  NAND22 U4731 ( .A(\u_cordic/cordic_to_rotation [12]), .B(n1216), .Q(
        \u_cordic/my_rotation/n77 ) );
  INV3 U4732 ( .A(\u_cordic/my_rotation/n78 ), .Q(n1860) );
  NAND22 U4733 ( .A(\u_cordic/cordic_to_rotation [11]), .B(n1216), .Q(
        \u_cordic/my_rotation/n78 ) );
  INV3 U4734 ( .A(\u_cordic/my_rotation/n79 ), .Q(n1861) );
  NAND22 U4735 ( .A(\u_cordic/cordic_to_rotation [10]), .B(n1216), .Q(
        \u_cordic/my_rotation/n79 ) );
  INV3 U4736 ( .A(\u_cordic/my_rotation/n80 ), .Q(n1862) );
  NAND22 U4737 ( .A(\u_cordic/cordic_to_rotation [9]), .B(n1216), .Q(
        \u_cordic/my_rotation/n80 ) );
  INV3 U4738 ( .A(\u_cordic/my_rotation/n81 ), .Q(n1863) );
  NAND22 U4739 ( .A(\u_cordic/cordic_to_rotation [8]), .B(n1216), .Q(
        \u_cordic/my_rotation/n81 ) );
  INV3 U4740 ( .A(\u_cordic/my_rotation/n82 ), .Q(n1864) );
  NAND22 U4741 ( .A(\u_cordic/cordic_to_rotation [7]), .B(n1216), .Q(
        \u_cordic/my_rotation/n82 ) );
  INV3 U4742 ( .A(\u_cordic/my_rotation/n83 ), .Q(n1865) );
  NAND22 U4743 ( .A(\u_cordic/cordic_to_rotation [6]), .B(n1215), .Q(
        \u_cordic/my_rotation/n83 ) );
  INV3 U4744 ( .A(\u_cordic/my_rotation/n84 ), .Q(n1866) );
  NAND22 U4745 ( .A(\u_cordic/cordic_to_rotation [5]), .B(n1215), .Q(
        \u_cordic/my_rotation/n84 ) );
  INV3 U4746 ( .A(\u_cordic/my_rotation/n85 ), .Q(n1867) );
  NAND22 U4747 ( .A(\u_cordic/cordic_to_rotation [4]), .B(n1215), .Q(
        \u_cordic/my_rotation/n85 ) );
  INV3 U4748 ( .A(\u_cordic/my_rotation/n50 ), .Q(n1852) );
  NAND22 U4749 ( .A(\u_cordic/cordic_to_rotation [2]), .B(n1216), .Q(
        \u_cordic/my_rotation/n50 ) );
  INV3 U4750 ( .A(\u_cordic/my_rotation/n51 ), .Q(n1853) );
  NAND22 U4751 ( .A(\u_cordic/cordic_to_rotation [1]), .B(n1216), .Q(
        \u_cordic/my_rotation/n51 ) );
  INV3 U4752 ( .A(\u_cordic/my_rotation/n52 ), .Q(n1854) );
  NAND22 U4753 ( .A(\u_cordic/cordic_to_rotation [0]), .B(n1216), .Q(
        \u_cordic/my_rotation/n52 ) );
  INV3 U4754 ( .A(\u_cordic/mycordic/n429 ), .Q(n1898) );
  NAND22 U4755 ( .A(\u_cordic/mycordic/present_C_table[1][2] ), .B(n1213), .Q(
        \u_cordic/mycordic/n429 ) );
  INV3 U4756 ( .A(\u_cordic/mycordic/n426 ), .Q(n1895) );
  NAND22 U4757 ( .A(\u_cordic/mycordic/present_C_table[2][2] ), .B(n1213), .Q(
        \u_cordic/mycordic/n426 ) );
  INV3 U4758 ( .A(\u_cordic/mycordic/n422 ), .Q(n1891) );
  NAND22 U4759 ( .A(\u_cordic/mycordic/present_C_table[3][2] ), .B(n1213), .Q(
        \u_cordic/mycordic/n422 ) );
  INV3 U4760 ( .A(\u_cordic/mycordic/n419 ), .Q(n1888) );
  NAND22 U4761 ( .A(\u_cordic/mycordic/present_C_table[4][2] ), .B(n1214), .Q(
        \u_cordic/mycordic/n419 ) );
  INV3 U4762 ( .A(\u_cordic/mycordic/n416 ), .Q(n1885) );
  NAND22 U4763 ( .A(\u_cordic/mycordic/present_C_table[5][2] ), .B(n1214), .Q(
        \u_cordic/mycordic/n416 ) );
  INV3 U4764 ( .A(\u_cordic/mycordic/n412 ), .Q(n1881) );
  NAND22 U4765 ( .A(\u_cordic/mycordic/present_C_table[6][2] ), .B(n1214), .Q(
        \u_cordic/mycordic/n412 ) );
  INV3 U4766 ( .A(\u_cordic/mycordic/n430 ), .Q(n1899) );
  NAND22 U4767 ( .A(\u_cordic/mycordic/present_C_table[1][1] ), .B(n1213), .Q(
        \u_cordic/mycordic/n430 ) );
  INV3 U4768 ( .A(\u_cordic/mycordic/n427 ), .Q(n1896) );
  NAND22 U4769 ( .A(\u_cordic/mycordic/present_C_table[2][1] ), .B(n1213), .Q(
        \u_cordic/mycordic/n427 ) );
  INV3 U4770 ( .A(\u_cordic/mycordic/n423 ), .Q(n1892) );
  NAND22 U4771 ( .A(\u_cordic/mycordic/present_C_table[3][1] ), .B(n1213), .Q(
        \u_cordic/mycordic/n423 ) );
  INV3 U4772 ( .A(\u_cordic/mycordic/n420 ), .Q(n1889) );
  NAND22 U4773 ( .A(\u_cordic/mycordic/present_C_table[4][1] ), .B(n1214), .Q(
        \u_cordic/mycordic/n420 ) );
  INV3 U4774 ( .A(\u_cordic/mycordic/n417 ), .Q(n1886) );
  NAND22 U4775 ( .A(\u_cordic/mycordic/present_C_table[5][1] ), .B(n1214), .Q(
        \u_cordic/mycordic/n417 ) );
  INV3 U4776 ( .A(\u_cordic/mycordic/n414 ), .Q(n1883) );
  NAND22 U4777 ( .A(\u_cordic/mycordic/present_C_table[6][1] ), .B(n1214), .Q(
        \u_cordic/mycordic/n414 ) );
  INV3 U4778 ( .A(\u_cordic/mycordic/n431 ), .Q(n1900) );
  NAND22 U4779 ( .A(\u_cordic/mycordic/present_C_table[1][0] ), .B(n1213), .Q(
        \u_cordic/mycordic/n431 ) );
  INV3 U4780 ( .A(\u_cordic/mycordic/n428 ), .Q(n1897) );
  NAND22 U4781 ( .A(\u_cordic/mycordic/present_C_table[2][0] ), .B(n1213), .Q(
        \u_cordic/mycordic/n428 ) );
  INV3 U4782 ( .A(\u_cordic/mycordic/n425 ), .Q(n1894) );
  NAND22 U4783 ( .A(\u_cordic/mycordic/present_C_table[3][0] ), .B(n1213), .Q(
        \u_cordic/mycordic/n425 ) );
  INV3 U4784 ( .A(\u_cordic/mycordic/n421 ), .Q(n1890) );
  NAND22 U4785 ( .A(\u_cordic/mycordic/present_C_table[4][0] ), .B(n1214), .Q(
        \u_cordic/mycordic/n421 ) );
  INV3 U4786 ( .A(\u_cordic/mycordic/n418 ), .Q(n1887) );
  NAND22 U4787 ( .A(\u_cordic/mycordic/present_C_table[5][0] ), .B(n1214), .Q(
        \u_cordic/mycordic/n418 ) );
  INV3 U4788 ( .A(\u_cordic/mycordic/n415 ), .Q(n1884) );
  NAND22 U4789 ( .A(\u_cordic/mycordic/present_C_table[6][0] ), .B(n1214), .Q(
        \u_cordic/mycordic/n415 ) );
  NOR21 U4790 ( .A(\u_decoder/iq_demod/state [0]), .B(\u_decoder/iq_demod/n69 ), .Q(\u_decoder/iq_demod/N13 ) );
  NOR21 U4791 ( .A(n1239), .B(\u_coder/n131 ), .Q(\u_coder/N501 ) );
  NOR21 U4792 ( .A(n1239), .B(\u_coder/n130 ), .Q(\u_coder/N499 ) );
  INV3 U4793 ( .A(\u_decoder/iq_demod/n68 ), .Q(n1573) );
  AOI221 U4794 ( .A(\u_decoder/iq_demod/I_if_buff[3] ), .B(
        \u_decoder/iq_demod/n61 ), .C(n1910), .D(sig_DEMUX_outDEMUX18[3]), .Q(
        \u_decoder/iq_demod/n68 ) );
  NOR21 U4795 ( .A(in_DEMUX_inSEL17), .B(n2118), .Q(sig_DEMUX_outDEMUX18[3])
         );
  INV3 U4796 ( .A(\u_decoder/iq_demod/n64 ), .Q(n1577) );
  AOI221 U4797 ( .A(\u_decoder/iq_demod/Q_if_buff[3] ), .B(
        \u_decoder/iq_demod/n61 ), .C(n1910), .D(sig_DEMUX_outDEMUX17[3]), .Q(
        \u_decoder/iq_demod/n64 ) );
  NOR21 U4798 ( .A(in_DEMUX_inSEL17), .B(n2110), .Q(sig_DEMUX_outDEMUX17[3])
         );
  INV3 U4799 ( .A(n3073), .Q(n1841) );
  NAND22 U4800 ( .A(n1219), .B(\u_outFIFO/os1/sigQout1 ), .Q(n3073) );
  INV3 U4801 ( .A(n3069), .Q(n1837) );
  NAND22 U4802 ( .A(n1218), .B(\u_inFIFO/os1/sigQout1 ), .Q(n3069) );
  INV3 U4803 ( .A(n3071), .Q(n1839) );
  NAND22 U4804 ( .A(n1218), .B(\u_inFIFO/os2/sigQout1 ), .Q(n3071) );
  INV3 U4805 ( .A(n3075), .Q(n1843) );
  NAND22 U4806 ( .A(n1218), .B(\u_outFIFO/os2/sigQout1 ), .Q(n3075) );
  INV3 U4807 ( .A(\u_cordic/my_rotation/n49 ), .Q(n1851) );
  NAND22 U4808 ( .A(n1218), .B(\u_cordic/cordic_to_rotation [3]), .Q(
        \u_cordic/my_rotation/n49 ) );
  INV3 U4809 ( .A(in_DEMUX_inSEL17), .Q(n2140) );
  INV3 U4810 ( .A(in_MUX_inSEL6[0]), .Q(n2133) );
  INV3 U4811 ( .A(\u_inFIFO/n222 ), .Q(n1958) );
  NAND22 U4812 ( .A(in_inFIFO_inData[3]), .B(n1217), .Q(\u_inFIFO/n222 ) );
  INV3 U4813 ( .A(\u_inFIFO/n221 ), .Q(n1957) );
  NAND22 U4814 ( .A(in_inFIFO_inData[2]), .B(n1217), .Q(\u_inFIFO/n221 ) );
  INV3 U4815 ( .A(\u_inFIFO/n220 ), .Q(n1956) );
  NAND22 U4816 ( .A(in_inFIFO_inData[1]), .B(n1217), .Q(\u_inFIFO/n220 ) );
  INV3 U4817 ( .A(\u_inFIFO/n219 ), .Q(n1955) );
  NAND22 U4818 ( .A(in_inFIFO_inData[0]), .B(n1217), .Q(\u_inFIFO/n219 ) );
  NAND22 U4819 ( .A(in_DEMUX_inDEMUX1), .B(n2127), .Q(\u_demux1/n5 ) );
  INV3 U4820 ( .A(in_DEMUX_inSEL1[0]), .Q(n2127) );
  NAND22 U4821 ( .A(in_DEMUX_inDEMUX2), .B(n2130), .Q(n3118) );
  INV3 U4822 ( .A(in_DEMUX_inSEL2[0]), .Q(n2130) );
  INV3 U4823 ( .A(in_MUX_inSEL9[0]), .Q(n2135) );
  INV3 U4824 ( .A(in_MUX_inSEL9[1]), .Q(n2134) );
  NOR31 U4825 ( .A(\u_demux1/n5 ), .B(in_DEMUX_inSEL1[2]), .C(
        in_DEMUX_inSEL1[1]), .Q(sig_DEMUX_outDEMUX1[0]) );
  NAND22 U4826 ( .A(in_DEMUX_inSEL1[0]), .B(in_DEMUX_inDEMUX1), .Q(
        \u_demux1/n4 ) );
  NAND22 U4827 ( .A(in_DEMUX_inSEL2[0]), .B(in_DEMUX_inDEMUX2), .Q(n3117) );
  INV3 U4828 ( .A(inReset), .Q(n1235) );
  INV3 U4829 ( .A(inReset), .Q(n1233) );
  INV3 U4830 ( .A(inReset), .Q(n1234) );
  INV3 U4831 ( .A(inReset), .Q(n1232) );
  AOI221 U4832 ( .A(\sig_MUX_inMUX14[0] ), .B(n2139), .C(\sig_MUX_inMUX13[0] ), 
        .D(in_MUX_inSEL15[0]), .Q(n3076) );
  AOI221 U4833 ( .A(\sig_MUX_inMUX5[0] ), .B(n2139), .C(in_MUX_inSEL15[0]), 
        .D(\sig_MUX_inMUX8[0] ), .Q(n3077) );
  NAND22 U4834 ( .A(sig_decod_outQ[0]), .B(n2135), .Q(n3088) );
  AOI221 U4835 ( .A(sig_coder_outSinQ[0]), .B(n2135), .C(in_MUX_inSEL9[0]), 
        .D(sig_coder_outSinQMasked[0]), .Q(n3089) );
  NAND22 U4836 ( .A(sig_decod_outQ[1]), .B(n2135), .Q(n3090) );
  AOI221 U4837 ( .A(sig_coder_outSinQ[1]), .B(n2135), .C(in_MUX_inSEL9[0]), 
        .D(sig_coder_outSinQMasked[1]), .Q(n3091) );
  NAND22 U4838 ( .A(sig_decod_outQ[2]), .B(n2135), .Q(n3092) );
  AOI221 U4839 ( .A(sig_coder_outSinQ[2]), .B(n2135), .C(in_MUX_inSEL9[0]), 
        .D(sig_coder_outSinQMasked[2]), .Q(n3093) );
  AOI221 U4840 ( .A(sig_decod_outI[0]), .B(n2135), .C(sig_outFIFO_outData[0]), 
        .D(in_MUX_inSEL9[0]), .Q(n3080) );
  AOI221 U4841 ( .A(sig_coder_outSinI[0]), .B(n2135), .C(in_MUX_inSEL9[0]), 
        .D(sig_coder_outSinIMasked[0]), .Q(n3081) );
  NAND22 U4842 ( .A(sig_decod_outQ[3]), .B(n2135), .Q(n3094) );
  AOI221 U4843 ( .A(sig_coder_outSinQ[3]), .B(n2135), .C(in_MUX_inSEL9[0]), 
        .D(sig_coder_outSinQMasked[3]), .Q(n3095) );
  AOI221 U4844 ( .A(n2139), .B(\sig_MUX_inMUX11[0] ), .C(in_MUX_inSEL15[0]), 
        .D(\sig_MUX_inMUX12[0] ), .Q(n3078) );
  AOI221 U4845 ( .A(\sig_MUX_inMUX4[0] ), .B(n2139), .C(in_MUX_inSEL15[0]), 
        .D(\sig_MUX_inMUX3[0] ), .Q(n3079) );
  AOI221 U4846 ( .A(sig_decod_outI[1]), .B(n2135), .C(sig_outFIFO_outData[1]), 
        .D(in_MUX_inSEL9[0]), .Q(n3082) );
  AOI221 U4847 ( .A(sig_coder_outSinI[1]), .B(n2135), .C(in_MUX_inSEL9[0]), 
        .D(sig_coder_outSinIMasked[1]), .Q(n3083) );
  AOI221 U4848 ( .A(sig_decod_outI[2]), .B(n2135), .C(sig_outFIFO_outData[2]), 
        .D(in_MUX_inSEL9[0]), .Q(n3084) );
  AOI221 U4849 ( .A(sig_coder_outSinI[2]), .B(n2135), .C(in_MUX_inSEL9[0]), 
        .D(sig_coder_outSinIMasked[2]), .Q(n3085) );
  AOI221 U4850 ( .A(sig_decod_outI[3]), .B(n2135), .C(sig_outFIFO_outData[3]), 
        .D(in_MUX_inSEL9[0]), .Q(n3086) );
  AOI221 U4851 ( .A(sig_coder_outSinI[3]), .B(n2135), .C(in_MUX_inSEL9[0]), 
        .D(sig_coder_outSinIMasked[3]), .Q(n3087) );
  INV3 U4852 ( .A(inReset), .Q(n1236) );
  INV3 U4853 ( .A(inReset), .Q(n1240) );
  INV3 U4854 ( .A(inReset), .Q(n1237) );
  INV3 U4855 ( .A(inReset), .Q(n1238) );
  NOR31 U4856 ( .A(\u_demux1/n5 ), .B(in_DEMUX_inSEL1[2]), .C(n2126), .Q(
        sig_DEMUX_outDEMUX1[2]) );
  INV3 U4857 ( .A(inReset), .Q(n1239) );
  INV3 U4858 ( .A(inReset), .Q(n1241) );
  INV3 U4859 ( .A(in_MUX_inSEL15[0]), .Q(n2139) );
  NOR31 U4860 ( .A(n2129), .B(in_DEMUX_inSEL2[2]), .C(n3117), .Q(
        sig_DEMUX_outDEMUX2[3]) );
  NOR31 U4861 ( .A(\u_demux1/n5 ), .B(in_DEMUX_inSEL1[1]), .C(n2125), .Q(
        sig_DEMUX_outDEMUX1[4]) );
  INV3 U4862 ( .A(in_DEMUX_inSEL1[2]), .Q(n2125) );
  INV3 U4863 ( .A(in_MUX_inSEL6[1]), .Q(n2132) );
  INV3 U4864 ( .A(in_MUX_inSEL3), .Q(n2131) );
  INV3 U4865 ( .A(in_DEMUX_inSEL1[1]), .Q(n2126) );
  INV3 U4866 ( .A(in_DEMUX_inSEL2[1]), .Q(n2129) );
  INV3 U4867 ( .A(in_DEMUX_inDEMUX18[3]), .Q(n2118) );
  INV3 U4868 ( .A(in_DEMUX_inDEMUX18[2]), .Q(n2120) );
  INV3 U4869 ( .A(in_DEMUX_inDEMUX18[1]), .Q(n2122) );
  INV3 U4870 ( .A(in_DEMUX_inDEMUX18[0]), .Q(n2124) );
  INV3 U4871 ( .A(in_DEMUX_inDEMUX17[3]), .Q(n2110) );
  INV3 U4872 ( .A(in_DEMUX_inDEMUX17[2]), .Q(n2112) );
  INV3 U4873 ( .A(in_DEMUX_inDEMUX17[1]), .Q(n2114) );
  INV3 U4874 ( .A(in_DEMUX_inDEMUX17[0]), .Q(n2116) );
  INV3 U4875 ( .A(in_MUX_inSEL11), .Q(n2136) );
  INV3 U4876 ( .A(in_MUX_inSEL12), .Q(n2137) );
  INV3 U4877 ( .A(in_MUX_inSEL15[1]), .Q(n2138) );
  INV3 U4878 ( .A(in_DEMUX_inSEL2[2]), .Q(n2128) );
  INV3 U4879 ( .A(n3070), .Q(n1838) );
  NAND22 U4880 ( .A(n1218), .B(sig_DEMUX_outDEMUX2[0]), .Q(n3070) );
  NOR31 U4881 ( .A(n3118), .B(in_DEMUX_inSEL2[2]), .C(in_DEMUX_inSEL2[1]), .Q(
        sig_DEMUX_outDEMUX2[0]) );
  INV3 U4882 ( .A(n3072), .Q(n1840) );
  NAND22 U4883 ( .A(n1218), .B(in_outFIFO_inReadEnable), .Q(n3072) );
  NAND22 U4884 ( .A(\u_cdr/div1/N35 ), .B(\u_cdr/w_nb_P [1]), .Q(n1302) );
  CLKIN3 U4885 ( .A(n1302), .Q(n1242) );
  NAND22 U4886 ( .A(n1257), .B(n1261), .Q(\u_cdr/div1/n32 ) );
  NAND22 U4887 ( .A(\u_cdr/div1/n32 ), .B(\u_cdr/div1/n10 ), .Q(n1245) );
  OAI212 U4888 ( .A(\u_cdr/cnt_d [1]), .B(\u_cdr/cnt_d [0]), .C(n1244), .Q(
        n1281) );
  OAI222 U4889 ( .A(\u_cdr/div1/n27 ), .B(n1245), .C(\u_cdr/div1/n10 ), .D(
        n1281), .Q(\u_cdr/div1/n38 ) );
  CLKIN3 U4890 ( .A(inClock), .Q(n1401) );
  NAND22 U4891 ( .A(n1281), .B(n221), .Q(n1253) );
  CLKIN3 U4892 ( .A(n1253), .Q(n1272) );
  NAND22 U4893 ( .A(\u_cdr/div1/n9 ), .B(\u_cdr/div1/n8 ), .Q(n1328) );
  CLKIN3 U4894 ( .A(n1328), .Q(n1322) );
  NAND22 U4895 ( .A(n1322), .B(\u_cdr/div1/n10 ), .Q(n1246) );
  CLKIN3 U4896 ( .A(n1246), .Q(n1282) );
  NAND22 U4897 ( .A(n1272), .B(n1282), .Q(n1251) );
  NAND22 U4898 ( .A(\u_cdr/div1/n31 ), .B(n1281), .Q(n1274) );
  CLKIN3 U4899 ( .A(n1281), .Q(n1271) );
  NAND22 U4900 ( .A(\u_cdr/w_nb_P [2]), .B(\u_cdr/w_nb_P [1]), .Q(n1313) );
  CLKIN3 U4901 ( .A(n1313), .Q(n1276) );
  NAND22 U4902 ( .A(\u_cdr/div1/n10 ), .B(\u_cdr/div1/n9 ), .Q(n1275) );
  OAI212 U4903 ( .A(n221), .B(n1276), .C(n1247), .Q(n1248) );
  NAND22 U4904 ( .A(n1276), .B(\u_cdr/w_nb_P [3]), .Q(n1265) );
  OAI212 U4905 ( .A(n1282), .B(n1253), .C(n1252), .Q(n1254) );
  NAND22 U4906 ( .A(n1274), .B(n1256), .Q(\u_cdr/div1/n35 ) );
  CLKIN3 U4907 ( .A(n1257), .Q(n1258) );
  CLKIN3 U4908 ( .A(\u_cdr/div1/n27 ), .Q(n1262) );
  NAND22 U4909 ( .A(n1258), .B(n1262), .Q(n1259) );
  CLKIN3 U4910 ( .A(n1259), .Q(n1279) );
  NAND22 U4911 ( .A(n1282), .B(n60), .Q(n1260) );
  XNR21 U4912 ( .A(n1260), .B(\u_cdr/w_nb_P [5]), .Q(n1269) );
  CLKIN3 U4913 ( .A(n1261), .Q(n1263) );
  NAND22 U4914 ( .A(n1263), .B(n1262), .Q(n1264) );
  CLKIN3 U4915 ( .A(n1264), .Q(n1278) );
  CLKIN3 U4916 ( .A(n1265), .Q(n1266) );
  NAND22 U4917 ( .A(n1266), .B(\u_cdr/w_nb_P [4]), .Q(n1267) );
  XNR21 U4918 ( .A(n1267), .B(\u_cdr/w_nb_P [5]), .Q(n1268) );
  OAI212 U4919 ( .A(\u_cdr/div1/n7 ), .B(n1281), .C(n1270), .Q(
        \u_cdr/div1/n39 ) );
  NAND22 U4920 ( .A(n1274), .B(n1273), .Q(\u_cdr/div1/n40 ) );
  CLKIN3 U4921 ( .A(n1275), .Q(n1284) );
  OAI212 U4922 ( .A(\u_cdr/div1/n9 ), .B(n1281), .C(n1280), .Q(
        \u_cdr/div1/n37 ) );
  NAND22 U4923 ( .A(n1282), .B(n59), .Q(n1285) );
  CLKIN3 U4924 ( .A(n1285), .Q(n1289) );
  NAND22 U4925 ( .A(n1289), .B(n60), .Q(n1288) );
  CLKIN3 U4926 ( .A(n1288), .Q(n1283) );
  OAI212 U4927 ( .A(n1283), .B(\u_cdr/div1/n7 ), .C(n1388), .Q(n1344) );
  CLKIN3 U4928 ( .A(n1344), .Q(n1378) );
  NAND22 U4929 ( .A(n1284), .B(n59), .Q(n1287) );
  CLKIN3 U4930 ( .A(n1287), .Q(n1286) );
  OAI212 U4931 ( .A(n1286), .B(\u_cdr/div1/n8 ), .C(n1285), .Q(n1292) );
  CLKIN3 U4932 ( .A(n1292), .Q(n1381) );
  CLKIN3 U4933 ( .A(n1349), .Q(n1380) );
  OAI212 U4934 ( .A(\u_cdr/div1/N35 ), .B(\u_cdr/w_nb_P [1]), .C(n1302), .Q(
        n1377) );
  CLKIN3 U4935 ( .A(n1377), .Q(n1363) );
  CLKIN3 U4936 ( .A(n1293), .Q(n1291) );
  OAI212 U4937 ( .A(n1289), .B(n60), .C(n1288), .Q(n1338) );
  CLKIN3 U4938 ( .A(n1338), .Q(n1379) );
  OAI212 U4939 ( .A(n1293), .B(n1338), .C(n1344), .Q(n1290) );
  NAND22 U4940 ( .A(n1295), .B(n1290), .Q(\u_cdr/phd1/cnt_phd/N14 ) );
  XNR21 U4941 ( .A(n1379), .B(n1291), .Q(\u_cdr/phd1/cnt_phd/N13 ) );
  NAND22 U4942 ( .A(n1349), .B(n1292), .Q(n1337) );
  NAND22 U4943 ( .A(n1388), .B(n1295), .Q(n2678) );
  NAND22 U4944 ( .A(\u_cdr/phd1/cnt_phd/cnt [0]), .B(n1377), .Q(n3047) );
  XNR21 U4945 ( .A(n1380), .B(n1363), .Q(n1400) );
  NAND22 U4946 ( .A(n1363), .B(n3055), .Q(n1294) );
  CLKIN3 U4947 ( .A(n1294), .Q(n1399) );
  NAND22 U4948 ( .A(n1388), .B(n1295), .Q(n2677) );
  CLKIN3 U4949 ( .A(n1295), .Q(\u_cdr/phd1/cnt_phd/N41 ) );
  CLKIN3 U4950 ( .A(\u_cdr/dec1/n33 ), .Q(n1420) );
  CLKIN3 U4951 ( .A(\u_cdr/dec1/n32 ), .Q(n1421) );
  CLKIN3 U4952 ( .A(\u_cdr/dec1/n26 ), .Q(n1425) );
  CLKIN3 U4953 ( .A(\u_cdr/dec1/n29 ), .Q(n1424) );
  CLKIN3 U4954 ( .A(\u_cdr/dec1/n30 ), .Q(n1423) );
  CLKIN3 U4955 ( .A(\u_cdr/dec1/n31 ), .Q(n1422) );
  XNR21 U4956 ( .A(n3055), .B(\u_cdr/div1/N35 ), .Q(n1320) );
  XNR21 U4957 ( .A(\u_cdr/phd1/cnt_phd/cnt [5]), .B(n1378), .Q(n1299) );
  XNR21 U4958 ( .A(\u_cdr/phd1/cnt_phd/cnt [4]), .B(n1379), .Q(n1298) );
  XNR21 U4959 ( .A(\u_cdr/phd1/cnt_phd/cnt [2]), .B(n1380), .Q(n1297) );
  XNR21 U4960 ( .A(\u_cdr/phd1/cnt_phd/cnt [3]), .B(n1381), .Q(n1296) );
  CLKIN3 U4961 ( .A(n1301), .Q(n1398) );
  NAND22 U4962 ( .A(n1302), .B(\u_cdr/div1/n9 ), .Q(n1312) );
  CLKIN3 U4963 ( .A(n1312), .Q(n1310) );
  NAND22 U4964 ( .A(n1310), .B(\u_cdr/div1/n8 ), .Q(n1309) );
  CLKIN3 U4965 ( .A(n1309), .Q(n1303) );
  NAND22 U4966 ( .A(n1303), .B(n60), .Q(n1305) );
  OAI212 U4967 ( .A(\u_cdr/w_nb_P [5]), .B(n1305), .C(n1320), .Q(n1319) );
  OAI212 U4968 ( .A(n1303), .B(n60), .C(n1305), .Q(n1304) );
  XNR21 U4969 ( .A(n1304), .B(\u_cdr/phd1/cnt_phd/cnt [4]), .Q(n1308) );
  NAND22 U4970 ( .A(\u_cdr/w_nb_P [5]), .B(n1305), .Q(n1306) );
  XNR21 U4971 ( .A(n255), .B(n1306), .Q(n1307) );
  NAND22 U4972 ( .A(n1308), .B(n1307), .Q(n1318) );
  OAI212 U4973 ( .A(n1310), .B(\u_cdr/div1/n8 ), .C(n1309), .Q(n1311) );
  XNR21 U4974 ( .A(n1311), .B(\u_cdr/phd1/cnt_phd/cnt [3]), .Q(n1316) );
  OAI212 U4975 ( .A(n59), .B(n1313), .C(n1312), .Q(n1314) );
  XNR21 U4976 ( .A(n1314), .B(\u_cdr/phd1/cnt_phd/cnt [2]), .Q(n1315) );
  NAND22 U4977 ( .A(n1316), .B(n1315), .Q(n1317) );
  XNR21 U4978 ( .A(\u_cdr/div1/n10 ), .B(\u_cdr/phd1/cnt_phd/cnt [1]), .Q(
        n1335) );
  NAND22 U4979 ( .A(n1322), .B(n60), .Q(n1324) );
  CLKIN3 U4980 ( .A(n1320), .Q(n1321) );
  OAI212 U4981 ( .A(\u_cdr/w_nb_P [5]), .B(n1324), .C(n1321), .Q(n1334) );
  OAI212 U4982 ( .A(n1322), .B(n60), .C(n1324), .Q(n1323) );
  XNR21 U4983 ( .A(n1323), .B(\u_cdr/phd1/cnt_phd/cnt [4]), .Q(n1327) );
  NAND22 U4984 ( .A(\u_cdr/w_nb_P [5]), .B(n1324), .Q(n1325) );
  XNR21 U4985 ( .A(n255), .B(n1325), .Q(n1326) );
  NAND22 U4986 ( .A(n1327), .B(n1326), .Q(n1333) );
  OAI212 U4987 ( .A(\u_cdr/div1/n8 ), .B(\u_cdr/div1/n9 ), .C(n1328), .Q(n1329) );
  XNR21 U4988 ( .A(n1329), .B(\u_cdr/phd1/cnt_phd/cnt [3]), .Q(n1331) );
  XNR21 U4989 ( .A(\u_cdr/div1/n9 ), .B(\u_cdr/phd1/cnt_phd/cnt [2]), .Q(n1330) );
  NAND22 U4990 ( .A(n1331), .B(n1330), .Q(n1332) );
  NAND22 U4991 ( .A(\u_cdr/dec1/w_s_r ), .B(n52), .Q(n1336) );
  CLKIN3 U4992 ( .A(n1337), .Q(n1339) );
  XOR31 U4993 ( .A(\u_cdr/dec1/cnt_r [3]), .B(n1379), .C(n1339), .Q(n1343) );
  NAND22 U4994 ( .A(n1339), .B(n1338), .Q(n1340) );
  CLKIN3 U4995 ( .A(n1340), .Q(n1345) );
  XOR31 U4996 ( .A(\u_cdr/dec1/cnt_r [4]), .B(n1378), .C(n1345), .Q(n1342) );
  NAND22 U4997 ( .A(\u_cdr/cnt_d [1]), .B(\u_cdr/cnt_d [0]), .Q(n1391) );
  NAND22 U4998 ( .A(n1345), .B(n1344), .Q(n1346) );
  XNR21 U4999 ( .A(n301), .B(n1346), .Q(n1348) );
  XOR31 U5000 ( .A(\u_cdr/dec1/cnt_r [2]), .B(n1381), .C(n1349), .Q(n1347) );
  NAND22 U5001 ( .A(n1348), .B(n1347), .Q(n1352) );
  XNR21 U5002 ( .A(n1349), .B(\u_cdr/dec1/cnt_r [1]), .Q(n1351) );
  XNR21 U5003 ( .A(n1377), .B(n248), .Q(n1350) );
  NAND22 U5004 ( .A(sig_DEMUX_outDEMUX1[4]), .B(in_MUX_inSEL12), .Q(n1354) );
  OAI212 U5005 ( .A(n52), .B(in_MUX_inSEL12), .C(n1354), .Q(n2101) );
  XNR21 U5006 ( .A(n1377), .B(\u_cdr/dec1/cnt_dec/cnt_dec [1]), .Q(n1361) );
  XNR21 U5007 ( .A(n263), .B(\u_cdr/div1/N35 ), .Q(n1360) );
  XNR21 U5008 ( .A(\u_cdr/dec1/cnt_dec/cnt_dec [5]), .B(n1378), .Q(n1358) );
  XNR21 U5009 ( .A(\u_cdr/dec1/cnt_dec/cnt_dec [4]), .B(n1379), .Q(n1357) );
  XNR21 U5010 ( .A(\u_cdr/dec1/cnt_dec/cnt_dec [2]), .B(n1380), .Q(n1356) );
  XNR21 U5011 ( .A(\u_cdr/dec1/cnt_dec/cnt_dec [3]), .B(n1381), .Q(n1355) );
  CLKIN3 U5012 ( .A(n1362), .Q(n1397) );
  XNR21 U5013 ( .A(n302), .B(n1380), .Q(n1369) );
  XNR21 U5014 ( .A(\u_cdr/dec1/cnt_dec/cnt_dec [0]), .B(n1363), .Q(n1367) );
  XNR21 U5015 ( .A(\u_cdr/dec1/cnt_dec/cnt_dec [4]), .B(n1378), .Q(n1366) );
  XNR21 U5016 ( .A(\u_cdr/dec1/cnt_dec/cnt_dec [2]), .B(n1381), .Q(n1365) );
  XNR21 U5017 ( .A(\u_cdr/dec1/cnt_dec/cnt_dec [3]), .B(n1379), .Q(n1364) );
  XNR21 U5018 ( .A(n1377), .B(\u_cdr/div1/cnt_div/cnt [1]), .Q(n1376) );
  XNR21 U5019 ( .A(n262), .B(\u_cdr/div1/N35 ), .Q(n1375) );
  XNR21 U5020 ( .A(\u_cdr/div1/cnt_div/cnt [3]), .B(n1381), .Q(n1373) );
  XNR21 U5021 ( .A(\u_cdr/div1/cnt_div/cnt [2]), .B(n1380), .Q(n1372) );
  XNR21 U5022 ( .A(\u_cdr/div1/cnt_div/cnt [4]), .B(n1379), .Q(n1371) );
  XNR21 U5023 ( .A(\u_cdr/div1/cnt_div/cnt [5]), .B(n1378), .Q(n1370) );
  CLKIN3 U5024 ( .A(n2675), .Q(n1396) );
  XNR21 U5025 ( .A(n1377), .B(\u_cdr/dec1/cnt_r [1]), .Q(n1389) );
  XNR21 U5026 ( .A(n248), .B(\u_cdr/div1/N35 ), .Q(n1387) );
  XNR21 U5027 ( .A(\u_cdr/dec1/cnt_r [5]), .B(n1378), .Q(n1385) );
  XNR21 U5028 ( .A(\u_cdr/dec1/cnt_r [4]), .B(n1379), .Q(n1384) );
  XNR21 U5029 ( .A(\u_cdr/dec1/cnt_r [2]), .B(n1380), .Q(n1383) );
  XNR21 U5030 ( .A(\u_cdr/dec1/cnt_r [3]), .B(n1381), .Q(n1382) );
  CLKIN3 U5031 ( .A(n1390), .Q(n1395) );
  CLKIN3 U5032 ( .A(n1393), .Q(n1394) );
  OAI212 U5033 ( .A(\u_inFIFO/outReadCount[2] ), .B(\u_inFIFO/n186 ), .C(n2696), .Q(n2699) );
  OAI212 U5034 ( .A(\u_inFIFO/outReadCount[6] ), .B(\u_inFIFO/n182 ), .C(n2705), .Q(n2711) );
  OAI212 U5035 ( .A(\u_outFIFO/outReadCount[2] ), .B(\u_outFIFO/n264 ), .C(
        n2749), .Q(n2752) );
  OAI212 U5036 ( .A(\u_outFIFO/outReadCount[6] ), .B(\u_outFIFO/n260 ), .C(
        n2758), .Q(n2764) );
  XNR31 U5037 ( .A(\u_decoder/iq_demod/dp_cluster_1/mult_149/A2[5] ), .B(n2396), .C(n2765), .Q(\u_decoder/iq_demod/dp_cluster_1/mult_I_sin_out [7]) );
  OAI212 U5038 ( .A(\u_decoder/iq_demod/dp_cluster_1/mult_149/A1[4] ), .B(
        n2766), .C(\u_decoder/iq_demod/dp_cluster_1/mult_149/A2[4] ), .Q(n2767) );
  XOR31 U5039 ( .A(\u_decoder/iq_demod/dp_cluster_1/mult_149/A2[4] ), .B(
        \u_decoder/iq_demod/dp_cluster_1/mult_149/A1[4] ), .C(n2766), .Q(
        \u_decoder/iq_demod/dp_cluster_1/mult_I_sin_out [6]) );
  XNR31 U5040 ( .A(\u_decoder/iq_demod/dp_cluster_1/mult_150/A2[5] ), .B(n2389), .C(n2772), .Q(\u_decoder/iq_demod/dp_cluster_1/mult_Q_cos_out [7]) );
  OAI212 U5041 ( .A(\u_decoder/iq_demod/dp_cluster_1/mult_150/A1[4] ), .B(
        n2773), .C(\u_decoder/iq_demod/dp_cluster_1/mult_150/A2[4] ), .Q(n2774) );
  XOR31 U5042 ( .A(\u_decoder/iq_demod/dp_cluster_1/mult_150/A2[4] ), .B(
        \u_decoder/iq_demod/dp_cluster_1/mult_150/A1[4] ), .C(n2773), .Q(
        \u_decoder/iq_demod/dp_cluster_1/mult_Q_cos_out [6]) );
  XNR31 U5043 ( .A(\u_decoder/iq_demod/dp_cluster_0/mult_148/A2[5] ), .B(n2397), .C(n2779), .Q(\u_decoder/iq_demod/dp_cluster_0/mult_I_cos_out [7]) );
  OAI212 U5044 ( .A(\u_decoder/iq_demod/dp_cluster_0/mult_148/A1[4] ), .B(
        n2780), .C(\u_decoder/iq_demod/dp_cluster_0/mult_148/A2[4] ), .Q(n2781) );
  XOR31 U5045 ( .A(\u_decoder/iq_demod/dp_cluster_0/mult_148/A2[4] ), .B(
        \u_decoder/iq_demod/dp_cluster_0/mult_148/A1[4] ), .C(n2780), .Q(
        \u_decoder/iq_demod/dp_cluster_0/mult_I_cos_out [6]) );
  OAI212 U5046 ( .A(\u_decoder/iq_demod/dp_cluster_0/mult_151/A1[4] ), .B(
        n2787), .C(\u_decoder/iq_demod/dp_cluster_0/mult_151/A2[4] ), .Q(n2788) );
  OAI212 U5047 ( .A(\u_decoder/fir_filter/dp_cluster_0/r177/A1[6] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r177/A2[6] ), .C(n2798), .Q(n2797)
         );
  OAI212 U5048 ( .A(\u_decoder/fir_filter/dp_cluster_0/r177/A2[6] ), .B(n2799), 
        .C(n2800), .Q(\u_decoder/fir_filter/Q_data_mult_0 [8]) );
  OAI212 U5049 ( .A(\u_decoder/fir_filter/dp_cluster_0/r177/PROD1[4] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r177/A1[3] ), .C(n2802), .Q(n2804)
         );
  OAI212 U5050 ( .A(n2376), .B(n2793), .C(
        \u_decoder/fir_filter/dp_cluster_0/r177/A2[9] ), .Q(n2806) );
  OAI212 U5051 ( .A(n2794), .B(n2368), .C(n2807), .Q(n2793) );
  OAI212 U5052 ( .A(\u_decoder/fir_filter/dp_cluster_0/r177/A1[8] ), .B(n2361), 
        .C(\u_decoder/fir_filter/dp_cluster_0/r177/A2[8] ), .Q(n2807) );
  OAI222 U5053 ( .A(\u_decoder/fir_filter/dp_cluster_0/r177/A1[6] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r177/A2[6] ), .C(
        \u_decoder/fir_filter/dp_cluster_0/r177/A1[7] ), .D(
        \u_decoder/fir_filter/dp_cluster_0/r177/A2[7] ), .Q(n2810) );
  OAI212 U5054 ( .A(\u_decoder/fir_filter/dp_cluster_0/r178/PROD1[5] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r178/A1[4] ), .C(n2816), .Q(n2818)
         );
  OAI212 U5055 ( .A(n2376), .B(n2820), .C(
        \u_decoder/fir_filter/dp_cluster_0/r178/A2[10] ), .Q(n2821) );
  OAI212 U5056 ( .A(n2310), .B(n2309), .C(n2822), .Q(n2820) );
  OAI212 U5057 ( .A(\u_decoder/fir_filter/dp_cluster_0/r178/A1[9] ), .B(n2811), 
        .C(\u_decoder/fir_filter/dp_cluster_0/r178/A2[9] ), .Q(n2822) );
  OAI212 U5058 ( .A(n2812), .B(n2311), .C(n2823), .Q(n2811) );
  OAI212 U5059 ( .A(\u_decoder/fir_filter/dp_cluster_0/r178/A1[8] ), .B(n2312), 
        .C(\u_decoder/fir_filter/dp_cluster_0/r178/A2[8] ), .Q(n2823) );
  OAI212 U5060 ( .A(\u_decoder/fir_filter/dp_cluster_0/r178/A1[7] ), .B(n2813), 
        .C(\u_decoder/fir_filter/dp_cluster_0/r178/A2[7] ), .Q(n2824) );
  OAI212 U5061 ( .A(n2317), .B(n2316), .C(n2831), .Q(n2830) );
  OAI212 U5062 ( .A(\u_decoder/fir_filter/dp_cluster_0/r179/CARRYB[7][3] ), 
        .B(n2826), .C(\u_decoder/fir_filter/dp_cluster_0/r179/A2[9] ), .Q(
        n2831) );
  OAI212 U5063 ( .A(n2827), .B(n2318), .C(n2832), .Q(n2826) );
  OAI212 U5064 ( .A(\u_decoder/fir_filter/dp_cluster_0/r179/A1[8] ), .B(n2319), 
        .C(\u_decoder/fir_filter/dp_cluster_0/r179/A2[8] ), .Q(n2832) );
  OAI212 U5065 ( .A(\u_decoder/fir_filter/dp_cluster_0/r179/A1[7] ), .B(n2322), 
        .C(\u_decoder/fir_filter/dp_cluster_0/r179/A2[7] ), .Q(n2833) );
  OAI212 U5066 ( .A(n2838), .B(n2839), .C(n2840), .Q(
        \u_decoder/fir_filter/Q_data_mult_3 [10]) );
  OAI222 U5067 ( .A(\u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[7][5] ), 
        .B(\u_decoder/fir_filter/dp_cluster_0/r180/A2[11] ), .C(
        \u_decoder/fir_filter/dp_cluster_0/r180/A1[8] ), .D(
        \u_decoder/fir_filter/dp_cluster_0/r180/A2[8] ), .Q(n2849) );
  OAI212 U5068 ( .A(\u_decoder/fir_filter/dp_cluster_0/r180/CARRYB[7][5] ), 
        .B(n2845), .C(\u_decoder/fir_filter/dp_cluster_0/r180/A2[11] ), .Q(
        n2850) );
  OAI212 U5069 ( .A(n2848), .B(n2350), .C(n2851), .Q(n2845) );
  OAI212 U5070 ( .A(n2839), .B(n2847), .C(n2837), .Q(n2852) );
  OAI212 U5071 ( .A(n2848), .B(n2854), .C(n2851), .Q(n2853) );
  OAI212 U5072 ( .A(n2838), .B(n2856), .C(n2839), .Q(n2835) );
  IMAJ31 U5073 ( .A(\u_decoder/fir_filter/dp_cluster_0/r180/A2[7] ), .B(n2843), 
        .C(\u_decoder/fir_filter/dp_cluster_0/r180/A1[7] ), .Q(n2838) );
  OAI212 U5074 ( .A(n2860), .B(n2861), .C(n2862), .Q(
        \u_decoder/fir_filter/Q_data_mult_4 [10]) );
  XOR31 U5075 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_308/A1[7] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/A2[7] ), .C(n2865), .Q(
        \u_decoder/fir_filter/Q_data_mult_4 [9]) );
  OAI222 U5076 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[7][5] ), 
        .B(\u_decoder/fir_filter/dp_cluster_0/mult_308/A2[11] ), .C(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/A1[8] ), .D(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/A2[8] ), .Q(n2871) );
  OAI212 U5077 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[7][5] ), 
        .B(n2867), .C(\u_decoder/fir_filter/dp_cluster_0/mult_308/A2[11] ), 
        .Q(n2872) );
  OAI212 U5078 ( .A(n2870), .B(n2334), .C(n2873), .Q(n2867) );
  OAI212 U5079 ( .A(n2861), .B(n2869), .C(n2859), .Q(n2874) );
  XOR31 U5080 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_308/A2[11] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/mult_308/CARRYB[7][5] ), .C(n2875), 
        .Q(\u_decoder/fir_filter/Q_data_mult_4 [13]) );
  OAI212 U5081 ( .A(n2870), .B(n2876), .C(n2873), .Q(n2875) );
  OAI212 U5082 ( .A(n2860), .B(n2878), .C(n2861), .Q(n2857) );
  IMAJ31 U5083 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_308/A2[7] ), .B(
        n2865), .C(\u_decoder/fir_filter/dp_cluster_0/mult_308/A1[7] ), .Q(
        n2860) );
  OAI212 U5084 ( .A(\u_decoder/fir_filter/dp_cluster_0/r164/A1[6] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r164/A2[6] ), .C(n2884), .Q(n2883)
         );
  OAI212 U5085 ( .A(\u_decoder/fir_filter/dp_cluster_0/r164/A2[6] ), .B(n2885), 
        .C(n2886), .Q(\u_decoder/fir_filter/I_data_mult_0 [8]) );
  OAI212 U5086 ( .A(\u_decoder/fir_filter/dp_cluster_0/r164/PROD1[4] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r164/A1[3] ), .C(n2888), .Q(n2890)
         );
  OAI212 U5087 ( .A(n2305), .B(n2879), .C(
        \u_decoder/fir_filter/dp_cluster_0/r164/A2[9] ), .Q(n2892) );
  OAI212 U5088 ( .A(n2880), .B(n2297), .C(n2893), .Q(n2879) );
  OAI212 U5089 ( .A(\u_decoder/fir_filter/dp_cluster_0/r164/A1[8] ), .B(n2290), 
        .C(\u_decoder/fir_filter/dp_cluster_0/r164/A2[8] ), .Q(n2893) );
  OAI222 U5090 ( .A(\u_decoder/fir_filter/dp_cluster_0/r164/A1[6] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r164/A2[6] ), .C(
        \u_decoder/fir_filter/dp_cluster_0/r164/A1[7] ), .D(
        \u_decoder/fir_filter/dp_cluster_0/r164/A2[7] ), .Q(n2896) );
  OAI212 U5091 ( .A(\u_decoder/fir_filter/dp_cluster_0/r165/PROD1[5] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/r165/A1[4] ), .C(n2902), .Q(n2904)
         );
  OAI212 U5092 ( .A(n2305), .B(n2906), .C(
        \u_decoder/fir_filter/dp_cluster_0/r165/A2[10] ), .Q(n2907) );
  OAI212 U5093 ( .A(n2239), .B(n2238), .C(n2908), .Q(n2906) );
  OAI212 U5094 ( .A(\u_decoder/fir_filter/dp_cluster_0/r165/A1[9] ), .B(n2897), 
        .C(\u_decoder/fir_filter/dp_cluster_0/r165/A2[9] ), .Q(n2908) );
  OAI212 U5095 ( .A(n2898), .B(n2240), .C(n2909), .Q(n2897) );
  OAI212 U5096 ( .A(\u_decoder/fir_filter/dp_cluster_0/r165/A1[8] ), .B(n2241), 
        .C(\u_decoder/fir_filter/dp_cluster_0/r165/A2[8] ), .Q(n2909) );
  OAI212 U5097 ( .A(\u_decoder/fir_filter/dp_cluster_0/r165/A1[7] ), .B(n2899), 
        .C(\u_decoder/fir_filter/dp_cluster_0/r165/A2[7] ), .Q(n2910) );
  OAI212 U5098 ( .A(n2246), .B(n2245), .C(n2917), .Q(n2916) );
  OAI212 U5099 ( .A(\u_decoder/fir_filter/dp_cluster_0/r166/CARRYB[7][3] ), 
        .B(n2912), .C(\u_decoder/fir_filter/dp_cluster_0/r166/A2[9] ), .Q(
        n2917) );
  OAI212 U5100 ( .A(n2913), .B(n2247), .C(n2918), .Q(n2912) );
  OAI212 U5101 ( .A(\u_decoder/fir_filter/dp_cluster_0/r166/A1[8] ), .B(n2248), 
        .C(\u_decoder/fir_filter/dp_cluster_0/r166/A2[8] ), .Q(n2918) );
  OAI212 U5102 ( .A(\u_decoder/fir_filter/dp_cluster_0/r166/A1[7] ), .B(n2251), 
        .C(\u_decoder/fir_filter/dp_cluster_0/r166/A2[7] ), .Q(n2919) );
  OAI212 U5103 ( .A(n2924), .B(n2925), .C(n2926), .Q(
        \u_decoder/fir_filter/I_data_mult_3 [10]) );
  OAI222 U5104 ( .A(\u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[7][5] ), 
        .B(\u_decoder/fir_filter/dp_cluster_0/r167/A2[11] ), .C(
        \u_decoder/fir_filter/dp_cluster_0/r167/A1[8] ), .D(
        \u_decoder/fir_filter/dp_cluster_0/r167/A2[8] ), .Q(n2935) );
  OAI212 U5105 ( .A(\u_decoder/fir_filter/dp_cluster_0/r167/CARRYB[7][5] ), 
        .B(n2931), .C(\u_decoder/fir_filter/dp_cluster_0/r167/A2[11] ), .Q(
        n2936) );
  OAI212 U5106 ( .A(n2934), .B(n2279), .C(n2937), .Q(n2931) );
  OAI212 U5107 ( .A(n2925), .B(n2933), .C(n2923), .Q(n2938) );
  OAI212 U5108 ( .A(n2934), .B(n2940), .C(n2937), .Q(n2939) );
  OAI212 U5109 ( .A(n2924), .B(n2942), .C(n2925), .Q(n2921) );
  IMAJ31 U5110 ( .A(\u_decoder/fir_filter/dp_cluster_0/r167/A2[7] ), .B(n2929), 
        .C(\u_decoder/fir_filter/dp_cluster_0/r167/A1[7] ), .Q(n2924) );
  OAI212 U5111 ( .A(n2946), .B(n2947), .C(n2948), .Q(
        \u_decoder/fir_filter/I_data_mult_4 [10]) );
  XOR31 U5112 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_276/A1[7] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/A2[7] ), .C(n2951), .Q(
        \u_decoder/fir_filter/I_data_mult_4 [9]) );
  OAI222 U5113 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[7][5] ), 
        .B(\u_decoder/fir_filter/dp_cluster_0/mult_276/A2[11] ), .C(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/A1[8] ), .D(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/A2[8] ), .Q(n2957) );
  OAI212 U5114 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[7][5] ), 
        .B(n2953), .C(\u_decoder/fir_filter/dp_cluster_0/mult_276/A2[11] ), 
        .Q(n2958) );
  OAI212 U5115 ( .A(n2956), .B(n2263), .C(n2959), .Q(n2953) );
  OAI212 U5116 ( .A(n2947), .B(n2955), .C(n2945), .Q(n2960) );
  XOR31 U5117 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_276/A2[11] ), .B(
        \u_decoder/fir_filter/dp_cluster_0/mult_276/CARRYB[7][5] ), .C(n2961), 
        .Q(\u_decoder/fir_filter/I_data_mult_4 [13]) );
  OAI212 U5118 ( .A(n2956), .B(n2962), .C(n2959), .Q(n2961) );
  OAI212 U5119 ( .A(n2946), .B(n2964), .C(n2947), .Q(n2943) );
  IMAJ31 U5120 ( .A(\u_decoder/fir_filter/dp_cluster_0/mult_276/A2[7] ), .B(
        n2951), .C(\u_decoder/fir_filter/dp_cluster_0/mult_276/A1[7] ), .Q(
        n2946) );
  OAI212 U5121 ( .A(n93), .B(n24), .C(n2965), .Q(n2966) );
  OAI212 U5122 ( .A(\u_decoder/fir_filter/Q_data_mult_0_buff [2]), .B(n2966), 
        .C(\u_decoder/fir_filter/Q_data_add_1_buff [2]), .Q(n2967) );
  OAI212 U5123 ( .A(n2424), .B(n91), .C(n2967), .Q(n2968) );
  OAI212 U5124 ( .A(\u_decoder/fir_filter/Q_data_mult_0_buff [3]), .B(n2968), 
        .C(\u_decoder/fir_filter/Q_data_add_1_buff [3]), .Q(n2969) );
  OAI212 U5125 ( .A(n2422), .B(n135), .C(n2969), .Q(n2970) );
  OAI212 U5126 ( .A(\u_decoder/fir_filter/Q_data_mult_0_buff [4]), .B(n2970), 
        .C(\u_decoder/fir_filter/Q_data_add_1_buff [4]), .Q(n2971) );
  OAI212 U5127 ( .A(n2420), .B(n136), .C(n2971), .Q(n2972) );
  OAI212 U5128 ( .A(\u_decoder/fir_filter/Q_data_mult_0_buff [5]), .B(n2972), 
        .C(\u_decoder/fir_filter/Q_data_add_1_buff [5]), .Q(n2973) );
  OAI212 U5129 ( .A(n2418), .B(n137), .C(n2973), .Q(n2974) );
  OAI212 U5130 ( .A(\u_decoder/fir_filter/Q_data_mult_0_buff [6]), .B(n2974), 
        .C(\u_decoder/fir_filter/Q_data_add_1_buff [6]), .Q(n2975) );
  OAI212 U5131 ( .A(n2416), .B(n177), .C(n2975), .Q(n2977) );
  OAI212 U5132 ( .A(\u_decoder/fir_filter/Q_data_mult_0_buff [7]), .B(n2977), 
        .C(\u_decoder/fir_filter/Q_data_add_1_buff [7]), .Q(n2976) );
  OAI212 U5133 ( .A(\u_decoder/fir_filter/Q_data_mult_0_buff [8]), .B(n2412), 
        .C(\u_decoder/fir_filter/Q_data_add_1_buff [8]), .Q(n2978) );
  OAI212 U5134 ( .A(n2979), .B(n223), .C(n2978), .Q(n2981) );
  OAI212 U5135 ( .A(\u_decoder/fir_filter/Q_data_mult_0_buff [9]), .B(n2981), 
        .C(\u_decoder/fir_filter/Q_data_add_1_buff [9]), .Q(n2980) );
  OAI212 U5136 ( .A(\u_decoder/fir_filter/Q_data_mult_0_buff [10]), .B(n2408), 
        .C(\u_decoder/fir_filter/Q_data_add_1_buff [10]), .Q(n2982) );
  OAI212 U5137 ( .A(n2983), .B(n264), .C(n2982), .Q(
        \u_decoder/fir_filter/add_326/carry [11]) );
  OAI212 U5138 ( .A(n94), .B(n25), .C(n2984), .Q(n2985) );
  OAI212 U5139 ( .A(\u_decoder/fir_filter/I_data_mult_0_buff [2]), .B(n2985), 
        .C(\u_decoder/fir_filter/I_data_add_1_buff [2]), .Q(n2986) );
  OAI212 U5140 ( .A(n2544), .B(n92), .C(n2986), .Q(n2987) );
  OAI212 U5141 ( .A(\u_decoder/fir_filter/I_data_mult_0_buff [3]), .B(n2987), 
        .C(\u_decoder/fir_filter/I_data_add_1_buff [3]), .Q(n2988) );
  OAI212 U5142 ( .A(n2542), .B(n138), .C(n2988), .Q(n2989) );
  OAI212 U5143 ( .A(\u_decoder/fir_filter/I_data_mult_0_buff [4]), .B(n2989), 
        .C(\u_decoder/fir_filter/I_data_add_1_buff [4]), .Q(n2990) );
  OAI212 U5144 ( .A(n2540), .B(n139), .C(n2990), .Q(n2991) );
  OAI212 U5145 ( .A(\u_decoder/fir_filter/I_data_mult_0_buff [5]), .B(n2991), 
        .C(\u_decoder/fir_filter/I_data_add_1_buff [5]), .Q(n2992) );
  OAI212 U5146 ( .A(n2538), .B(n140), .C(n2992), .Q(n2993) );
  OAI212 U5147 ( .A(\u_decoder/fir_filter/I_data_mult_0_buff [6]), .B(n2993), 
        .C(\u_decoder/fir_filter/I_data_add_1_buff [6]), .Q(n2994) );
  OAI212 U5148 ( .A(n2536), .B(n178), .C(n2994), .Q(n2996) );
  OAI212 U5149 ( .A(\u_decoder/fir_filter/I_data_mult_0_buff [7]), .B(n2996), 
        .C(\u_decoder/fir_filter/I_data_add_1_buff [7]), .Q(n2995) );
  OAI212 U5150 ( .A(\u_decoder/fir_filter/I_data_mult_0_buff [8]), .B(n2532), 
        .C(\u_decoder/fir_filter/I_data_add_1_buff [8]), .Q(n2997) );
  OAI212 U5151 ( .A(n2998), .B(n224), .C(n2997), .Q(n3000) );
  OAI212 U5152 ( .A(\u_decoder/fir_filter/I_data_mult_0_buff [9]), .B(n3000), 
        .C(\u_decoder/fir_filter/I_data_add_1_buff [9]), .Q(n2999) );
  OAI212 U5153 ( .A(\u_decoder/fir_filter/I_data_mult_0_buff [10]), .B(n2528), 
        .C(\u_decoder/fir_filter/I_data_add_1_buff [10]), .Q(n3001) );
  OAI212 U5154 ( .A(n3002), .B(n265), .C(n3001), .Q(
        \u_decoder/fir_filter/add_294/carry [11]) );
  OAI212 U5155 ( .A(n225), .B(n46), .C(n3003), .Q(n3004) );
  OAI212 U5156 ( .A(\u_cordic/mycordic/present_Q_table[5][2] ), .B(n3004), .C(
        \u_cordic/mycordic/present_I_table[5][6] ), .Q(n3005) );
  OAI212 U5157 ( .A(n2649), .B(n197), .C(n3005), .Q(n3007) );
  OAI212 U5158 ( .A(\u_cordic/mycordic/present_Q_table[5][3] ), .B(n3007), .C(
        \u_cordic/mycordic/present_I_table[5][7] ), .Q(n3006) );
  OAI212 U5159 ( .A(\u_cordic/mycordic/present_Q_table[5][4] ), .B(n2645), .C(
        \u_cordic/mycordic/present_I_table[5][7] ), .Q(n3008) );
  OAI212 U5160 ( .A(n3009), .B(n247), .C(n3008), .Q(n3011) );
  OAI212 U5161 ( .A(\u_cordic/mycordic/present_Q_table[5][5] ), .B(n3011), .C(
        \u_cordic/mycordic/present_I_table[5][7] ), .Q(n3010) );
  OAI212 U5162 ( .A(\u_cordic/mycordic/present_Q_table[5][6] ), .B(n2641), .C(
        \u_cordic/mycordic/present_I_table[5][7] ), .Q(n3012) );
  OAI212 U5163 ( .A(n3013), .B(n286), .C(n3012), .Q(
        \u_cordic/mycordic/add_228/carry[7] ) );
  OAI222 U5164 ( .A(n3017), .B(n197), .C(
        \u_cordic/mycordic/present_I_table[5][6] ), .D(n2648), .Q(n3019) );
  OAI212 U5165 ( .A(\u_cordic/mycordic/present_Q_table[5][3] ), .B(n3019), .C(
        n199), .Q(n3018) );
  OAI212 U5166 ( .A(n3021), .B(n247), .C(n2644), .Q(n3023) );
  OAI212 U5167 ( .A(\u_cordic/mycordic/present_Q_table[5][5] ), .B(n3023), .C(
        n199), .Q(n3022) );
  OAI212 U5168 ( .A(n3025), .B(n286), .C(n2640), .Q(
        \u_cordic/mycordic/sub_223/carry[7] ) );
  OAI222 U5169 ( .A(n3027), .B(n226), .C(
        \u_cordic/mycordic/present_Q_table[4][4] ), .D(n3026), .Q(n3029) );
  OAI222 U5170 ( .A(n3031), .B(n163), .C(
        \u_cordic/mycordic/present_Q_table[4][6] ), .D(n3030), .Q(
        \u_cordic/mycordic/sub_216/carry [4]) );
  OAI212 U5171 ( .A(\u_cordic/mycordic/present_I_table[4][2] ), .B(n2656), .C(
        \u_cordic/mycordic/present_Q_table[4][5] ), .Q(n3033) );
  OAI212 U5172 ( .A(n3034), .B(n222), .C(n3033), .Q(n3036) );
  OAI212 U5173 ( .A(\u_cordic/mycordic/present_I_table[4][3] ), .B(n3036), .C(
        \u_cordic/mycordic/present_Q_table[4][6] ), .Q(n3035) );
  OAI222 U5174 ( .A(n1399), .B(n293), .C(n1400), .D(n1399), .Q(n3049) );
  OAI212 U5175 ( .A(\u_coder/n241 ), .B(\u_coder/n88 ), .C(\u_coder/stateQ[0] ), .Q(\u_coder/N1149 ) );
  OAI212 U5176 ( .A(\u_coder/n242 ), .B(\u_coder/n88 ), .C(\u_coder/stateI[0] ), .Q(\u_coder/N1143 ) );
endmodule

